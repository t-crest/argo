module Xbar
  (input  [19:0] func,
   input  [179:0] inPort,
   output [179:0] outPort);
  wire [3:0] sel0;
  wire [3:0] sel1;
  wire [3:0] sel2;
  wire [3:0] sel3;
  wire [3:0] sel4;
  wire [3:0] n1_o;
  wire [3:0] n2_o;
  wire [3:0] n3_o;
  wire [3:0] n4_o;
  wire [3:0] n5_o;
  wire [35:0] n6_o;
  wire [34:0] n7_o;
  wire n8_o;
  wire n9_o;
  wire n10_o;
  wire n11_o;
  wire n12_o;
  wire n13_o;
  wire n14_o;
  wire n15_o;
  wire n16_o;
  wire n17_o;
  wire n18_o;
  wire n19_o;
  wire n20_o;
  wire n21_o;
  wire n22_o;
  wire n23_o;
  wire n24_o;
  wire n25_o;
  wire n26_o;
  wire n27_o;
  wire n28_o;
  wire n29_o;
  wire n30_o;
  wire n31_o;
  wire n32_o;
  wire n33_o;
  wire n34_o;
  wire n35_o;
  wire n36_o;
  wire n37_o;
  wire n38_o;
  wire n39_o;
  wire n40_o;
  wire n41_o;
  wire n42_o;
  wire [3:0] n43_o;
  wire [3:0] n44_o;
  wire [3:0] n45_o;
  wire [3:0] n46_o;
  wire [3:0] n47_o;
  wire [3:0] n48_o;
  wire [3:0] n49_o;
  wire [3:0] n50_o;
  wire [2:0] n51_o;
  wire [15:0] n52_o;
  wire [15:0] n53_o;
  wire [34:0] n54_o;
  wire [34:0] n55_o;
  wire [35:0] n56_o;
  wire [34:0] n57_o;
  wire n58_o;
  wire n59_o;
  wire n60_o;
  wire n61_o;
  wire n62_o;
  wire n63_o;
  wire n64_o;
  wire n65_o;
  wire n66_o;
  wire n67_o;
  wire n68_o;
  wire n69_o;
  wire n70_o;
  wire n71_o;
  wire n72_o;
  wire n73_o;
  wire n74_o;
  wire n75_o;
  wire n76_o;
  wire n77_o;
  wire n78_o;
  wire n79_o;
  wire n80_o;
  wire n81_o;
  wire n82_o;
  wire n83_o;
  wire n84_o;
  wire n85_o;
  wire n86_o;
  wire n87_o;
  wire n88_o;
  wire n89_o;
  wire n90_o;
  wire n91_o;
  wire n92_o;
  wire [3:0] n93_o;
  wire [3:0] n94_o;
  wire [3:0] n95_o;
  wire [3:0] n96_o;
  wire [3:0] n97_o;
  wire [3:0] n98_o;
  wire [3:0] n99_o;
  wire [3:0] n100_o;
  wire [2:0] n101_o;
  wire [15:0] n102_o;
  wire [15:0] n103_o;
  wire [34:0] n104_o;
  wire [34:0] n105_o;
  wire [34:0] n106_o;
  wire [35:0] n107_o;
  wire [34:0] n108_o;
  wire n109_o;
  wire n110_o;
  wire n111_o;
  wire n112_o;
  wire n113_o;
  wire n114_o;
  wire n115_o;
  wire n116_o;
  wire n117_o;
  wire n118_o;
  wire n119_o;
  wire n120_o;
  wire n121_o;
  wire n122_o;
  wire n123_o;
  wire n124_o;
  wire n125_o;
  wire n126_o;
  wire n127_o;
  wire n128_o;
  wire n129_o;
  wire n130_o;
  wire n131_o;
  wire n132_o;
  wire n133_o;
  wire n134_o;
  wire n135_o;
  wire n136_o;
  wire n137_o;
  wire n138_o;
  wire n139_o;
  wire n140_o;
  wire n141_o;
  wire n142_o;
  wire n143_o;
  wire [3:0] n144_o;
  wire [3:0] n145_o;
  wire [3:0] n146_o;
  wire [3:0] n147_o;
  wire [3:0] n148_o;
  wire [3:0] n149_o;
  wire [3:0] n150_o;
  wire [3:0] n151_o;
  wire [2:0] n152_o;
  wire [15:0] n153_o;
  wire [15:0] n154_o;
  wire [34:0] n155_o;
  wire [34:0] n156_o;
  wire [34:0] n157_o;
  wire [35:0] n158_o;
  wire [34:0] n159_o;
  wire n160_o;
  wire n161_o;
  wire n162_o;
  wire n163_o;
  wire n164_o;
  wire n165_o;
  wire n166_o;
  wire n167_o;
  wire n168_o;
  wire n169_o;
  wire n170_o;
  wire n171_o;
  wire n172_o;
  wire n173_o;
  wire n174_o;
  wire n175_o;
  wire n176_o;
  wire n177_o;
  wire n178_o;
  wire n179_o;
  wire n180_o;
  wire n181_o;
  wire n182_o;
  wire n183_o;
  wire n184_o;
  wire n185_o;
  wire n186_o;
  wire n187_o;
  wire n188_o;
  wire n189_o;
  wire n190_o;
  wire n191_o;
  wire n192_o;
  wire n193_o;
  wire n194_o;
  wire [3:0] n195_o;
  wire [3:0] n196_o;
  wire [3:0] n197_o;
  wire [3:0] n198_o;
  wire [3:0] n199_o;
  wire [3:0] n200_o;
  wire [3:0] n201_o;
  wire [3:0] n202_o;
  wire [2:0] n203_o;
  wire [15:0] n204_o;
  wire [15:0] n205_o;
  wire [34:0] n206_o;
  wire [34:0] n207_o;
  wire [34:0] n208_o;
  wire [35:0] n209_o;
  wire [34:0] n210_o;
  wire n211_o;
  wire n212_o;
  wire n213_o;
  wire n214_o;
  wire n215_o;
  wire n216_o;
  wire n217_o;
  wire n218_o;
  wire n219_o;
  wire n220_o;
  wire n221_o;
  wire n222_o;
  wire n223_o;
  wire n224_o;
  wire n225_o;
  wire n226_o;
  wire n227_o;
  wire n228_o;
  wire n229_o;
  wire n230_o;
  wire n231_o;
  wire n232_o;
  wire n233_o;
  wire n234_o;
  wire n235_o;
  wire n236_o;
  wire n237_o;
  wire n238_o;
  wire n239_o;
  wire n240_o;
  wire n241_o;
  wire n242_o;
  wire n243_o;
  wire n244_o;
  wire n245_o;
  wire [3:0] n246_o;
  wire [3:0] n247_o;
  wire [3:0] n248_o;
  wire [3:0] n249_o;
  wire [3:0] n250_o;
  wire [3:0] n251_o;
  wire [3:0] n252_o;
  wire [3:0] n253_o;
  wire [2:0] n254_o;
  wire [15:0] n255_o;
  wire [15:0] n256_o;
  wire [34:0] n257_o;
  wire [34:0] n258_o;
  wire [35:0] n259_o;
  wire [34:0] n260_o;
  wire n261_o;
  wire n262_o;
  wire n263_o;
  wire n264_o;
  wire n265_o;
  wire n266_o;
  wire n267_o;
  wire n268_o;
  wire n269_o;
  wire n270_o;
  wire n271_o;
  wire n272_o;
  wire n273_o;
  wire n274_o;
  wire n275_o;
  wire n276_o;
  wire n277_o;
  wire n278_o;
  wire n279_o;
  wire n280_o;
  wire n281_o;
  wire n282_o;
  wire n283_o;
  wire n284_o;
  wire n285_o;
  wire n286_o;
  wire n287_o;
  wire n288_o;
  wire n289_o;
  wire n290_o;
  wire n291_o;
  wire n292_o;
  wire n293_o;
  wire n294_o;
  wire n295_o;
  wire [3:0] n296_o;
  wire [3:0] n297_o;
  wire [3:0] n298_o;
  wire [3:0] n299_o;
  wire [3:0] n300_o;
  wire [3:0] n301_o;
  wire [3:0] n302_o;
  wire [3:0] n303_o;
  wire [2:0] n304_o;
  wire [15:0] n305_o;
  wire [15:0] n306_o;
  wire [34:0] n307_o;
  wire [34:0] n308_o;
  wire [34:0] n309_o;
  wire [35:0] n310_o;
  wire [34:0] n311_o;
  wire n312_o;
  wire n313_o;
  wire n314_o;
  wire n315_o;
  wire n316_o;
  wire n317_o;
  wire n318_o;
  wire n319_o;
  wire n320_o;
  wire n321_o;
  wire n322_o;
  wire n323_o;
  wire n324_o;
  wire n325_o;
  wire n326_o;
  wire n327_o;
  wire n328_o;
  wire n329_o;
  wire n330_o;
  wire n331_o;
  wire n332_o;
  wire n333_o;
  wire n334_o;
  wire n335_o;
  wire n336_o;
  wire n337_o;
  wire n338_o;
  wire n339_o;
  wire n340_o;
  wire n341_o;
  wire n342_o;
  wire n343_o;
  wire n344_o;
  wire n345_o;
  wire n346_o;
  wire [3:0] n347_o;
  wire [3:0] n348_o;
  wire [3:0] n349_o;
  wire [3:0] n350_o;
  wire [3:0] n351_o;
  wire [3:0] n352_o;
  wire [3:0] n353_o;
  wire [3:0] n354_o;
  wire [2:0] n355_o;
  wire [15:0] n356_o;
  wire [15:0] n357_o;
  wire [34:0] n358_o;
  wire [34:0] n359_o;
  wire [34:0] n360_o;
  wire [35:0] n361_o;
  wire [34:0] n362_o;
  wire n363_o;
  wire n364_o;
  wire n365_o;
  wire n366_o;
  wire n367_o;
  wire n368_o;
  wire n369_o;
  wire n370_o;
  wire n371_o;
  wire n372_o;
  wire n373_o;
  wire n374_o;
  wire n375_o;
  wire n376_o;
  wire n377_o;
  wire n378_o;
  wire n379_o;
  wire n380_o;
  wire n381_o;
  wire n382_o;
  wire n383_o;
  wire n384_o;
  wire n385_o;
  wire n386_o;
  wire n387_o;
  wire n388_o;
  wire n389_o;
  wire n390_o;
  wire n391_o;
  wire n392_o;
  wire n393_o;
  wire n394_o;
  wire n395_o;
  wire n396_o;
  wire n397_o;
  wire [3:0] n398_o;
  wire [3:0] n399_o;
  wire [3:0] n400_o;
  wire [3:0] n401_o;
  wire [3:0] n402_o;
  wire [3:0] n403_o;
  wire [3:0] n404_o;
  wire [3:0] n405_o;
  wire [2:0] n406_o;
  wire [15:0] n407_o;
  wire [15:0] n408_o;
  wire [34:0] n409_o;
  wire [34:0] n410_o;
  wire [34:0] n411_o;
  wire [35:0] n412_o;
  wire [34:0] n413_o;
  wire n414_o;
  wire n415_o;
  wire n416_o;
  wire n417_o;
  wire n418_o;
  wire n419_o;
  wire n420_o;
  wire n421_o;
  wire n422_o;
  wire n423_o;
  wire n424_o;
  wire n425_o;
  wire n426_o;
  wire n427_o;
  wire n428_o;
  wire n429_o;
  wire n430_o;
  wire n431_o;
  wire n432_o;
  wire n433_o;
  wire n434_o;
  wire n435_o;
  wire n436_o;
  wire n437_o;
  wire n438_o;
  wire n439_o;
  wire n440_o;
  wire n441_o;
  wire n442_o;
  wire n443_o;
  wire n444_o;
  wire n445_o;
  wire n446_o;
  wire n447_o;
  wire n448_o;
  wire [3:0] n449_o;
  wire [3:0] n450_o;
  wire [3:0] n451_o;
  wire [3:0] n452_o;
  wire [3:0] n453_o;
  wire [3:0] n454_o;
  wire [3:0] n455_o;
  wire [3:0] n456_o;
  wire [2:0] n457_o;
  wire [15:0] n458_o;
  wire [15:0] n459_o;
  wire [34:0] n460_o;
  wire [34:0] n461_o;
  wire [35:0] n462_o;
  wire [34:0] n463_o;
  wire n464_o;
  wire n465_o;
  wire n466_o;
  wire n467_o;
  wire n468_o;
  wire n469_o;
  wire n470_o;
  wire n471_o;
  wire n472_o;
  wire n473_o;
  wire n474_o;
  wire n475_o;
  wire n476_o;
  wire n477_o;
  wire n478_o;
  wire n479_o;
  wire n480_o;
  wire n481_o;
  wire n482_o;
  wire n483_o;
  wire n484_o;
  wire n485_o;
  wire n486_o;
  wire n487_o;
  wire n488_o;
  wire n489_o;
  wire n490_o;
  wire n491_o;
  wire n492_o;
  wire n493_o;
  wire n494_o;
  wire n495_o;
  wire n496_o;
  wire n497_o;
  wire n498_o;
  wire [3:0] n499_o;
  wire [3:0] n500_o;
  wire [3:0] n501_o;
  wire [3:0] n502_o;
  wire [3:0] n503_o;
  wire [3:0] n504_o;
  wire [3:0] n505_o;
  wire [3:0] n506_o;
  wire [2:0] n507_o;
  wire [15:0] n508_o;
  wire [15:0] n509_o;
  wire [34:0] n510_o;
  wire [34:0] n511_o;
  wire [34:0] n512_o;
  wire [35:0] n513_o;
  wire [34:0] n514_o;
  wire n515_o;
  wire n516_o;
  wire n517_o;
  wire n518_o;
  wire n519_o;
  wire n520_o;
  wire n521_o;
  wire n522_o;
  wire n523_o;
  wire n524_o;
  wire n525_o;
  wire n526_o;
  wire n527_o;
  wire n528_o;
  wire n529_o;
  wire n530_o;
  wire n531_o;
  wire n532_o;
  wire n533_o;
  wire n534_o;
  wire n535_o;
  wire n536_o;
  wire n537_o;
  wire n538_o;
  wire n539_o;
  wire n540_o;
  wire n541_o;
  wire n542_o;
  wire n543_o;
  wire n544_o;
  wire n545_o;
  wire n546_o;
  wire n547_o;
  wire n548_o;
  wire n549_o;
  wire [3:0] n550_o;
  wire [3:0] n551_o;
  wire [3:0] n552_o;
  wire [3:0] n553_o;
  wire [3:0] n554_o;
  wire [3:0] n555_o;
  wire [3:0] n556_o;
  wire [3:0] n557_o;
  wire [2:0] n558_o;
  wire [15:0] n559_o;
  wire [15:0] n560_o;
  wire [34:0] n561_o;
  wire [34:0] n562_o;
  wire [34:0] n563_o;
  wire [35:0] n564_o;
  wire [34:0] n565_o;
  wire n566_o;
  wire n567_o;
  wire n568_o;
  wire n569_o;
  wire n570_o;
  wire n571_o;
  wire n572_o;
  wire n573_o;
  wire n574_o;
  wire n575_o;
  wire n576_o;
  wire n577_o;
  wire n578_o;
  wire n579_o;
  wire n580_o;
  wire n581_o;
  wire n582_o;
  wire n583_o;
  wire n584_o;
  wire n585_o;
  wire n586_o;
  wire n587_o;
  wire n588_o;
  wire n589_o;
  wire n590_o;
  wire n591_o;
  wire n592_o;
  wire n593_o;
  wire n594_o;
  wire n595_o;
  wire n596_o;
  wire n597_o;
  wire n598_o;
  wire n599_o;
  wire n600_o;
  wire [3:0] n601_o;
  wire [3:0] n602_o;
  wire [3:0] n603_o;
  wire [3:0] n604_o;
  wire [3:0] n605_o;
  wire [3:0] n606_o;
  wire [3:0] n607_o;
  wire [3:0] n608_o;
  wire [2:0] n609_o;
  wire [15:0] n610_o;
  wire [15:0] n611_o;
  wire [34:0] n612_o;
  wire [34:0] n613_o;
  wire [34:0] n614_o;
  wire [35:0] n615_o;
  wire [34:0] n616_o;
  wire n617_o;
  wire n618_o;
  wire n619_o;
  wire n620_o;
  wire n621_o;
  wire n622_o;
  wire n623_o;
  wire n624_o;
  wire n625_o;
  wire n626_o;
  wire n627_o;
  wire n628_o;
  wire n629_o;
  wire n630_o;
  wire n631_o;
  wire n632_o;
  wire n633_o;
  wire n634_o;
  wire n635_o;
  wire n636_o;
  wire n637_o;
  wire n638_o;
  wire n639_o;
  wire n640_o;
  wire n641_o;
  wire n642_o;
  wire n643_o;
  wire n644_o;
  wire n645_o;
  wire n646_o;
  wire n647_o;
  wire n648_o;
  wire n649_o;
  wire n650_o;
  wire n651_o;
  wire [3:0] n652_o;
  wire [3:0] n653_o;
  wire [3:0] n654_o;
  wire [3:0] n655_o;
  wire [3:0] n656_o;
  wire [3:0] n657_o;
  wire [3:0] n658_o;
  wire [3:0] n659_o;
  wire [2:0] n660_o;
  wire [15:0] n661_o;
  wire [15:0] n662_o;
  wire [34:0] n663_o;
  wire [34:0] n664_o;
  wire [35:0] n665_o;
  wire [34:0] n666_o;
  wire n667_o;
  wire n668_o;
  wire n669_o;
  wire n670_o;
  wire n671_o;
  wire n672_o;
  wire n673_o;
  wire n674_o;
  wire n675_o;
  wire n676_o;
  wire n677_o;
  wire n678_o;
  wire n679_o;
  wire n680_o;
  wire n681_o;
  wire n682_o;
  wire n683_o;
  wire n684_o;
  wire n685_o;
  wire n686_o;
  wire n687_o;
  wire n688_o;
  wire n689_o;
  wire n690_o;
  wire n691_o;
  wire n692_o;
  wire n693_o;
  wire n694_o;
  wire n695_o;
  wire n696_o;
  wire n697_o;
  wire n698_o;
  wire n699_o;
  wire n700_o;
  wire n701_o;
  wire [3:0] n702_o;
  wire [3:0] n703_o;
  wire [3:0] n704_o;
  wire [3:0] n705_o;
  wire [3:0] n706_o;
  wire [3:0] n707_o;
  wire [3:0] n708_o;
  wire [3:0] n709_o;
  wire [2:0] n710_o;
  wire [15:0] n711_o;
  wire [15:0] n712_o;
  wire [34:0] n713_o;
  wire [34:0] n714_o;
  wire [34:0] n715_o;
  wire [35:0] n716_o;
  wire [34:0] n717_o;
  wire n718_o;
  wire n719_o;
  wire n720_o;
  wire n721_o;
  wire n722_o;
  wire n723_o;
  wire n724_o;
  wire n725_o;
  wire n726_o;
  wire n727_o;
  wire n728_o;
  wire n729_o;
  wire n730_o;
  wire n731_o;
  wire n732_o;
  wire n733_o;
  wire n734_o;
  wire n735_o;
  wire n736_o;
  wire n737_o;
  wire n738_o;
  wire n739_o;
  wire n740_o;
  wire n741_o;
  wire n742_o;
  wire n743_o;
  wire n744_o;
  wire n745_o;
  wire n746_o;
  wire n747_o;
  wire n748_o;
  wire n749_o;
  wire n750_o;
  wire n751_o;
  wire n752_o;
  wire [3:0] n753_o;
  wire [3:0] n754_o;
  wire [3:0] n755_o;
  wire [3:0] n756_o;
  wire [3:0] n757_o;
  wire [3:0] n758_o;
  wire [3:0] n759_o;
  wire [3:0] n760_o;
  wire [2:0] n761_o;
  wire [15:0] n762_o;
  wire [15:0] n763_o;
  wire [34:0] n764_o;
  wire [34:0] n765_o;
  wire [34:0] n766_o;
  wire [35:0] n767_o;
  wire [34:0] n768_o;
  wire n769_o;
  wire n770_o;
  wire n771_o;
  wire n772_o;
  wire n773_o;
  wire n774_o;
  wire n775_o;
  wire n776_o;
  wire n777_o;
  wire n778_o;
  wire n779_o;
  wire n780_o;
  wire n781_o;
  wire n782_o;
  wire n783_o;
  wire n784_o;
  wire n785_o;
  wire n786_o;
  wire n787_o;
  wire n788_o;
  wire n789_o;
  wire n790_o;
  wire n791_o;
  wire n792_o;
  wire n793_o;
  wire n794_o;
  wire n795_o;
  wire n796_o;
  wire n797_o;
  wire n798_o;
  wire n799_o;
  wire n800_o;
  wire n801_o;
  wire n802_o;
  wire n803_o;
  wire [3:0] n804_o;
  wire [3:0] n805_o;
  wire [3:0] n806_o;
  wire [3:0] n807_o;
  wire [3:0] n808_o;
  wire [3:0] n809_o;
  wire [3:0] n810_o;
  wire [3:0] n811_o;
  wire [2:0] n812_o;
  wire [15:0] n813_o;
  wire [15:0] n814_o;
  wire [34:0] n815_o;
  wire [34:0] n816_o;
  wire [34:0] n817_o;
  wire [35:0] n818_o;
  wire [34:0] n819_o;
  wire n820_o;
  wire n821_o;
  wire n822_o;
  wire n823_o;
  wire n824_o;
  wire n825_o;
  wire n826_o;
  wire n827_o;
  wire n828_o;
  wire n829_o;
  wire n830_o;
  wire n831_o;
  wire n832_o;
  wire n833_o;
  wire n834_o;
  wire n835_o;
  wire n836_o;
  wire n837_o;
  wire n838_o;
  wire n839_o;
  wire n840_o;
  wire n841_o;
  wire n842_o;
  wire n843_o;
  wire n844_o;
  wire n845_o;
  wire n846_o;
  wire n847_o;
  wire n848_o;
  wire n849_o;
  wire n850_o;
  wire n851_o;
  wire n852_o;
  wire n853_o;
  wire n854_o;
  wire [3:0] n855_o;
  wire [3:0] n856_o;
  wire [3:0] n857_o;
  wire [3:0] n858_o;
  wire [3:0] n859_o;
  wire [3:0] n860_o;
  wire [3:0] n861_o;
  wire [3:0] n862_o;
  wire [2:0] n863_o;
  wire [15:0] n864_o;
  wire [15:0] n865_o;
  wire [34:0] n866_o;
  wire [34:0] n867_o;
  wire [35:0] n868_o;
  wire [34:0] n869_o;
  wire n870_o;
  wire n871_o;
  wire n872_o;
  wire n873_o;
  wire n874_o;
  wire n875_o;
  wire n876_o;
  wire n877_o;
  wire n878_o;
  wire n879_o;
  wire n880_o;
  wire n881_o;
  wire n882_o;
  wire n883_o;
  wire n884_o;
  wire n885_o;
  wire n886_o;
  wire n887_o;
  wire n888_o;
  wire n889_o;
  wire n890_o;
  wire n891_o;
  wire n892_o;
  wire n893_o;
  wire n894_o;
  wire n895_o;
  wire n896_o;
  wire n897_o;
  wire n898_o;
  wire n899_o;
  wire n900_o;
  wire n901_o;
  wire n902_o;
  wire n903_o;
  wire n904_o;
  wire [3:0] n905_o;
  wire [3:0] n906_o;
  wire [3:0] n907_o;
  wire [3:0] n908_o;
  wire [3:0] n909_o;
  wire [3:0] n910_o;
  wire [3:0] n911_o;
  wire [3:0] n912_o;
  wire [2:0] n913_o;
  wire [15:0] n914_o;
  wire [15:0] n915_o;
  wire [34:0] n916_o;
  wire [34:0] n917_o;
  wire [34:0] n918_o;
  wire [35:0] n919_o;
  wire [34:0] n920_o;
  wire n921_o;
  wire n922_o;
  wire n923_o;
  wire n924_o;
  wire n925_o;
  wire n926_o;
  wire n927_o;
  wire n928_o;
  wire n929_o;
  wire n930_o;
  wire n931_o;
  wire n932_o;
  wire n933_o;
  wire n934_o;
  wire n935_o;
  wire n936_o;
  wire n937_o;
  wire n938_o;
  wire n939_o;
  wire n940_o;
  wire n941_o;
  wire n942_o;
  wire n943_o;
  wire n944_o;
  wire n945_o;
  wire n946_o;
  wire n947_o;
  wire n948_o;
  wire n949_o;
  wire n950_o;
  wire n951_o;
  wire n952_o;
  wire n953_o;
  wire n954_o;
  wire n955_o;
  wire [3:0] n956_o;
  wire [3:0] n957_o;
  wire [3:0] n958_o;
  wire [3:0] n959_o;
  wire [3:0] n960_o;
  wire [3:0] n961_o;
  wire [3:0] n962_o;
  wire [3:0] n963_o;
  wire [2:0] n964_o;
  wire [15:0] n965_o;
  wire [15:0] n966_o;
  wire [34:0] n967_o;
  wire [34:0] n968_o;
  wire [34:0] n969_o;
  wire [35:0] n970_o;
  wire [34:0] n971_o;
  wire n972_o;
  wire n973_o;
  wire n974_o;
  wire n975_o;
  wire n976_o;
  wire n977_o;
  wire n978_o;
  wire n979_o;
  wire n980_o;
  wire n981_o;
  wire n982_o;
  wire n983_o;
  wire n984_o;
  wire n985_o;
  wire n986_o;
  wire n987_o;
  wire n988_o;
  wire n989_o;
  wire n990_o;
  wire n991_o;
  wire n992_o;
  wire n993_o;
  wire n994_o;
  wire n995_o;
  wire n996_o;
  wire n997_o;
  wire n998_o;
  wire n999_o;
  wire n1000_o;
  wire n1001_o;
  wire n1002_o;
  wire n1003_o;
  wire n1004_o;
  wire n1005_o;
  wire n1006_o;
  wire [3:0] n1007_o;
  wire [3:0] n1008_o;
  wire [3:0] n1009_o;
  wire [3:0] n1010_o;
  wire [3:0] n1011_o;
  wire [3:0] n1012_o;
  wire [3:0] n1013_o;
  wire [3:0] n1014_o;
  wire [2:0] n1015_o;
  wire [15:0] n1016_o;
  wire [15:0] n1017_o;
  wire [34:0] n1018_o;
  wire [34:0] n1019_o;
  wire [34:0] n1020_o;
  wire [179:0] n1026_o;
  assign outPort = n1026_o;
  /* routers/synchronous/xbar.vhd:59:16  */
  assign sel0 = n1_o; // (signal)
  /* routers/synchronous/xbar.vhd:59:22  */
  assign sel1 = n2_o; // (signal)
  /* routers/synchronous/xbar.vhd:59:28  */
  assign sel2 = n3_o; // (signal)
  /* routers/synchronous/xbar.vhd:59:34  */
  assign sel3 = n4_o; // (signal)
  /* routers/synchronous/xbar.vhd:59:40  */
  assign sel4 = n5_o; // (signal)
  /* routers/synchronous/xbar.vhd:61:21  */
  assign n1_o = func[3:0];
  /* routers/synchronous/xbar.vhd:62:21  */
  assign n2_o = func[7:4];
  /* routers/synchronous/xbar.vhd:63:21  */
  assign n3_o = func[11:8];
  /* routers/synchronous/xbar.vhd:64:21  */
  assign n4_o = func[15:12];
  /* routers/synchronous/xbar.vhd:65:21  */
  assign n5_o = func[19:16];
  /* routers/synchronous/xbar.vhd:67:35  */
  assign n6_o = inPort[71:36];
  /* routers/synchronous/xbar.vhd:67:39  */
  assign n7_o = n6_o[35:1];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n8_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n9_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n10_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n11_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n12_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n13_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n14_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n15_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n16_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n17_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n18_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n19_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n20_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n21_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n22_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n23_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n24_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n25_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n26_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n27_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n28_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n29_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n30_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n31_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n32_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n33_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n34_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n35_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n36_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n37_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n38_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n39_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n40_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n41_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n42_o = sel1[0];
  assign n43_o = {n42_o, n41_o, n40_o, n39_o};
  assign n44_o = {n38_o, n37_o, n36_o, n35_o};
  assign n45_o = {n34_o, n33_o, n32_o, n31_o};
  assign n46_o = {n30_o, n29_o, n28_o, n27_o};
  assign n47_o = {n26_o, n25_o, n24_o, n23_o};
  assign n48_o = {n22_o, n21_o, n20_o, n19_o};
  assign n49_o = {n18_o, n17_o, n16_o, n15_o};
  assign n50_o = {n14_o, n13_o, n12_o, n11_o};
  assign n51_o = {n10_o, n9_o, n8_o};
  assign n52_o = {n43_o, n44_o, n45_o, n46_o};
  assign n53_o = {n47_o, n48_o, n49_o, n50_o};
  assign n54_o = {n52_o, n53_o, n51_o};
  /* routers/synchronous/xbar.vhd:67:44  */
  assign n55_o = n7_o & n54_o;
  /* routers/synchronous/xbar.vhd:68:42  */
  assign n56_o = inPort[107:72];
  /* routers/synchronous/xbar.vhd:68:46  */
  assign n57_o = n56_o[35:1];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n58_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n59_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n60_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n61_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n62_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n63_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n64_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n65_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n66_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n67_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n68_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n69_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n70_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n71_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n72_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n73_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n74_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n75_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n76_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n77_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n78_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n79_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n80_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n81_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n82_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n83_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n84_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n85_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n86_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n87_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n88_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n89_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n90_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n91_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n92_o = sel2[0];
  assign n93_o = {n92_o, n91_o, n90_o, n89_o};
  assign n94_o = {n88_o, n87_o, n86_o, n85_o};
  assign n95_o = {n84_o, n83_o, n82_o, n81_o};
  assign n96_o = {n80_o, n79_o, n78_o, n77_o};
  assign n97_o = {n76_o, n75_o, n74_o, n73_o};
  assign n98_o = {n72_o, n71_o, n70_o, n69_o};
  assign n99_o = {n68_o, n67_o, n66_o, n65_o};
  assign n100_o = {n64_o, n63_o, n62_o, n61_o};
  assign n101_o = {n60_o, n59_o, n58_o};
  assign n102_o = {n93_o, n94_o, n95_o, n96_o};
  assign n103_o = {n97_o, n98_o, n99_o, n100_o};
  assign n104_o = {n102_o, n103_o, n101_o};
  /* routers/synchronous/xbar.vhd:68:51  */
  assign n105_o = n57_o & n104_o;
  /* routers/synchronous/xbar.vhd:67:73  */
  assign n106_o = n55_o | n105_o;
  /* routers/synchronous/xbar.vhd:69:42  */
  assign n107_o = inPort[143:108];
  /* routers/synchronous/xbar.vhd:69:46  */
  assign n108_o = n107_o[35:1];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n109_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n110_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n111_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n112_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n113_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n114_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n115_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n116_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n117_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n118_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n119_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n120_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n121_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n122_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n123_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n124_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n125_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n126_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n127_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n128_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n129_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n130_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n131_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n132_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n133_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n134_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n135_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n136_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n137_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n138_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n139_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n140_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n141_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n142_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n143_o = sel3[0];
  assign n144_o = {n143_o, n142_o, n141_o, n140_o};
  assign n145_o = {n139_o, n138_o, n137_o, n136_o};
  assign n146_o = {n135_o, n134_o, n133_o, n132_o};
  assign n147_o = {n131_o, n130_o, n129_o, n128_o};
  assign n148_o = {n127_o, n126_o, n125_o, n124_o};
  assign n149_o = {n123_o, n122_o, n121_o, n120_o};
  assign n150_o = {n119_o, n118_o, n117_o, n116_o};
  assign n151_o = {n115_o, n114_o, n113_o, n112_o};
  assign n152_o = {n111_o, n110_o, n109_o};
  assign n153_o = {n144_o, n145_o, n146_o, n147_o};
  assign n154_o = {n148_o, n149_o, n150_o, n151_o};
  assign n155_o = {n153_o, n154_o, n152_o};
  /* routers/synchronous/xbar.vhd:69:51  */
  assign n156_o = n108_o & n155_o;
  /* routers/synchronous/xbar.vhd:68:80  */
  assign n157_o = n106_o | n156_o;
  /* routers/synchronous/xbar.vhd:70:42  */
  assign n158_o = inPort[179:144];
  /* routers/synchronous/xbar.vhd:70:46  */
  assign n159_o = n158_o[35:1];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n160_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n161_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n162_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n163_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n164_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n165_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n166_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n167_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n168_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n169_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n170_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n171_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n172_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n173_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n174_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n175_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n176_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n177_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n178_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n179_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n180_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n181_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n182_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n183_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n184_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n185_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n186_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n187_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n188_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n189_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n190_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n191_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n192_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n193_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n194_o = sel4[0];
  assign n195_o = {n194_o, n193_o, n192_o, n191_o};
  assign n196_o = {n190_o, n189_o, n188_o, n187_o};
  assign n197_o = {n186_o, n185_o, n184_o, n183_o};
  assign n198_o = {n182_o, n181_o, n180_o, n179_o};
  assign n199_o = {n178_o, n177_o, n176_o, n175_o};
  assign n200_o = {n174_o, n173_o, n172_o, n171_o};
  assign n201_o = {n170_o, n169_o, n168_o, n167_o};
  assign n202_o = {n166_o, n165_o, n164_o, n163_o};
  assign n203_o = {n162_o, n161_o, n160_o};
  assign n204_o = {n195_o, n196_o, n197_o, n198_o};
  assign n205_o = {n199_o, n200_o, n201_o, n202_o};
  assign n206_o = {n204_o, n205_o, n203_o};
  /* routers/synchronous/xbar.vhd:70:51  */
  assign n207_o = n159_o & n206_o;
  /* routers/synchronous/xbar.vhd:69:80  */
  assign n208_o = n157_o | n207_o;
  /* routers/synchronous/xbar.vhd:71:35  */
  assign n209_o = inPort[35:0];
  /* routers/synchronous/xbar.vhd:71:39  */
  assign n210_o = n209_o[35:1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n211_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n212_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n213_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n214_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n215_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n216_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n217_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n218_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n219_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n220_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n221_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n222_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n223_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n224_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n225_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n226_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n227_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n228_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n229_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n230_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n231_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n232_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n233_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n234_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n235_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n236_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n237_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n238_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n239_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n240_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n241_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n242_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n243_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n244_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n245_o = sel0[1];
  assign n246_o = {n245_o, n244_o, n243_o, n242_o};
  assign n247_o = {n241_o, n240_o, n239_o, n238_o};
  assign n248_o = {n237_o, n236_o, n235_o, n234_o};
  assign n249_o = {n233_o, n232_o, n231_o, n230_o};
  assign n250_o = {n229_o, n228_o, n227_o, n226_o};
  assign n251_o = {n225_o, n224_o, n223_o, n222_o};
  assign n252_o = {n221_o, n220_o, n219_o, n218_o};
  assign n253_o = {n217_o, n216_o, n215_o, n214_o};
  assign n254_o = {n213_o, n212_o, n211_o};
  assign n255_o = {n246_o, n247_o, n248_o, n249_o};
  assign n256_o = {n250_o, n251_o, n252_o, n253_o};
  assign n257_o = {n255_o, n256_o, n254_o};
  /* routers/synchronous/xbar.vhd:71:44  */
  assign n258_o = n210_o & n257_o;
  /* routers/synchronous/xbar.vhd:72:42  */
  assign n259_o = inPort[107:72];
  /* routers/synchronous/xbar.vhd:72:46  */
  assign n260_o = n259_o[35:1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n261_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n262_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n263_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n264_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n265_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n266_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n267_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n268_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n269_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n270_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n271_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n272_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n273_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n274_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n275_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n276_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n277_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n278_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n279_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n280_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n281_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n282_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n283_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n284_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n285_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n286_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n287_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n288_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n289_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n290_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n291_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n292_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n293_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n294_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n295_o = sel2[1];
  assign n296_o = {n295_o, n294_o, n293_o, n292_o};
  assign n297_o = {n291_o, n290_o, n289_o, n288_o};
  assign n298_o = {n287_o, n286_o, n285_o, n284_o};
  assign n299_o = {n283_o, n282_o, n281_o, n280_o};
  assign n300_o = {n279_o, n278_o, n277_o, n276_o};
  assign n301_o = {n275_o, n274_o, n273_o, n272_o};
  assign n302_o = {n271_o, n270_o, n269_o, n268_o};
  assign n303_o = {n267_o, n266_o, n265_o, n264_o};
  assign n304_o = {n263_o, n262_o, n261_o};
  assign n305_o = {n296_o, n297_o, n298_o, n299_o};
  assign n306_o = {n300_o, n301_o, n302_o, n303_o};
  assign n307_o = {n305_o, n306_o, n304_o};
  /* routers/synchronous/xbar.vhd:72:51  */
  assign n308_o = n260_o & n307_o;
  /* routers/synchronous/xbar.vhd:71:73  */
  assign n309_o = n258_o | n308_o;
  /* routers/synchronous/xbar.vhd:73:42  */
  assign n310_o = inPort[143:108];
  /* routers/synchronous/xbar.vhd:73:46  */
  assign n311_o = n310_o[35:1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n312_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n313_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n314_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n315_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n316_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n317_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n318_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n319_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n320_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n321_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n322_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n323_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n324_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n325_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n326_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n327_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n328_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n329_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n330_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n331_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n332_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n333_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n334_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n335_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n336_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n337_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n338_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n339_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n340_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n341_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n342_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n343_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n344_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n345_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n346_o = sel3[1];
  assign n347_o = {n346_o, n345_o, n344_o, n343_o};
  assign n348_o = {n342_o, n341_o, n340_o, n339_o};
  assign n349_o = {n338_o, n337_o, n336_o, n335_o};
  assign n350_o = {n334_o, n333_o, n332_o, n331_o};
  assign n351_o = {n330_o, n329_o, n328_o, n327_o};
  assign n352_o = {n326_o, n325_o, n324_o, n323_o};
  assign n353_o = {n322_o, n321_o, n320_o, n319_o};
  assign n354_o = {n318_o, n317_o, n316_o, n315_o};
  assign n355_o = {n314_o, n313_o, n312_o};
  assign n356_o = {n347_o, n348_o, n349_o, n350_o};
  assign n357_o = {n351_o, n352_o, n353_o, n354_o};
  assign n358_o = {n356_o, n357_o, n355_o};
  /* routers/synchronous/xbar.vhd:73:51  */
  assign n359_o = n311_o & n358_o;
  /* routers/synchronous/xbar.vhd:72:80  */
  assign n360_o = n309_o | n359_o;
  /* routers/synchronous/xbar.vhd:74:42  */
  assign n361_o = inPort[179:144];
  /* routers/synchronous/xbar.vhd:74:46  */
  assign n362_o = n361_o[35:1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n363_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n364_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n365_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n366_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n367_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n368_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n369_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n370_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n371_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n372_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n373_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n374_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n375_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n376_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n377_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n378_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n379_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n380_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n381_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n382_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n383_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n384_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n385_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n386_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n387_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n388_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n389_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n390_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n391_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n392_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n393_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n394_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n395_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n396_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n397_o = sel4[1];
  assign n398_o = {n397_o, n396_o, n395_o, n394_o};
  assign n399_o = {n393_o, n392_o, n391_o, n390_o};
  assign n400_o = {n389_o, n388_o, n387_o, n386_o};
  assign n401_o = {n385_o, n384_o, n383_o, n382_o};
  assign n402_o = {n381_o, n380_o, n379_o, n378_o};
  assign n403_o = {n377_o, n376_o, n375_o, n374_o};
  assign n404_o = {n373_o, n372_o, n371_o, n370_o};
  assign n405_o = {n369_o, n368_o, n367_o, n366_o};
  assign n406_o = {n365_o, n364_o, n363_o};
  assign n407_o = {n398_o, n399_o, n400_o, n401_o};
  assign n408_o = {n402_o, n403_o, n404_o, n405_o};
  assign n409_o = {n407_o, n408_o, n406_o};
  /* routers/synchronous/xbar.vhd:74:51  */
  assign n410_o = n362_o & n409_o;
  /* routers/synchronous/xbar.vhd:73:80  */
  assign n411_o = n360_o | n410_o;
  /* routers/synchronous/xbar.vhd:75:35  */
  assign n412_o = inPort[35:0];
  /* routers/synchronous/xbar.vhd:75:39  */
  assign n413_o = n412_o[35:1];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n414_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n415_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n416_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n417_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n418_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n419_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n420_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n421_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n422_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n423_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n424_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n425_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n426_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n427_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n428_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n429_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n430_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n431_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n432_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n433_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n434_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n435_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n436_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n437_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n438_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n439_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n440_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n441_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n442_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n443_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n444_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n445_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n446_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n447_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n448_o = sel0[2];
  assign n449_o = {n448_o, n447_o, n446_o, n445_o};
  assign n450_o = {n444_o, n443_o, n442_o, n441_o};
  assign n451_o = {n440_o, n439_o, n438_o, n437_o};
  assign n452_o = {n436_o, n435_o, n434_o, n433_o};
  assign n453_o = {n432_o, n431_o, n430_o, n429_o};
  assign n454_o = {n428_o, n427_o, n426_o, n425_o};
  assign n455_o = {n424_o, n423_o, n422_o, n421_o};
  assign n456_o = {n420_o, n419_o, n418_o, n417_o};
  assign n457_o = {n416_o, n415_o, n414_o};
  assign n458_o = {n449_o, n450_o, n451_o, n452_o};
  assign n459_o = {n453_o, n454_o, n455_o, n456_o};
  assign n460_o = {n458_o, n459_o, n457_o};
  /* routers/synchronous/xbar.vhd:75:44  */
  assign n461_o = n413_o & n460_o;
  /* routers/synchronous/xbar.vhd:76:42  */
  assign n462_o = inPort[71:36];
  /* routers/synchronous/xbar.vhd:76:46  */
  assign n463_o = n462_o[35:1];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n464_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n465_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n466_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n467_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n468_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n469_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n470_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n471_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n472_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n473_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n474_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n475_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n476_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n477_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n478_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n479_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n480_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n481_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n482_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n483_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n484_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n485_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n486_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n487_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n488_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n489_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n490_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n491_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n492_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n493_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n494_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n495_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n496_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n497_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n498_o = sel1[2];
  assign n499_o = {n498_o, n497_o, n496_o, n495_o};
  assign n500_o = {n494_o, n493_o, n492_o, n491_o};
  assign n501_o = {n490_o, n489_o, n488_o, n487_o};
  assign n502_o = {n486_o, n485_o, n484_o, n483_o};
  assign n503_o = {n482_o, n481_o, n480_o, n479_o};
  assign n504_o = {n478_o, n477_o, n476_o, n475_o};
  assign n505_o = {n474_o, n473_o, n472_o, n471_o};
  assign n506_o = {n470_o, n469_o, n468_o, n467_o};
  assign n507_o = {n466_o, n465_o, n464_o};
  assign n508_o = {n499_o, n500_o, n501_o, n502_o};
  assign n509_o = {n503_o, n504_o, n505_o, n506_o};
  assign n510_o = {n508_o, n509_o, n507_o};
  /* routers/synchronous/xbar.vhd:76:51  */
  assign n511_o = n463_o & n510_o;
  /* routers/synchronous/xbar.vhd:75:73  */
  assign n512_o = n461_o | n511_o;
  /* routers/synchronous/xbar.vhd:77:42  */
  assign n513_o = inPort[143:108];
  /* routers/synchronous/xbar.vhd:77:46  */
  assign n514_o = n513_o[35:1];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n515_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n516_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n517_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n518_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n519_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n520_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n521_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n522_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n523_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n524_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n525_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n526_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n527_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n528_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n529_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n530_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n531_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n532_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n533_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n534_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n535_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n536_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n537_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n538_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n539_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n540_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n541_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n542_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n543_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n544_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n545_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n546_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n547_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n548_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n549_o = sel3[2];
  assign n550_o = {n549_o, n548_o, n547_o, n546_o};
  assign n551_o = {n545_o, n544_o, n543_o, n542_o};
  assign n552_o = {n541_o, n540_o, n539_o, n538_o};
  assign n553_o = {n537_o, n536_o, n535_o, n534_o};
  assign n554_o = {n533_o, n532_o, n531_o, n530_o};
  assign n555_o = {n529_o, n528_o, n527_o, n526_o};
  assign n556_o = {n525_o, n524_o, n523_o, n522_o};
  assign n557_o = {n521_o, n520_o, n519_o, n518_o};
  assign n558_o = {n517_o, n516_o, n515_o};
  assign n559_o = {n550_o, n551_o, n552_o, n553_o};
  assign n560_o = {n554_o, n555_o, n556_o, n557_o};
  assign n561_o = {n559_o, n560_o, n558_o};
  /* routers/synchronous/xbar.vhd:77:51  */
  assign n562_o = n514_o & n561_o;
  /* routers/synchronous/xbar.vhd:76:80  */
  assign n563_o = n512_o | n562_o;
  /* routers/synchronous/xbar.vhd:78:42  */
  assign n564_o = inPort[179:144];
  /* routers/synchronous/xbar.vhd:78:46  */
  assign n565_o = n564_o[35:1];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n566_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n567_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n568_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n569_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n570_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n571_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n572_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n573_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n574_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n575_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n576_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n577_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n578_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n579_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n580_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n581_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n582_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n583_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n584_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n585_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n586_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n587_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n588_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n589_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n590_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n591_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n592_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n593_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n594_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n595_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n596_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n597_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n598_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n599_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n600_o = sel4[2];
  assign n601_o = {n600_o, n599_o, n598_o, n597_o};
  assign n602_o = {n596_o, n595_o, n594_o, n593_o};
  assign n603_o = {n592_o, n591_o, n590_o, n589_o};
  assign n604_o = {n588_o, n587_o, n586_o, n585_o};
  assign n605_o = {n584_o, n583_o, n582_o, n581_o};
  assign n606_o = {n580_o, n579_o, n578_o, n577_o};
  assign n607_o = {n576_o, n575_o, n574_o, n573_o};
  assign n608_o = {n572_o, n571_o, n570_o, n569_o};
  assign n609_o = {n568_o, n567_o, n566_o};
  assign n610_o = {n601_o, n602_o, n603_o, n604_o};
  assign n611_o = {n605_o, n606_o, n607_o, n608_o};
  assign n612_o = {n610_o, n611_o, n609_o};
  /* routers/synchronous/xbar.vhd:78:51  */
  assign n613_o = n565_o & n612_o;
  /* routers/synchronous/xbar.vhd:77:80  */
  assign n614_o = n563_o | n613_o;
  /* routers/synchronous/xbar.vhd:79:35  */
  assign n615_o = inPort[35:0];
  /* routers/synchronous/xbar.vhd:79:39  */
  assign n616_o = n615_o[35:1];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n617_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n618_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n619_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n620_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n621_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n622_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n623_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n624_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n625_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n626_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n627_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n628_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n629_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n630_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n631_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n632_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n633_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n634_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n635_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n636_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n637_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n638_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n639_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n640_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n641_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n642_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n643_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n644_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n645_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n646_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n647_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n648_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n649_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n650_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n651_o = sel0[3];
  assign n652_o = {n651_o, n650_o, n649_o, n648_o};
  assign n653_o = {n647_o, n646_o, n645_o, n644_o};
  assign n654_o = {n643_o, n642_o, n641_o, n640_o};
  assign n655_o = {n639_o, n638_o, n637_o, n636_o};
  assign n656_o = {n635_o, n634_o, n633_o, n632_o};
  assign n657_o = {n631_o, n630_o, n629_o, n628_o};
  assign n658_o = {n627_o, n626_o, n625_o, n624_o};
  assign n659_o = {n623_o, n622_o, n621_o, n620_o};
  assign n660_o = {n619_o, n618_o, n617_o};
  assign n661_o = {n652_o, n653_o, n654_o, n655_o};
  assign n662_o = {n656_o, n657_o, n658_o, n659_o};
  assign n663_o = {n661_o, n662_o, n660_o};
  /* routers/synchronous/xbar.vhd:79:44  */
  assign n664_o = n616_o & n663_o;
  /* routers/synchronous/xbar.vhd:80:42  */
  assign n665_o = inPort[71:36];
  /* routers/synchronous/xbar.vhd:80:46  */
  assign n666_o = n665_o[35:1];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n667_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n668_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n669_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n670_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n671_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n672_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n673_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n674_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n675_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n676_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n677_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n678_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n679_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n680_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n681_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n682_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n683_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n684_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n685_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n686_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n687_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n688_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n689_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n690_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n691_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n692_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n693_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n694_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n695_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n696_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n697_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n698_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n699_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n700_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n701_o = sel1[3];
  assign n702_o = {n701_o, n700_o, n699_o, n698_o};
  assign n703_o = {n697_o, n696_o, n695_o, n694_o};
  assign n704_o = {n693_o, n692_o, n691_o, n690_o};
  assign n705_o = {n689_o, n688_o, n687_o, n686_o};
  assign n706_o = {n685_o, n684_o, n683_o, n682_o};
  assign n707_o = {n681_o, n680_o, n679_o, n678_o};
  assign n708_o = {n677_o, n676_o, n675_o, n674_o};
  assign n709_o = {n673_o, n672_o, n671_o, n670_o};
  assign n710_o = {n669_o, n668_o, n667_o};
  assign n711_o = {n702_o, n703_o, n704_o, n705_o};
  assign n712_o = {n706_o, n707_o, n708_o, n709_o};
  assign n713_o = {n711_o, n712_o, n710_o};
  /* routers/synchronous/xbar.vhd:80:51  */
  assign n714_o = n666_o & n713_o;
  /* routers/synchronous/xbar.vhd:79:73  */
  assign n715_o = n664_o | n714_o;
  /* routers/synchronous/xbar.vhd:81:42  */
  assign n716_o = inPort[107:72];
  /* routers/synchronous/xbar.vhd:81:46  */
  assign n717_o = n716_o[35:1];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n718_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n719_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n720_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n721_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n722_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n723_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n724_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n725_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n726_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n727_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n728_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n729_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n730_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n731_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n732_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n733_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n734_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n735_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n736_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n737_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n738_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n739_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n740_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n741_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n742_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n743_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n744_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n745_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n746_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n747_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n748_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n749_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n750_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n751_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n752_o = sel2[3];
  assign n753_o = {n752_o, n751_o, n750_o, n749_o};
  assign n754_o = {n748_o, n747_o, n746_o, n745_o};
  assign n755_o = {n744_o, n743_o, n742_o, n741_o};
  assign n756_o = {n740_o, n739_o, n738_o, n737_o};
  assign n757_o = {n736_o, n735_o, n734_o, n733_o};
  assign n758_o = {n732_o, n731_o, n730_o, n729_o};
  assign n759_o = {n728_o, n727_o, n726_o, n725_o};
  assign n760_o = {n724_o, n723_o, n722_o, n721_o};
  assign n761_o = {n720_o, n719_o, n718_o};
  assign n762_o = {n753_o, n754_o, n755_o, n756_o};
  assign n763_o = {n757_o, n758_o, n759_o, n760_o};
  assign n764_o = {n762_o, n763_o, n761_o};
  /* routers/synchronous/xbar.vhd:81:51  */
  assign n765_o = n717_o & n764_o;
  /* routers/synchronous/xbar.vhd:80:80  */
  assign n766_o = n715_o | n765_o;
  /* routers/synchronous/xbar.vhd:82:42  */
  assign n767_o = inPort[179:144];
  /* routers/synchronous/xbar.vhd:82:46  */
  assign n768_o = n767_o[35:1];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n769_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n770_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n771_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n772_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n773_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n774_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n775_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n776_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n777_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n778_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n779_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n780_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n781_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n782_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n783_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n784_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n785_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n786_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n787_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n788_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n789_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n790_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n791_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n792_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n793_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n794_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n795_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n796_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n797_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n798_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n799_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n800_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n801_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n802_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n803_o = sel4[3];
  assign n804_o = {n803_o, n802_o, n801_o, n800_o};
  assign n805_o = {n799_o, n798_o, n797_o, n796_o};
  assign n806_o = {n795_o, n794_o, n793_o, n792_o};
  assign n807_o = {n791_o, n790_o, n789_o, n788_o};
  assign n808_o = {n787_o, n786_o, n785_o, n784_o};
  assign n809_o = {n783_o, n782_o, n781_o, n780_o};
  assign n810_o = {n779_o, n778_o, n777_o, n776_o};
  assign n811_o = {n775_o, n774_o, n773_o, n772_o};
  assign n812_o = {n771_o, n770_o, n769_o};
  assign n813_o = {n804_o, n805_o, n806_o, n807_o};
  assign n814_o = {n808_o, n809_o, n810_o, n811_o};
  assign n815_o = {n813_o, n814_o, n812_o};
  /* routers/synchronous/xbar.vhd:82:51  */
  assign n816_o = n768_o & n815_o;
  /* routers/synchronous/xbar.vhd:81:80  */
  assign n817_o = n766_o | n816_o;
  /* routers/synchronous/xbar.vhd:83:35  */
  assign n818_o = inPort[35:0];
  /* routers/synchronous/xbar.vhd:83:39  */
  assign n819_o = n818_o[35:1];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n820_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n821_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n822_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n823_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n824_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n825_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n826_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n827_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n828_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n829_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n830_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n831_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n832_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n833_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n834_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n835_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n836_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n837_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n838_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n839_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n840_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n841_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n842_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n843_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n844_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n845_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n846_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n847_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n848_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n849_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n850_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n851_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n852_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n853_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n854_o = sel0[0];
  assign n855_o = {n854_o, n853_o, n852_o, n851_o};
  assign n856_o = {n850_o, n849_o, n848_o, n847_o};
  assign n857_o = {n846_o, n845_o, n844_o, n843_o};
  assign n858_o = {n842_o, n841_o, n840_o, n839_o};
  assign n859_o = {n838_o, n837_o, n836_o, n835_o};
  assign n860_o = {n834_o, n833_o, n832_o, n831_o};
  assign n861_o = {n830_o, n829_o, n828_o, n827_o};
  assign n862_o = {n826_o, n825_o, n824_o, n823_o};
  assign n863_o = {n822_o, n821_o, n820_o};
  assign n864_o = {n855_o, n856_o, n857_o, n858_o};
  assign n865_o = {n859_o, n860_o, n861_o, n862_o};
  assign n866_o = {n864_o, n865_o, n863_o};
  /* routers/synchronous/xbar.vhd:83:44  */
  assign n867_o = n819_o & n866_o;
  /* routers/synchronous/xbar.vhd:84:42  */
  assign n868_o = inPort[71:36];
  /* routers/synchronous/xbar.vhd:84:46  */
  assign n869_o = n868_o[35:1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n870_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n871_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n872_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n873_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n874_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n875_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n876_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n877_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n878_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n879_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n880_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n881_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n882_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n883_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n884_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n885_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n886_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n887_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n888_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n889_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n890_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n891_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n892_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n893_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n894_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n895_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n896_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n897_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n898_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n899_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n900_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n901_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n902_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n903_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n904_o = sel1[1];
  assign n905_o = {n904_o, n903_o, n902_o, n901_o};
  assign n906_o = {n900_o, n899_o, n898_o, n897_o};
  assign n907_o = {n896_o, n895_o, n894_o, n893_o};
  assign n908_o = {n892_o, n891_o, n890_o, n889_o};
  assign n909_o = {n888_o, n887_o, n886_o, n885_o};
  assign n910_o = {n884_o, n883_o, n882_o, n881_o};
  assign n911_o = {n880_o, n879_o, n878_o, n877_o};
  assign n912_o = {n876_o, n875_o, n874_o, n873_o};
  assign n913_o = {n872_o, n871_o, n870_o};
  assign n914_o = {n905_o, n906_o, n907_o, n908_o};
  assign n915_o = {n909_o, n910_o, n911_o, n912_o};
  assign n916_o = {n914_o, n915_o, n913_o};
  /* routers/synchronous/xbar.vhd:84:51  */
  assign n917_o = n869_o & n916_o;
  /* routers/synchronous/xbar.vhd:83:73  */
  assign n918_o = n867_o | n917_o;
  /* routers/synchronous/xbar.vhd:85:42  */
  assign n919_o = inPort[107:72];
  /* routers/synchronous/xbar.vhd:85:46  */
  assign n920_o = n919_o[35:1];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n921_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n922_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n923_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n924_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n925_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n926_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n927_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n928_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n929_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n930_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n931_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n932_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n933_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n934_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n935_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n936_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n937_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n938_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n939_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n940_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n941_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n942_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n943_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n944_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n945_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n946_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n947_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n948_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n949_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n950_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n951_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n952_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n953_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n954_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n955_o = sel2[2];
  assign n956_o = {n955_o, n954_o, n953_o, n952_o};
  assign n957_o = {n951_o, n950_o, n949_o, n948_o};
  assign n958_o = {n947_o, n946_o, n945_o, n944_o};
  assign n959_o = {n943_o, n942_o, n941_o, n940_o};
  assign n960_o = {n939_o, n938_o, n937_o, n936_o};
  assign n961_o = {n935_o, n934_o, n933_o, n932_o};
  assign n962_o = {n931_o, n930_o, n929_o, n928_o};
  assign n963_o = {n927_o, n926_o, n925_o, n924_o};
  assign n964_o = {n923_o, n922_o, n921_o};
  assign n965_o = {n956_o, n957_o, n958_o, n959_o};
  assign n966_o = {n960_o, n961_o, n962_o, n963_o};
  assign n967_o = {n965_o, n966_o, n964_o};
  /* routers/synchronous/xbar.vhd:85:51  */
  assign n968_o = n920_o & n967_o;
  /* routers/synchronous/xbar.vhd:84:80  */
  assign n969_o = n918_o | n968_o;
  /* routers/synchronous/xbar.vhd:86:42  */
  assign n970_o = inPort[143:108];
  /* routers/synchronous/xbar.vhd:86:46  */
  assign n971_o = n970_o[35:1];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n972_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n973_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n974_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n975_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n976_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n977_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n978_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n979_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n980_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n981_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n982_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n983_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n984_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n985_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n986_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n987_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n988_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n989_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n990_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n991_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n992_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n993_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n994_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n995_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n996_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n997_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n998_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n999_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n1000_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n1001_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n1002_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n1003_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n1004_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n1005_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n1006_o = sel3[3];
  assign n1007_o = {n1006_o, n1005_o, n1004_o, n1003_o};
  assign n1008_o = {n1002_o, n1001_o, n1000_o, n999_o};
  assign n1009_o = {n998_o, n997_o, n996_o, n995_o};
  assign n1010_o = {n994_o, n993_o, n992_o, n991_o};
  assign n1011_o = {n990_o, n989_o, n988_o, n987_o};
  assign n1012_o = {n986_o, n985_o, n984_o, n983_o};
  assign n1013_o = {n982_o, n981_o, n980_o, n979_o};
  assign n1014_o = {n978_o, n977_o, n976_o, n975_o};
  assign n1015_o = {n974_o, n973_o, n972_o};
  assign n1016_o = {n1007_o, n1008_o, n1009_o, n1010_o};
  assign n1017_o = {n1011_o, n1012_o, n1013_o, n1014_o};
  assign n1018_o = {n1016_o, n1017_o, n1015_o};
  /* routers/synchronous/xbar.vhd:86:51  */
  assign n1019_o = n971_o & n1018_o;
  /* routers/synchronous/xbar.vhd:85:80  */
  assign n1020_o = n969_o | n1019_o;
  assign n1026_o = {n1020_o, 1'bZ, n817_o, 1'bZ, n614_o, 1'bZ, n411_o, 1'bZ, n208_o, 1'bZ};
endmodule

