
module counter_WIDTH3_0 ( clk, reset, enable, cnt );
  output [2:0] cnt;
  input clk, reset, enable;
  wire   n6, n7, n10, n11, n13, n1, n2, n3, n4;

  HS65_LS_DFPRQX9 \reg_reg[0]  ( .D(n13), .CP(clk), .RN(n1), .Q(cnt[0]) );
  HS65_LS_DFPRQX9 \reg_reg[2]  ( .D(n11), .CP(clk), .RN(n1), .Q(cnt[2]) );
  HS65_LS_DFPRQX9 \reg_reg[1]  ( .D(n10), .CP(clk), .RN(n1), .Q(cnt[1]) );
  HS65_LH_OAI22X1 U3 ( .A(enable), .B(n2), .C(cnt[0]), .D(n6), .Z(n13) );
  HS65_LH_OA12X4 U4 ( .A(cnt[0]), .B(cnt[2]), .C(enable), .Z(n7) );
  HS65_LH_NAND2X2 U5 ( .A(enable), .B(n3), .Z(n6) );
  HS65_LH_OAI32X2 U6 ( .A(n4), .B(n6), .C(n2), .D(enable), .E(n3), .Z(n11) );
  HS65_LS_IVX9 U7 ( .A(reset), .Z(n1) );
  HS65_LS_OAI32X5 U8 ( .A(n2), .B(cnt[1]), .C(n6), .D(n7), .E(n4), .Z(n10) );
  HS65_LS_IVX9 U9 ( .A(cnt[0]), .Z(n2) );
  HS65_LS_IVX9 U10 ( .A(cnt[1]), .Z(n4) );
  HS65_LS_IVX9 U11 ( .A(cnt[2]), .Z(n3) );
endmodule


module bram_DATA16_ADDR2_0 ( clk, reset, rd_addr, wr_addr, wr_data, wr_ena, 
        rd_data );
  input [1:0] rd_addr;
  input [1:0] wr_addr;
  input [15:0] wr_data;
  output [15:0] rd_data;
  input clk, reset, wr_ena;
  wire   \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] ,
         \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][15] , \mem[1][14] , \mem[1][13] ,
         \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] , \mem[1][8] ,
         \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] ,
         \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][15] , \mem[0][14] ,
         \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] ,
         \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] ,
         \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n1, n2, n3, n4, n5, n6, n7, n8, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90;

  HS65_LS_DFPRQX9 \mem_reg[3][15]  ( .D(n80), .CP(clk), .RN(n1), .Q(
        \mem[3][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][14]  ( .D(n79), .CP(clk), .RN(n1), .Q(
        \mem[3][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][13]  ( .D(n78), .CP(clk), .RN(n1), .Q(
        \mem[3][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][12]  ( .D(n77), .CP(clk), .RN(n1), .Q(
        \mem[3][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][11]  ( .D(n76), .CP(clk), .RN(n1), .Q(
        \mem[3][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][10]  ( .D(n75), .CP(clk), .RN(n1), .Q(
        \mem[3][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][9]  ( .D(n74), .CP(clk), .RN(n1), .Q(\mem[3][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][8]  ( .D(n73), .CP(clk), .RN(n1), .Q(\mem[3][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][7]  ( .D(n72), .CP(clk), .RN(n1), .Q(\mem[3][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][6]  ( .D(n71), .CP(clk), .RN(n1), .Q(\mem[3][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][5]  ( .D(n70), .CP(clk), .RN(n1), .Q(\mem[3][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][4]  ( .D(n69), .CP(clk), .RN(n1), .Q(\mem[3][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][3]  ( .D(n68), .CP(clk), .RN(n1), .Q(\mem[3][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][2]  ( .D(n67), .CP(clk), .RN(n2), .Q(\mem[3][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][1]  ( .D(n66), .CP(clk), .RN(n2), .Q(\mem[3][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][0]  ( .D(n65), .CP(clk), .RN(n2), .Q(\mem[3][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][15]  ( .D(n64), .CP(clk), .RN(n2), .Q(
        \mem[2][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][14]  ( .D(n63), .CP(clk), .RN(n2), .Q(
        \mem[2][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][13]  ( .D(n62), .CP(clk), .RN(n2), .Q(
        \mem[2][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][12]  ( .D(n61), .CP(clk), .RN(n2), .Q(
        \mem[2][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][11]  ( .D(n60), .CP(clk), .RN(n2), .Q(
        \mem[2][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][10]  ( .D(n59), .CP(clk), .RN(n2), .Q(
        \mem[2][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][9]  ( .D(n58), .CP(clk), .RN(n2), .Q(\mem[2][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][8]  ( .D(n57), .CP(clk), .RN(n2), .Q(\mem[2][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][7]  ( .D(n56), .CP(clk), .RN(n2), .Q(\mem[2][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][6]  ( .D(n55), .CP(clk), .RN(n2), .Q(\mem[2][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][5]  ( .D(n54), .CP(clk), .RN(n3), .Q(\mem[2][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][4]  ( .D(n53), .CP(clk), .RN(n3), .Q(\mem[2][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][3]  ( .D(n52), .CP(clk), .RN(n3), .Q(\mem[2][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][2]  ( .D(n51), .CP(clk), .RN(n3), .Q(\mem[2][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][1]  ( .D(n50), .CP(clk), .RN(n3), .Q(\mem[2][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][0]  ( .D(n49), .CP(clk), .RN(n3), .Q(\mem[2][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][15]  ( .D(n48), .CP(clk), .RN(n3), .Q(
        \mem[1][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][14]  ( .D(n47), .CP(clk), .RN(n3), .Q(
        \mem[1][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][13]  ( .D(n46), .CP(clk), .RN(n3), .Q(
        \mem[1][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][12]  ( .D(n45), .CP(clk), .RN(n3), .Q(
        \mem[1][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][11]  ( .D(n44), .CP(clk), .RN(n3), .Q(
        \mem[1][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][10]  ( .D(n43), .CP(clk), .RN(n3), .Q(
        \mem[1][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][9]  ( .D(n42), .CP(clk), .RN(n3), .Q(\mem[1][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][8]  ( .D(n41), .CP(clk), .RN(n4), .Q(\mem[1][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][7]  ( .D(n40), .CP(clk), .RN(n4), .Q(\mem[1][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][6]  ( .D(n39), .CP(clk), .RN(n4), .Q(\mem[1][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][5]  ( .D(n38), .CP(clk), .RN(n4), .Q(\mem[1][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][4]  ( .D(n37), .CP(clk), .RN(n4), .Q(\mem[1][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][3]  ( .D(n36), .CP(clk), .RN(n4), .Q(\mem[1][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][2]  ( .D(n35), .CP(clk), .RN(n4), .Q(\mem[1][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][1]  ( .D(n34), .CP(clk), .RN(n4), .Q(\mem[1][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][0]  ( .D(n33), .CP(clk), .RN(n4), .Q(\mem[1][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][15]  ( .D(n32), .CP(clk), .RN(n4), .Q(
        \mem[0][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][14]  ( .D(n31), .CP(clk), .RN(n4), .Q(
        \mem[0][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][13]  ( .D(n30), .CP(clk), .RN(n4), .Q(
        \mem[0][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][12]  ( .D(n29), .CP(clk), .RN(n4), .Q(
        \mem[0][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][11]  ( .D(n28), .CP(clk), .RN(n5), .Q(
        \mem[0][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][10]  ( .D(n27), .CP(clk), .RN(n5), .Q(
        \mem[0][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][9]  ( .D(n26), .CP(clk), .RN(n5), .Q(\mem[0][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][8]  ( .D(n25), .CP(clk), .RN(n5), .Q(\mem[0][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][7]  ( .D(n24), .CP(clk), .RN(n5), .Q(\mem[0][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][6]  ( .D(n23), .CP(clk), .RN(n5), .Q(\mem[0][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][5]  ( .D(n22), .CP(clk), .RN(n5), .Q(\mem[0][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][4]  ( .D(n21), .CP(clk), .RN(n5), .Q(\mem[0][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][3]  ( .D(n20), .CP(clk), .RN(n5), .Q(\mem[0][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][2]  ( .D(n19), .CP(clk), .RN(n5), .Q(\mem[0][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][1]  ( .D(n18), .CP(clk), .RN(n5), .Q(\mem[0][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][0]  ( .D(n17), .CP(clk), .RN(n5), .Q(\mem[0][0] ) );
  HS65_LS_DFPRQX9 \rd_data_reg[15]  ( .D(N17), .CP(clk), .RN(n5), .Q(
        rd_data[15]) );
  HS65_LS_DFPRQX9 \rd_data_reg[14]  ( .D(N18), .CP(clk), .RN(n6), .Q(
        rd_data[14]) );
  HS65_LS_DFPRQX9 \rd_data_reg[13]  ( .D(N19), .CP(clk), .RN(n6), .Q(
        rd_data[13]) );
  HS65_LS_DFPRQX9 \rd_data_reg[12]  ( .D(N20), .CP(clk), .RN(n6), .Q(
        rd_data[12]) );
  HS65_LS_DFPRQX9 \rd_data_reg[11]  ( .D(N21), .CP(clk), .RN(n6), .Q(
        rd_data[11]) );
  HS65_LS_DFPRQX9 \rd_data_reg[10]  ( .D(N22), .CP(clk), .RN(n6), .Q(
        rd_data[10]) );
  HS65_LS_DFPRQX9 \rd_data_reg[9]  ( .D(N23), .CP(clk), .RN(n6), .Q(rd_data[9]) );
  HS65_LS_DFPRQX9 \rd_data_reg[8]  ( .D(N24), .CP(clk), .RN(n6), .Q(rd_data[8]) );
  HS65_LS_DFPRQX9 \rd_data_reg[7]  ( .D(N25), .CP(clk), .RN(n6), .Q(rd_data[7]) );
  HS65_LS_DFPRQX9 \rd_data_reg[6]  ( .D(N26), .CP(clk), .RN(n6), .Q(rd_data[6]) );
  HS65_LS_DFPRQX9 \rd_data_reg[5]  ( .D(N27), .CP(clk), .RN(n6), .Q(rd_data[5]) );
  HS65_LS_DFPRQX9 \rd_data_reg[4]  ( .D(N28), .CP(clk), .RN(n6), .Q(rd_data[4]) );
  HS65_LS_DFPRQX9 \rd_data_reg[3]  ( .D(N29), .CP(clk), .RN(n6), .Q(rd_data[3]) );
  HS65_LS_DFPRQX9 \rd_data_reg[2]  ( .D(N30), .CP(clk), .RN(n6), .Q(rd_data[2]) );
  HS65_LS_DFPRQX9 \rd_data_reg[1]  ( .D(N31), .CP(clk), .RN(n7), .Q(rd_data[1]) );
  HS65_LS_DFPRQX9 \rd_data_reg[0]  ( .D(N32), .CP(clk), .RN(n7), .Q(rd_data[0]) );
  HS65_LS_BFX9 U3 ( .A(n81), .Z(n4) );
  HS65_LS_BFX9 U4 ( .A(n81), .Z(n3) );
  HS65_LS_BFX9 U5 ( .A(n81), .Z(n2) );
  HS65_LS_BFX9 U6 ( .A(n83), .Z(n81) );
  HS65_LS_BFX9 U7 ( .A(n8), .Z(n6) );
  HS65_LS_BFX9 U8 ( .A(n8), .Z(n5) );
  HS65_LS_BFX9 U9 ( .A(n82), .Z(n1) );
  HS65_LS_BFX9 U10 ( .A(n83), .Z(n82) );
  HS65_LS_BFX9 U11 ( .A(n8), .Z(n7) );
  HS65_LS_BFX9 U12 ( .A(n83), .Z(n8) );
  HS65_LS_IVX9 U13 ( .A(reset), .Z(n83) );
  HS65_LS_IVX9 U14 ( .A(n10), .Z(n86) );
  HS65_LS_IVX9 U15 ( .A(n9), .Z(n87) );
  HS65_LS_NAND3X5 U16 ( .A(wr_ena), .B(n88), .C(wr_addr[0]), .Z(n10) );
  HS65_LS_IVX9 U17 ( .A(wr_addr[0]), .Z(n89) );
  HS65_LS_NAND3X5 U18 ( .A(n89), .B(n88), .C(wr_ena), .Z(n9) );
  HS65_LS_IVX9 U19 ( .A(n11), .Z(n85) );
  HS65_LS_IVX9 U20 ( .A(n12), .Z(n84) );
  HS65_LS_NAND3X5 U21 ( .A(wr_ena), .B(n89), .C(wr_addr[1]), .Z(n11) );
  HS65_LS_NOR2X6 U22 ( .A(n90), .B(rd_addr[1]), .Z(n14) );
  HS65_LS_NOR2X6 U23 ( .A(rd_addr[0]), .B(rd_addr[1]), .Z(n13) );
  HS65_LS_IVX9 U24 ( .A(wr_addr[1]), .Z(n88) );
  HS65_LS_NAND3X5 U25 ( .A(wr_addr[0]), .B(wr_ena), .C(wr_addr[1]), .Z(n12) );
  HS65_LS_AND2X4 U26 ( .A(rd_addr[1]), .B(n90), .Z(n15) );
  HS65_LH_AND2X4 U27 ( .A(rd_addr[1]), .B(rd_addr[0]), .Z(n16) );
  HS65_LS_IVX9 U28 ( .A(rd_addr[0]), .Z(n90) );
  HS65_LS_MX41X7 U29 ( .D0(n13), .S0(\mem[0][0] ), .D1(n14), .S1(\mem[1][0] ), 
        .D2(n15), .S2(\mem[2][0] ), .D3(n16), .S3(\mem[3][0] ), .Z(N32) );
  HS65_LS_MX41X7 U30 ( .D0(n13), .S0(\mem[0][1] ), .D1(n14), .S1(\mem[1][1] ), 
        .D2(n15), .S2(\mem[2][1] ), .D3(n16), .S3(\mem[3][1] ), .Z(N31) );
  HS65_LS_MX41X7 U31 ( .D0(n13), .S0(\mem[0][2] ), .D1(n14), .S1(\mem[1][2] ), 
        .D2(n15), .S2(\mem[2][2] ), .D3(n16), .S3(\mem[3][2] ), .Z(N30) );
  HS65_LS_MX41X7 U32 ( .D0(n13), .S0(\mem[0][3] ), .D1(n14), .S1(\mem[1][3] ), 
        .D2(n15), .S2(\mem[2][3] ), .D3(n16), .S3(\mem[3][3] ), .Z(N29) );
  HS65_LS_MX41X7 U33 ( .D0(n13), .S0(\mem[0][4] ), .D1(n14), .S1(\mem[1][4] ), 
        .D2(n15), .S2(\mem[2][4] ), .D3(n16), .S3(\mem[3][4] ), .Z(N28) );
  HS65_LS_MX41X7 U34 ( .D0(n13), .S0(\mem[0][5] ), .D1(n14), .S1(\mem[1][5] ), 
        .D2(n15), .S2(\mem[2][5] ), .D3(n16), .S3(\mem[3][5] ), .Z(N27) );
  HS65_LS_MX41X7 U35 ( .D0(n13), .S0(\mem[0][6] ), .D1(n14), .S1(\mem[1][6] ), 
        .D2(n15), .S2(\mem[2][6] ), .D3(n16), .S3(\mem[3][6] ), .Z(N26) );
  HS65_LS_MX41X7 U36 ( .D0(n13), .S0(\mem[0][7] ), .D1(n14), .S1(\mem[1][7] ), 
        .D2(n15), .S2(\mem[2][7] ), .D3(n16), .S3(\mem[3][7] ), .Z(N25) );
  HS65_LS_MX41X7 U37 ( .D0(n13), .S0(\mem[0][8] ), .D1(n14), .S1(\mem[1][8] ), 
        .D2(n15), .S2(\mem[2][8] ), .D3(n16), .S3(\mem[3][8] ), .Z(N24) );
  HS65_LS_MX41X7 U38 ( .D0(n13), .S0(\mem[0][9] ), .D1(n14), .S1(\mem[1][9] ), 
        .D2(n15), .S2(\mem[2][9] ), .D3(n16), .S3(\mem[3][9] ), .Z(N23) );
  HS65_LS_MX41X7 U39 ( .D0(n13), .S0(\mem[0][10] ), .D1(n14), .S1(\mem[1][10] ), .D2(n15), .S2(\mem[2][10] ), .D3(n16), .S3(\mem[3][10] ), .Z(N22) );
  HS65_LS_MX41X7 U40 ( .D0(n13), .S0(\mem[0][11] ), .D1(n14), .S1(\mem[1][11] ), .D2(n15), .S2(\mem[2][11] ), .D3(n16), .S3(\mem[3][11] ), .Z(N21) );
  HS65_LS_MX41X7 U41 ( .D0(n13), .S0(\mem[0][12] ), .D1(n14), .S1(\mem[1][12] ), .D2(n15), .S2(\mem[2][12] ), .D3(n16), .S3(\mem[3][12] ), .Z(N20) );
  HS65_LS_MX41X7 U42 ( .D0(n13), .S0(\mem[0][13] ), .D1(n14), .S1(\mem[1][13] ), .D2(n15), .S2(\mem[2][13] ), .D3(n16), .S3(\mem[3][13] ), .Z(N19) );
  HS65_LS_MX41X7 U43 ( .D0(n13), .S0(\mem[0][14] ), .D1(n14), .S1(\mem[1][14] ), .D2(n15), .S2(\mem[2][14] ), .D3(n16), .S3(\mem[3][14] ), .Z(N18) );
  HS65_LS_MX41X7 U44 ( .D0(n13), .S0(\mem[0][15] ), .D1(n14), .S1(\mem[1][15] ), .D2(n15), .S2(\mem[2][15] ), .D3(n16), .S3(\mem[3][15] ), .Z(N17) );
  HS65_LS_AO22X9 U45 ( .A(wr_data[0]), .B(n86), .C(n10), .D(\mem[1][0] ), .Z(
        n33) );
  HS65_LS_AO22X9 U46 ( .A(wr_data[1]), .B(n86), .C(n10), .D(\mem[1][1] ), .Z(
        n34) );
  HS65_LS_AO22X9 U47 ( .A(wr_data[2]), .B(n86), .C(n10), .D(\mem[1][2] ), .Z(
        n35) );
  HS65_LS_AO22X9 U48 ( .A(wr_data[3]), .B(n86), .C(n10), .D(\mem[1][3] ), .Z(
        n36) );
  HS65_LS_AO22X9 U49 ( .A(wr_data[4]), .B(n86), .C(n10), .D(\mem[1][4] ), .Z(
        n37) );
  HS65_LS_AO22X9 U50 ( .A(wr_data[5]), .B(n86), .C(n10), .D(\mem[1][5] ), .Z(
        n38) );
  HS65_LS_AO22X9 U51 ( .A(wr_data[6]), .B(n86), .C(n10), .D(\mem[1][6] ), .Z(
        n39) );
  HS65_LS_AO22X9 U52 ( .A(wr_data[7]), .B(n86), .C(n10), .D(\mem[1][7] ), .Z(
        n40) );
  HS65_LS_AO22X9 U53 ( .A(wr_data[8]), .B(n86), .C(n10), .D(\mem[1][8] ), .Z(
        n41) );
  HS65_LS_AO22X9 U54 ( .A(wr_data[9]), .B(n86), .C(n10), .D(\mem[1][9] ), .Z(
        n42) );
  HS65_LS_AO22X9 U55 ( .A(wr_data[10]), .B(n86), .C(n10), .D(\mem[1][10] ), 
        .Z(n43) );
  HS65_LS_AO22X9 U56 ( .A(wr_data[11]), .B(n86), .C(n10), .D(\mem[1][11] ), 
        .Z(n44) );
  HS65_LS_AO22X9 U57 ( .A(wr_data[12]), .B(n86), .C(n10), .D(\mem[1][12] ), 
        .Z(n45) );
  HS65_LS_AO22X9 U58 ( .A(wr_data[13]), .B(n86), .C(n10), .D(\mem[1][13] ), 
        .Z(n46) );
  HS65_LS_AO22X9 U59 ( .A(wr_data[14]), .B(n86), .C(n10), .D(\mem[1][14] ), 
        .Z(n47) );
  HS65_LS_AO22X9 U60 ( .A(wr_data[15]), .B(n86), .C(n10), .D(\mem[1][15] ), 
        .Z(n48) );
  HS65_LS_AO22X9 U61 ( .A(wr_data[0]), .B(n85), .C(n11), .D(\mem[2][0] ), .Z(
        n49) );
  HS65_LS_AO22X9 U62 ( .A(wr_data[1]), .B(n85), .C(n11), .D(\mem[2][1] ), .Z(
        n50) );
  HS65_LS_AO22X9 U63 ( .A(wr_data[2]), .B(n85), .C(n11), .D(\mem[2][2] ), .Z(
        n51) );
  HS65_LS_AO22X9 U64 ( .A(wr_data[3]), .B(n85), .C(n11), .D(\mem[2][3] ), .Z(
        n52) );
  HS65_LS_AO22X9 U65 ( .A(wr_data[4]), .B(n85), .C(n11), .D(\mem[2][4] ), .Z(
        n53) );
  HS65_LS_AO22X9 U66 ( .A(wr_data[5]), .B(n85), .C(n11), .D(\mem[2][5] ), .Z(
        n54) );
  HS65_LS_AO22X9 U67 ( .A(wr_data[6]), .B(n85), .C(n11), .D(\mem[2][6] ), .Z(
        n55) );
  HS65_LS_AO22X9 U68 ( .A(wr_data[7]), .B(n85), .C(n11), .D(\mem[2][7] ), .Z(
        n56) );
  HS65_LS_AO22X9 U69 ( .A(wr_data[8]), .B(n85), .C(n11), .D(\mem[2][8] ), .Z(
        n57) );
  HS65_LS_AO22X9 U70 ( .A(wr_data[9]), .B(n85), .C(n11), .D(\mem[2][9] ), .Z(
        n58) );
  HS65_LS_AO22X9 U71 ( .A(wr_data[10]), .B(n85), .C(n11), .D(\mem[2][10] ), 
        .Z(n59) );
  HS65_LS_AO22X9 U72 ( .A(wr_data[11]), .B(n85), .C(n11), .D(\mem[2][11] ), 
        .Z(n60) );
  HS65_LS_AO22X9 U73 ( .A(wr_data[12]), .B(n85), .C(n11), .D(\mem[2][12] ), 
        .Z(n61) );
  HS65_LS_AO22X9 U74 ( .A(wr_data[13]), .B(n85), .C(n11), .D(\mem[2][13] ), 
        .Z(n62) );
  HS65_LS_AO22X9 U75 ( .A(wr_data[14]), .B(n85), .C(n11), .D(\mem[2][14] ), 
        .Z(n63) );
  HS65_LS_AO22X9 U76 ( .A(wr_data[15]), .B(n85), .C(n11), .D(\mem[2][15] ), 
        .Z(n64) );
  HS65_LS_AO22X9 U77 ( .A(n87), .B(wr_data[0]), .C(n9), .D(\mem[0][0] ), .Z(
        n17) );
  HS65_LS_AO22X9 U78 ( .A(n87), .B(wr_data[1]), .C(n9), .D(\mem[0][1] ), .Z(
        n18) );
  HS65_LS_AO22X9 U79 ( .A(n87), .B(wr_data[2]), .C(n9), .D(\mem[0][2] ), .Z(
        n19) );
  HS65_LS_AO22X9 U80 ( .A(n87), .B(wr_data[3]), .C(n9), .D(\mem[0][3] ), .Z(
        n20) );
  HS65_LS_AO22X9 U81 ( .A(n87), .B(wr_data[4]), .C(n9), .D(\mem[0][4] ), .Z(
        n21) );
  HS65_LS_AO22X9 U82 ( .A(n87), .B(wr_data[5]), .C(n9), .D(\mem[0][5] ), .Z(
        n22) );
  HS65_LS_AO22X9 U83 ( .A(n87), .B(wr_data[6]), .C(n9), .D(\mem[0][6] ), .Z(
        n23) );
  HS65_LS_AO22X9 U84 ( .A(n87), .B(wr_data[7]), .C(n9), .D(\mem[0][7] ), .Z(
        n24) );
  HS65_LS_AO22X9 U85 ( .A(n87), .B(wr_data[8]), .C(n9), .D(\mem[0][8] ), .Z(
        n25) );
  HS65_LS_AO22X9 U86 ( .A(n87), .B(wr_data[9]), .C(n9), .D(\mem[0][9] ), .Z(
        n26) );
  HS65_LS_AO22X9 U87 ( .A(n87), .B(wr_data[10]), .C(n9), .D(\mem[0][10] ), .Z(
        n27) );
  HS65_LS_AO22X9 U88 ( .A(n87), .B(wr_data[11]), .C(n9), .D(\mem[0][11] ), .Z(
        n28) );
  HS65_LS_AO22X9 U89 ( .A(n87), .B(wr_data[12]), .C(n9), .D(\mem[0][12] ), .Z(
        n29) );
  HS65_LS_AO22X9 U90 ( .A(n87), .B(wr_data[13]), .C(n9), .D(\mem[0][13] ), .Z(
        n30) );
  HS65_LS_AO22X9 U91 ( .A(n87), .B(wr_data[14]), .C(n9), .D(\mem[0][14] ), .Z(
        n31) );
  HS65_LS_AO22X9 U92 ( .A(n87), .B(wr_data[15]), .C(n9), .D(\mem[0][15] ), .Z(
        n32) );
  HS65_LS_AO22X9 U93 ( .A(wr_data[0]), .B(n84), .C(n12), .D(\mem[3][0] ), .Z(
        n65) );
  HS65_LS_AO22X9 U94 ( .A(wr_data[1]), .B(n84), .C(n12), .D(\mem[3][1] ), .Z(
        n66) );
  HS65_LS_AO22X9 U95 ( .A(wr_data[2]), .B(n84), .C(n12), .D(\mem[3][2] ), .Z(
        n67) );
  HS65_LS_AO22X9 U96 ( .A(wr_data[3]), .B(n84), .C(n12), .D(\mem[3][3] ), .Z(
        n68) );
  HS65_LS_AO22X9 U97 ( .A(wr_data[4]), .B(n84), .C(n12), .D(\mem[3][4] ), .Z(
        n69) );
  HS65_LS_AO22X9 U98 ( .A(wr_data[5]), .B(n84), .C(n12), .D(\mem[3][5] ), .Z(
        n70) );
  HS65_LS_AO22X9 U99 ( .A(wr_data[6]), .B(n84), .C(n12), .D(\mem[3][6] ), .Z(
        n71) );
  HS65_LS_AO22X9 U100 ( .A(wr_data[7]), .B(n84), .C(n12), .D(\mem[3][7] ), .Z(
        n72) );
  HS65_LS_AO22X9 U101 ( .A(wr_data[8]), .B(n84), .C(n12), .D(\mem[3][8] ), .Z(
        n73) );
  HS65_LS_AO22X9 U102 ( .A(wr_data[9]), .B(n84), .C(n12), .D(\mem[3][9] ), .Z(
        n74) );
  HS65_LS_AO22X9 U103 ( .A(wr_data[10]), .B(n84), .C(n12), .D(\mem[3][10] ), 
        .Z(n75) );
  HS65_LS_AO22X9 U104 ( .A(wr_data[11]), .B(n84), .C(n12), .D(\mem[3][11] ), 
        .Z(n76) );
  HS65_LS_AO22X9 U105 ( .A(wr_data[12]), .B(n84), .C(n12), .D(\mem[3][12] ), 
        .Z(n77) );
  HS65_LS_AO22X9 U106 ( .A(wr_data[13]), .B(n84), .C(n12), .D(\mem[3][13] ), 
        .Z(n78) );
  HS65_LS_AO22X9 U107 ( .A(wr_data[14]), .B(n84), .C(n12), .D(\mem[3][14] ), 
        .Z(n79) );
  HS65_LS_AO22X9 U108 ( .A(wr_data[15]), .B(n84), .C(n12), .D(\mem[3][15] ), 
        .Z(n80) );
endmodule


module bram_DATA32_ADDR2_0 ( clk, reset, rd_addr, wr_addr, wr_data, wr_ena, 
        rd_data );
  input [1:0] rd_addr;
  input [1:0] wr_addr;
  input [31:0] wr_data;
  output [31:0] rd_data;
  input clk, reset, wr_ena;
  wire   \mem[3][31] , \mem[3][30] , \mem[3][29] , \mem[3][28] , \mem[3][27] ,
         \mem[3][26] , \mem[3][25] , \mem[3][24] , \mem[3][23] , \mem[3][22] ,
         \mem[3][21] , \mem[3][20] , \mem[3][19] , \mem[3][18] , \mem[3][17] ,
         \mem[3][16] , \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] ,
         \mem[3][11] , \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] ,
         \mem[3][6] , \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] ,
         \mem[3][1] , \mem[3][0] , \mem[2][31] , \mem[2][30] , \mem[2][29] ,
         \mem[2][28] , \mem[2][27] , \mem[2][26] , \mem[2][25] , \mem[2][24] ,
         \mem[2][23] , \mem[2][22] , \mem[2][21] , \mem[2][20] , \mem[2][19] ,
         \mem[2][18] , \mem[2][17] , \mem[2][16] , \mem[2][15] , \mem[2][14] ,
         \mem[2][13] , \mem[2][12] , \mem[2][11] , \mem[2][10] , \mem[2][9] ,
         \mem[2][8] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][31] ,
         \mem[1][30] , \mem[1][29] , \mem[1][28] , \mem[1][27] , \mem[1][26] ,
         \mem[1][25] , \mem[1][24] , \mem[1][23] , \mem[1][22] , \mem[1][21] ,
         \mem[1][20] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][31] , \mem[0][30] , \mem[0][29] , \mem[0][28] ,
         \mem[0][27] , \mem[0][26] , \mem[0][25] , \mem[0][24] , \mem[0][23] ,
         \mem[0][22] , \mem[0][21] , \mem[0][20] , \mem[0][19] , \mem[0][18] ,
         \mem[0][17] , \mem[0][16] , \mem[0][15] , \mem[0][14] , \mem[0][13] ,
         \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] , \mem[0][8] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N17, N18, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36,
         N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n1, n2, n3, n4, n5, n6, n7, n8, n9, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192;

  HS65_LS_DFPRQX9 \mem_reg[3][31]  ( .D(n144), .CP(clk), .RN(n171), .Q(
        \mem[3][31] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][30]  ( .D(n143), .CP(clk), .RN(n171), .Q(
        \mem[3][30] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][29]  ( .D(n142), .CP(clk), .RN(n171), .Q(
        \mem[3][29] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][28]  ( .D(n141), .CP(clk), .RN(n171), .Q(
        \mem[3][28] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][27]  ( .D(n140), .CP(clk), .RN(n171), .Q(
        \mem[3][27] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][26]  ( .D(n139), .CP(clk), .RN(n171), .Q(
        \mem[3][26] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][25]  ( .D(n138), .CP(clk), .RN(n171), .Q(
        \mem[3][25] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][24]  ( .D(n137), .CP(clk), .RN(n171), .Q(
        \mem[3][24] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][23]  ( .D(n136), .CP(clk), .RN(n171), .Q(
        \mem[3][23] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][22]  ( .D(n135), .CP(clk), .RN(n171), .Q(
        \mem[3][22] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][21]  ( .D(n134), .CP(clk), .RN(n171), .Q(
        \mem[3][21] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][20]  ( .D(n133), .CP(clk), .RN(n171), .Q(
        \mem[3][20] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][19]  ( .D(n132), .CP(clk), .RN(n171), .Q(
        \mem[3][19] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][18]  ( .D(n131), .CP(clk), .RN(n172), .Q(
        \mem[3][18] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][17]  ( .D(n130), .CP(clk), .RN(n172), .Q(
        \mem[3][17] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][16]  ( .D(n129), .CP(clk), .RN(n172), .Q(
        \mem[3][16] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][15]  ( .D(n128), .CP(clk), .RN(n172), .Q(
        \mem[3][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][14]  ( .D(n127), .CP(clk), .RN(n172), .Q(
        \mem[3][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][13]  ( .D(n126), .CP(clk), .RN(n172), .Q(
        \mem[3][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][12]  ( .D(n125), .CP(clk), .RN(n172), .Q(
        \mem[3][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][11]  ( .D(n124), .CP(clk), .RN(n172), .Q(
        \mem[3][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][10]  ( .D(n123), .CP(clk), .RN(n172), .Q(
        \mem[3][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][9]  ( .D(n122), .CP(clk), .RN(n172), .Q(
        \mem[3][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][8]  ( .D(n121), .CP(clk), .RN(n172), .Q(
        \mem[3][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][7]  ( .D(n120), .CP(clk), .RN(n172), .Q(
        \mem[3][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][6]  ( .D(n119), .CP(clk), .RN(n172), .Q(
        \mem[3][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][5]  ( .D(n118), .CP(clk), .RN(n173), .Q(
        \mem[3][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][4]  ( .D(n117), .CP(clk), .RN(n173), .Q(
        \mem[3][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][3]  ( .D(n116), .CP(clk), .RN(n173), .Q(
        \mem[3][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][2]  ( .D(n115), .CP(clk), .RN(n173), .Q(
        \mem[3][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][1]  ( .D(n114), .CP(clk), .RN(n173), .Q(
        \mem[3][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][0]  ( .D(n113), .CP(clk), .RN(n173), .Q(
        \mem[3][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][31]  ( .D(n112), .CP(clk), .RN(n173), .Q(
        \mem[2][31] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][30]  ( .D(n111), .CP(clk), .RN(n173), .Q(
        \mem[2][30] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][29]  ( .D(n110), .CP(clk), .RN(n173), .Q(
        \mem[2][29] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][28]  ( .D(n109), .CP(clk), .RN(n173), .Q(
        \mem[2][28] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][27]  ( .D(n108), .CP(clk), .RN(n173), .Q(
        \mem[2][27] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][26]  ( .D(n107), .CP(clk), .RN(n173), .Q(
        \mem[2][26] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][25]  ( .D(n106), .CP(clk), .RN(n173), .Q(
        \mem[2][25] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][24]  ( .D(n105), .CP(clk), .RN(n174), .Q(
        \mem[2][24] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][23]  ( .D(n104), .CP(clk), .RN(n174), .Q(
        \mem[2][23] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][22]  ( .D(n103), .CP(clk), .RN(n174), .Q(
        \mem[2][22] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][21]  ( .D(n102), .CP(clk), .RN(n174), .Q(
        \mem[2][21] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][20]  ( .D(n101), .CP(clk), .RN(n174), .Q(
        \mem[2][20] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][19]  ( .D(n100), .CP(clk), .RN(n174), .Q(
        \mem[2][19] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][18]  ( .D(n99), .CP(clk), .RN(n174), .Q(
        \mem[2][18] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][17]  ( .D(n98), .CP(clk), .RN(n174), .Q(
        \mem[2][17] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][16]  ( .D(n97), .CP(clk), .RN(n174), .Q(
        \mem[2][16] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][15]  ( .D(n96), .CP(clk), .RN(n174), .Q(
        \mem[2][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][14]  ( .D(n95), .CP(clk), .RN(n174), .Q(
        \mem[2][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][13]  ( .D(n94), .CP(clk), .RN(n174), .Q(
        \mem[2][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][12]  ( .D(n93), .CP(clk), .RN(n174), .Q(
        \mem[2][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][11]  ( .D(n92), .CP(clk), .RN(n175), .Q(
        \mem[2][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][10]  ( .D(n91), .CP(clk), .RN(n175), .Q(
        \mem[2][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][9]  ( .D(n90), .CP(clk), .RN(n175), .Q(
        \mem[2][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][8]  ( .D(n89), .CP(clk), .RN(n175), .Q(
        \mem[2][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][7]  ( .D(n88), .CP(clk), .RN(n175), .Q(
        \mem[2][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][6]  ( .D(n87), .CP(clk), .RN(n175), .Q(
        \mem[2][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][5]  ( .D(n86), .CP(clk), .RN(n175), .Q(
        \mem[2][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][4]  ( .D(n85), .CP(clk), .RN(n175), .Q(
        \mem[2][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][3]  ( .D(n84), .CP(clk), .RN(n175), .Q(
        \mem[2][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][2]  ( .D(n83), .CP(clk), .RN(n175), .Q(
        \mem[2][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][1]  ( .D(n82), .CP(clk), .RN(n175), .Q(
        \mem[2][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][0]  ( .D(n81), .CP(clk), .RN(n175), .Q(
        \mem[2][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][31]  ( .D(n80), .CP(clk), .RN(n175), .Q(
        \mem[1][31] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][30]  ( .D(n79), .CP(clk), .RN(n176), .Q(
        \mem[1][30] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][29]  ( .D(n78), .CP(clk), .RN(n176), .Q(
        \mem[1][29] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][28]  ( .D(n77), .CP(clk), .RN(n176), .Q(
        \mem[1][28] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][27]  ( .D(n76), .CP(clk), .RN(n176), .Q(
        \mem[1][27] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][26]  ( .D(n75), .CP(clk), .RN(n176), .Q(
        \mem[1][26] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][25]  ( .D(n74), .CP(clk), .RN(n176), .Q(
        \mem[1][25] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][24]  ( .D(n73), .CP(clk), .RN(n176), .Q(
        \mem[1][24] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][23]  ( .D(n72), .CP(clk), .RN(n176), .Q(
        \mem[1][23] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][22]  ( .D(n71), .CP(clk), .RN(n176), .Q(
        \mem[1][22] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][21]  ( .D(n70), .CP(clk), .RN(n176), .Q(
        \mem[1][21] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][20]  ( .D(n69), .CP(clk), .RN(n176), .Q(
        \mem[1][20] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][19]  ( .D(n68), .CP(clk), .RN(n176), .Q(
        \mem[1][19] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][18]  ( .D(n67), .CP(clk), .RN(n176), .Q(
        \mem[1][18] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][17]  ( .D(n66), .CP(clk), .RN(n177), .Q(
        \mem[1][17] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][16]  ( .D(n65), .CP(clk), .RN(n177), .Q(
        \mem[1][16] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][15]  ( .D(n64), .CP(clk), .RN(n177), .Q(
        \mem[1][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][14]  ( .D(n63), .CP(clk), .RN(n177), .Q(
        \mem[1][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][13]  ( .D(n62), .CP(clk), .RN(n177), .Q(
        \mem[1][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][12]  ( .D(n61), .CP(clk), .RN(n177), .Q(
        \mem[1][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][11]  ( .D(n60), .CP(clk), .RN(n177), .Q(
        \mem[1][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][10]  ( .D(n59), .CP(clk), .RN(n177), .Q(
        \mem[1][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][9]  ( .D(n58), .CP(clk), .RN(n177), .Q(
        \mem[1][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][8]  ( .D(n57), .CP(clk), .RN(n177), .Q(
        \mem[1][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][7]  ( .D(n56), .CP(clk), .RN(n177), .Q(
        \mem[1][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][6]  ( .D(n55), .CP(clk), .RN(n177), .Q(
        \mem[1][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][5]  ( .D(n54), .CP(clk), .RN(n177), .Q(
        \mem[1][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][4]  ( .D(n53), .CP(clk), .RN(n178), .Q(
        \mem[1][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][3]  ( .D(n52), .CP(clk), .RN(n178), .Q(
        \mem[1][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][2]  ( .D(n51), .CP(clk), .RN(n178), .Q(
        \mem[1][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][1]  ( .D(n50), .CP(clk), .RN(n178), .Q(
        \mem[1][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][0]  ( .D(n49), .CP(clk), .RN(n178), .Q(
        \mem[1][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][31]  ( .D(n48), .CP(clk), .RN(n178), .Q(
        \mem[0][31] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][30]  ( .D(n47), .CP(clk), .RN(n178), .Q(
        \mem[0][30] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][29]  ( .D(n46), .CP(clk), .RN(n178), .Q(
        \mem[0][29] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][28]  ( .D(n45), .CP(clk), .RN(n178), .Q(
        \mem[0][28] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][27]  ( .D(n44), .CP(clk), .RN(n178), .Q(
        \mem[0][27] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][26]  ( .D(n43), .CP(clk), .RN(n178), .Q(
        \mem[0][26] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][25]  ( .D(n42), .CP(clk), .RN(n178), .Q(
        \mem[0][25] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][24]  ( .D(n41), .CP(clk), .RN(n178), .Q(
        \mem[0][24] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][23]  ( .D(n40), .CP(clk), .RN(n179), .Q(
        \mem[0][23] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][22]  ( .D(n39), .CP(clk), .RN(n179), .Q(
        \mem[0][22] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][21]  ( .D(n38), .CP(clk), .RN(n179), .Q(
        \mem[0][21] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][20]  ( .D(n37), .CP(clk), .RN(n179), .Q(
        \mem[0][20] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][19]  ( .D(n36), .CP(clk), .RN(n179), .Q(
        \mem[0][19] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][18]  ( .D(n35), .CP(clk), .RN(n179), .Q(
        \mem[0][18] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][17]  ( .D(n34), .CP(clk), .RN(n179), .Q(
        \mem[0][17] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][16]  ( .D(n33), .CP(clk), .RN(n179), .Q(
        \mem[0][16] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][15]  ( .D(n32), .CP(clk), .RN(n179), .Q(
        \mem[0][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][14]  ( .D(n31), .CP(clk), .RN(n179), .Q(
        \mem[0][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][13]  ( .D(n30), .CP(clk), .RN(n179), .Q(
        \mem[0][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][12]  ( .D(n29), .CP(clk), .RN(n179), .Q(
        \mem[0][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][11]  ( .D(n28), .CP(clk), .RN(n179), .Q(
        \mem[0][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][10]  ( .D(n27), .CP(clk), .RN(n180), .Q(
        \mem[0][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][9]  ( .D(n26), .CP(clk), .RN(n180), .Q(
        \mem[0][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][8]  ( .D(n25), .CP(clk), .RN(n180), .Q(
        \mem[0][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][7]  ( .D(n24), .CP(clk), .RN(n180), .Q(
        \mem[0][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][6]  ( .D(n23), .CP(clk), .RN(n180), .Q(
        \mem[0][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][5]  ( .D(n22), .CP(clk), .RN(n180), .Q(
        \mem[0][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][4]  ( .D(n21), .CP(clk), .RN(n180), .Q(
        \mem[0][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][3]  ( .D(n20), .CP(clk), .RN(n180), .Q(
        \mem[0][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][2]  ( .D(n19), .CP(clk), .RN(n180), .Q(
        \mem[0][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][1]  ( .D(n18), .CP(clk), .RN(n180), .Q(
        \mem[0][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][0]  ( .D(n17), .CP(clk), .RN(n180), .Q(
        \mem[0][0] ) );
  HS65_LS_DFPRQX9 \rd_data_reg[31]  ( .D(N17), .CP(clk), .RN(n180), .Q(
        rd_data[31]) );
  HS65_LS_DFPRQX9 \rd_data_reg[30]  ( .D(N18), .CP(clk), .RN(n180), .Q(
        rd_data[30]) );
  HS65_LS_DFPRQX9 \rd_data_reg[29]  ( .D(N19), .CP(clk), .RN(n181), .Q(
        rd_data[29]) );
  HS65_LS_DFPRQX9 \rd_data_reg[28]  ( .D(N20), .CP(clk), .RN(n181), .Q(
        rd_data[28]) );
  HS65_LS_DFPRQX9 \rd_data_reg[27]  ( .D(N21), .CP(clk), .RN(n181), .Q(
        rd_data[27]) );
  HS65_LS_DFPRQX9 \rd_data_reg[26]  ( .D(N22), .CP(clk), .RN(n181), .Q(
        rd_data[26]) );
  HS65_LS_DFPRQX9 \rd_data_reg[25]  ( .D(N23), .CP(clk), .RN(n181), .Q(
        rd_data[25]) );
  HS65_LS_DFPRQX9 \rd_data_reg[24]  ( .D(N24), .CP(clk), .RN(n181), .Q(
        rd_data[24]) );
  HS65_LS_DFPRQX9 \rd_data_reg[23]  ( .D(N25), .CP(clk), .RN(n181), .Q(
        rd_data[23]) );
  HS65_LS_DFPRQX9 \rd_data_reg[22]  ( .D(N26), .CP(clk), .RN(n181), .Q(
        rd_data[22]) );
  HS65_LS_DFPRQX9 \rd_data_reg[21]  ( .D(N27), .CP(clk), .RN(n181), .Q(
        rd_data[21]) );
  HS65_LS_DFPRQX9 \rd_data_reg[20]  ( .D(N28), .CP(clk), .RN(n181), .Q(
        rd_data[20]) );
  HS65_LS_DFPRQX9 \rd_data_reg[19]  ( .D(N29), .CP(clk), .RN(n181), .Q(
        rd_data[19]) );
  HS65_LS_DFPRQX9 \rd_data_reg[18]  ( .D(N30), .CP(clk), .RN(n181), .Q(
        rd_data[18]) );
  HS65_LS_DFPRQX9 \rd_data_reg[17]  ( .D(N31), .CP(clk), .RN(n181), .Q(
        rd_data[17]) );
  HS65_LS_DFPRQX9 \rd_data_reg[16]  ( .D(N32), .CP(clk), .RN(n182), .Q(
        rd_data[16]) );
  HS65_LS_DFPRQX9 \rd_data_reg[15]  ( .D(N33), .CP(clk), .RN(n182), .Q(
        rd_data[15]) );
  HS65_LS_DFPRQX9 \rd_data_reg[14]  ( .D(N34), .CP(clk), .RN(n182), .Q(
        rd_data[14]) );
  HS65_LS_DFPRQX9 \rd_data_reg[13]  ( .D(N35), .CP(clk), .RN(n182), .Q(
        rd_data[13]) );
  HS65_LS_DFPRQX9 \rd_data_reg[12]  ( .D(N36), .CP(clk), .RN(n182), .Q(
        rd_data[12]) );
  HS65_LS_DFPRQX9 \rd_data_reg[11]  ( .D(N37), .CP(clk), .RN(n182), .Q(
        rd_data[11]) );
  HS65_LS_DFPRQX9 \rd_data_reg[10]  ( .D(N38), .CP(clk), .RN(n182), .Q(
        rd_data[10]) );
  HS65_LS_DFPRQX9 \rd_data_reg[9]  ( .D(N39), .CP(clk), .RN(n182), .Q(
        rd_data[9]) );
  HS65_LS_DFPRQX9 \rd_data_reg[8]  ( .D(N40), .CP(clk), .RN(n182), .Q(
        rd_data[8]) );
  HS65_LS_DFPRQX9 \rd_data_reg[7]  ( .D(N41), .CP(clk), .RN(n182), .Q(
        rd_data[7]) );
  HS65_LS_DFPRQX9 \rd_data_reg[6]  ( .D(N42), .CP(clk), .RN(n182), .Q(
        rd_data[6]) );
  HS65_LS_DFPRQX9 \rd_data_reg[5]  ( .D(N43), .CP(clk), .RN(n182), .Q(
        rd_data[5]) );
  HS65_LS_DFPRQX9 \rd_data_reg[4]  ( .D(N44), .CP(clk), .RN(n182), .Q(
        rd_data[4]) );
  HS65_LS_DFPRQX9 \rd_data_reg[3]  ( .D(N45), .CP(clk), .RN(n183), .Q(
        rd_data[3]) );
  HS65_LS_DFPRQX9 \rd_data_reg[2]  ( .D(N46), .CP(clk), .RN(n183), .Q(
        rd_data[2]) );
  HS65_LS_DFPRQX9 \rd_data_reg[1]  ( .D(N47), .CP(clk), .RN(n183), .Q(
        rd_data[1]) );
  HS65_LS_DFPRQX9 \rd_data_reg[0]  ( .D(N48), .CP(clk), .RN(n183), .Q(
        rd_data[0]) );
  HS65_LS_AND3X9 U3 ( .A(n191), .B(n190), .C(wr_ena), .Z(n1) );
  HS65_LS_BFX9 U4 ( .A(n165), .Z(n162) );
  HS65_LS_BFX9 U5 ( .A(n1), .Z(n168) );
  HS65_LS_BFX9 U6 ( .A(n160), .Z(n157) );
  HS65_LS_BFX9 U7 ( .A(n155), .Z(n152) );
  HS65_LS_AND2X4 U8 ( .A(rd_addr[1]), .B(rd_addr[0]), .Z(n16) );
  HS65_LS_AND2X4 U9 ( .A(rd_addr[1]), .B(n192), .Z(n15) );
  HS65_LS_BFX9 U10 ( .A(n185), .Z(n180) );
  HS65_LS_BFX9 U11 ( .A(n185), .Z(n179) );
  HS65_LS_BFX9 U12 ( .A(n185), .Z(n178) );
  HS65_LS_BFX9 U13 ( .A(n186), .Z(n177) );
  HS65_LS_BFX9 U14 ( .A(n186), .Z(n176) );
  HS65_LS_BFX9 U15 ( .A(n186), .Z(n175) );
  HS65_LS_BFX9 U16 ( .A(n187), .Z(n174) );
  HS65_LS_BFX9 U17 ( .A(n187), .Z(n173) );
  HS65_LS_BFX9 U18 ( .A(n187), .Z(n172) );
  HS65_LS_BFX9 U19 ( .A(n188), .Z(n185) );
  HS65_LS_BFX9 U20 ( .A(n188), .Z(n186) );
  HS65_LS_BFX9 U21 ( .A(n189), .Z(n187) );
  HS65_LS_BFX9 U22 ( .A(n184), .Z(n182) );
  HS65_LS_BFX9 U23 ( .A(n184), .Z(n181) );
  HS65_LS_BFX9 U24 ( .A(n188), .Z(n171) );
  HS65_LS_BFX9 U25 ( .A(n189), .Z(n188) );
  HS65_LS_BFX9 U26 ( .A(n184), .Z(n183) );
  HS65_LS_BFX9 U27 ( .A(n189), .Z(n184) );
  HS65_LS_IVX9 U28 ( .A(reset), .Z(n189) );
  HS65_LS_IVX9 U29 ( .A(n168), .Z(n167) );
  HS65_LS_IVX9 U30 ( .A(n168), .Z(n166) );
  HS65_LS_IVX9 U31 ( .A(n162), .Z(n161) );
  HS65_LS_BFX9 U32 ( .A(n1), .Z(n169) );
  HS65_LS_BFX9 U33 ( .A(n165), .Z(n163) );
  HS65_LS_BFX9 U34 ( .A(n1), .Z(n170) );
  HS65_LS_BFX9 U35 ( .A(n162), .Z(n164) );
  HS65_LS_IVX9 U36 ( .A(n157), .Z(n156) );
  HS65_LS_IVX9 U37 ( .A(n152), .Z(n151) );
  HS65_LS_BFX9 U38 ( .A(n160), .Z(n158) );
  HS65_LS_BFX9 U39 ( .A(n155), .Z(n153) );
  HS65_LS_BFX9 U40 ( .A(n157), .Z(n159) );
  HS65_LS_BFX9 U41 ( .A(n152), .Z(n154) );
  HS65_LS_IVX9 U42 ( .A(n10), .Z(n165) );
  HS65_LS_IVX9 U43 ( .A(wr_addr[0]), .Z(n191) );
  HS65_LS_NAND3X5 U44 ( .A(wr_ena), .B(n190), .C(wr_addr[0]), .Z(n10) );
  HS65_LS_BFX9 U45 ( .A(n15), .Z(n6) );
  HS65_LS_BFX9 U46 ( .A(n15), .Z(n5) );
  HS65_LS_BFX9 U47 ( .A(n16), .Z(n3) );
  HS65_LS_BFX9 U48 ( .A(n16), .Z(n2) );
  HS65_LS_BFX9 U49 ( .A(n8), .Z(n145) );
  HS65_LS_BFX9 U50 ( .A(n8), .Z(n9) );
  HS65_LS_BFX9 U51 ( .A(n147), .Z(n149) );
  HS65_LS_BFX9 U52 ( .A(n147), .Z(n148) );
  HS65_LS_BFX9 U53 ( .A(n16), .Z(n4) );
  HS65_LS_BFX9 U54 ( .A(n15), .Z(n7) );
  HS65_LS_BFX9 U55 ( .A(n8), .Z(n146) );
  HS65_LS_BFX9 U56 ( .A(n147), .Z(n150) );
  HS65_LS_IVX9 U57 ( .A(n11), .Z(n160) );
  HS65_LS_IVX9 U58 ( .A(n12), .Z(n155) );
  HS65_LS_BFX9 U59 ( .A(n13), .Z(n147) );
  HS65_LS_NOR2X6 U60 ( .A(rd_addr[0]), .B(rd_addr[1]), .Z(n13) );
  HS65_LS_BFX9 U61 ( .A(n14), .Z(n8) );
  HS65_LS_NOR2X6 U62 ( .A(n192), .B(rd_addr[1]), .Z(n14) );
  HS65_LS_IVX9 U63 ( .A(wr_addr[1]), .Z(n190) );
  HS65_LS_IVX9 U64 ( .A(rd_addr[0]), .Z(n192) );
  HS65_LS_NAND3X5 U65 ( .A(wr_addr[0]), .B(wr_ena), .C(wr_addr[1]), .Z(n12) );
  HS65_LS_NAND3X5 U66 ( .A(wr_ena), .B(n191), .C(wr_addr[1]), .Z(n11) );
  HS65_LS_MX41X7 U67 ( .D0(n150), .S0(\mem[0][0] ), .D1(n146), .S1(\mem[1][0] ), .D2(n7), .S2(\mem[2][0] ), .D3(n4), .S3(\mem[3][0] ), .Z(N48) );
  HS65_LS_MX41X7 U68 ( .D0(n150), .S0(\mem[0][1] ), .D1(n146), .S1(\mem[1][1] ), .D2(n7), .S2(\mem[2][1] ), .D3(n4), .S3(\mem[3][1] ), .Z(N47) );
  HS65_LS_MX41X7 U69 ( .D0(n150), .S0(\mem[0][2] ), .D1(n146), .S1(\mem[1][2] ), .D2(n7), .S2(\mem[2][2] ), .D3(n4), .S3(\mem[3][2] ), .Z(N46) );
  HS65_LS_MX41X7 U70 ( .D0(n150), .S0(\mem[0][3] ), .D1(n146), .S1(\mem[1][3] ), .D2(n7), .S2(\mem[2][3] ), .D3(n4), .S3(\mem[3][3] ), .Z(N45) );
  HS65_LS_MX41X7 U71 ( .D0(n150), .S0(\mem[0][4] ), .D1(n146), .S1(\mem[1][4] ), .D2(n7), .S2(\mem[2][4] ), .D3(n4), .S3(\mem[3][4] ), .Z(N44) );
  HS65_LS_MX41X7 U72 ( .D0(n150), .S0(\mem[0][5] ), .D1(n146), .S1(\mem[1][5] ), .D2(n7), .S2(\mem[2][5] ), .D3(n4), .S3(\mem[3][5] ), .Z(N43) );
  HS65_LS_MX41X7 U73 ( .D0(n150), .S0(\mem[0][6] ), .D1(n146), .S1(\mem[1][6] ), .D2(n6), .S2(\mem[2][6] ), .D3(n4), .S3(\mem[3][6] ), .Z(N42) );
  HS65_LS_MX41X7 U74 ( .D0(n150), .S0(\mem[0][7] ), .D1(n146), .S1(\mem[1][7] ), .D2(n6), .S2(\mem[2][7] ), .D3(n4), .S3(\mem[3][7] ), .Z(N41) );
  HS65_LS_MX41X7 U75 ( .D0(n149), .S0(\mem[0][8] ), .D1(n145), .S1(\mem[1][8] ), .D2(n6), .S2(\mem[2][8] ), .D3(n3), .S3(\mem[3][8] ), .Z(N40) );
  HS65_LS_MX41X7 U76 ( .D0(n149), .S0(\mem[0][9] ), .D1(n145), .S1(\mem[1][9] ), .D2(n6), .S2(\mem[2][9] ), .D3(n3), .S3(\mem[3][9] ), .Z(N39) );
  HS65_LS_MX41X7 U77 ( .D0(n149), .S0(\mem[0][10] ), .D1(n145), .S1(
        \mem[1][10] ), .D2(n6), .S2(\mem[2][10] ), .D3(n3), .S3(\mem[3][10] ), 
        .Z(N38) );
  HS65_LS_MX41X7 U78 ( .D0(n149), .S0(\mem[0][11] ), .D1(n145), .S1(
        \mem[1][11] ), .D2(n6), .S2(\mem[2][11] ), .D3(n3), .S3(\mem[3][11] ), 
        .Z(N37) );
  HS65_LS_MX41X7 U79 ( .D0(n149), .S0(\mem[0][12] ), .D1(n145), .S1(
        \mem[1][12] ), .D2(n6), .S2(\mem[2][12] ), .D3(n3), .S3(\mem[3][12] ), 
        .Z(N36) );
  HS65_LS_MX41X7 U80 ( .D0(n149), .S0(\mem[0][13] ), .D1(n145), .S1(
        \mem[1][13] ), .D2(n6), .S2(\mem[2][13] ), .D3(n3), .S3(\mem[3][13] ), 
        .Z(N35) );
  HS65_LS_MX41X7 U81 ( .D0(n149), .S0(\mem[0][14] ), .D1(n145), .S1(
        \mem[1][14] ), .D2(n6), .S2(\mem[2][14] ), .D3(n3), .S3(\mem[3][14] ), 
        .Z(N34) );
  HS65_LS_MX41X7 U82 ( .D0(n149), .S0(\mem[0][15] ), .D1(n145), .S1(
        \mem[1][15] ), .D2(n6), .S2(\mem[2][15] ), .D3(n3), .S3(\mem[3][15] ), 
        .Z(N33) );
  HS65_LS_MX41X7 U83 ( .D0(n149), .S0(\mem[0][16] ), .D1(n145), .S1(
        \mem[1][16] ), .D2(n6), .S2(\mem[2][16] ), .D3(n3), .S3(\mem[3][16] ), 
        .Z(N32) );
  HS65_LS_MX41X7 U84 ( .D0(n149), .S0(\mem[0][17] ), .D1(n145), .S1(
        \mem[1][17] ), .D2(n6), .S2(\mem[2][17] ), .D3(n3), .S3(\mem[3][17] ), 
        .Z(N31) );
  HS65_LS_MX41X7 U85 ( .D0(n149), .S0(\mem[0][18] ), .D1(n145), .S1(
        \mem[1][18] ), .D2(n6), .S2(\mem[2][18] ), .D3(n3), .S3(\mem[3][18] ), 
        .Z(N30) );
  HS65_LS_MX41X7 U86 ( .D0(n149), .S0(\mem[0][19] ), .D1(n145), .S1(
        \mem[1][19] ), .D2(n5), .S2(\mem[2][19] ), .D3(n3), .S3(\mem[3][19] ), 
        .Z(N29) );
  HS65_LS_MX41X7 U87 ( .D0(n148), .S0(\mem[0][20] ), .D1(n9), .S1(\mem[1][20] ), .D2(n5), .S2(\mem[2][20] ), .D3(n2), .S3(\mem[3][20] ), .Z(N28) );
  HS65_LS_MX41X7 U88 ( .D0(n148), .S0(\mem[0][21] ), .D1(n9), .S1(\mem[1][21] ), .D2(n5), .S2(\mem[2][21] ), .D3(n2), .S3(\mem[3][21] ), .Z(N27) );
  HS65_LS_MX41X7 U89 ( .D0(n148), .S0(\mem[0][22] ), .D1(n9), .S1(\mem[1][22] ), .D2(n5), .S2(\mem[2][22] ), .D3(n2), .S3(\mem[3][22] ), .Z(N26) );
  HS65_LS_MX41X7 U90 ( .D0(n148), .S0(\mem[0][23] ), .D1(n9), .S1(\mem[1][23] ), .D2(n5), .S2(\mem[2][23] ), .D3(n2), .S3(\mem[3][23] ), .Z(N25) );
  HS65_LS_MX41X7 U91 ( .D0(n148), .S0(\mem[0][24] ), .D1(n9), .S1(\mem[1][24] ), .D2(n5), .S2(\mem[2][24] ), .D3(n2), .S3(\mem[3][24] ), .Z(N24) );
  HS65_LS_MX41X7 U92 ( .D0(n148), .S0(\mem[0][25] ), .D1(n9), .S1(\mem[1][25] ), .D2(n5), .S2(\mem[2][25] ), .D3(n2), .S3(\mem[3][25] ), .Z(N23) );
  HS65_LS_MX41X7 U93 ( .D0(n148), .S0(\mem[0][26] ), .D1(n9), .S1(\mem[1][26] ), .D2(n5), .S2(\mem[2][26] ), .D3(n2), .S3(\mem[3][26] ), .Z(N22) );
  HS65_LS_MX41X7 U94 ( .D0(n148), .S0(\mem[0][27] ), .D1(n9), .S1(\mem[1][27] ), .D2(n5), .S2(\mem[2][27] ), .D3(n2), .S3(\mem[3][27] ), .Z(N21) );
  HS65_LS_MX41X7 U95 ( .D0(n148), .S0(\mem[0][28] ), .D1(n9), .S1(\mem[1][28] ), .D2(n5), .S2(\mem[2][28] ), .D3(n2), .S3(\mem[3][28] ), .Z(N20) );
  HS65_LS_MX41X7 U96 ( .D0(n148), .S0(\mem[0][29] ), .D1(n9), .S1(\mem[1][29] ), .D2(n5), .S2(\mem[2][29] ), .D3(n2), .S3(\mem[3][29] ), .Z(N19) );
  HS65_LS_MX41X7 U97 ( .D0(n148), .S0(\mem[0][30] ), .D1(n9), .S1(\mem[1][30] ), .D2(n5), .S2(\mem[2][30] ), .D3(n2), .S3(\mem[3][30] ), .Z(N18) );
  HS65_LS_MX41X7 U98 ( .D0(n148), .S0(\mem[0][31] ), .D1(n9), .S1(\mem[1][31] ), .D2(n5), .S2(\mem[2][31] ), .D3(n2), .S3(\mem[3][31] ), .Z(N17) );
  HS65_LS_AO22X9 U99 ( .A(wr_data[0]), .B(n154), .C(n151), .D(\mem[3][0] ), 
        .Z(n113) );
  HS65_LS_AO22X9 U100 ( .A(wr_data[1]), .B(n154), .C(n151), .D(\mem[3][1] ), 
        .Z(n114) );
  HS65_LS_AO22X9 U101 ( .A(wr_data[2]), .B(n154), .C(n151), .D(\mem[3][2] ), 
        .Z(n115) );
  HS65_LS_AO22X9 U102 ( .A(wr_data[3]), .B(n154), .C(n151), .D(\mem[3][3] ), 
        .Z(n116) );
  HS65_LS_AO22X9 U103 ( .A(wr_data[4]), .B(n154), .C(n151), .D(\mem[3][4] ), 
        .Z(n117) );
  HS65_LS_AO22X9 U104 ( .A(wr_data[5]), .B(n154), .C(n151), .D(\mem[3][5] ), 
        .Z(n118) );
  HS65_LS_AO22X9 U105 ( .A(wr_data[6]), .B(n154), .C(n151), .D(\mem[3][6] ), 
        .Z(n119) );
  HS65_LS_AO22X9 U106 ( .A(wr_data[7]), .B(n154), .C(n151), .D(\mem[3][7] ), 
        .Z(n120) );
  HS65_LS_AO22X9 U107 ( .A(wr_data[8]), .B(n154), .C(n151), .D(\mem[3][8] ), 
        .Z(n121) );
  HS65_LS_AO22X9 U108 ( .A(wr_data[9]), .B(n154), .C(n151), .D(\mem[3][9] ), 
        .Z(n122) );
  HS65_LS_AO22X9 U109 ( .A(wr_data[10]), .B(n154), .C(n151), .D(\mem[3][10] ), 
        .Z(n123) );
  HS65_LS_AO22X9 U110 ( .A(wr_data[11]), .B(n153), .C(n151), .D(\mem[3][11] ), 
        .Z(n124) );
  HS65_LS_AO22X9 U111 ( .A(wr_data[12]), .B(n153), .C(n151), .D(\mem[3][12] ), 
        .Z(n125) );
  HS65_LS_AO22X9 U112 ( .A(wr_data[13]), .B(n153), .C(n151), .D(\mem[3][13] ), 
        .Z(n126) );
  HS65_LS_AO22X9 U113 ( .A(wr_data[14]), .B(n153), .C(n151), .D(\mem[3][14] ), 
        .Z(n127) );
  HS65_LS_AO22X9 U114 ( .A(wr_data[15]), .B(n153), .C(n151), .D(\mem[3][15] ), 
        .Z(n128) );
  HS65_LS_AO22X9 U115 ( .A(wr_data[16]), .B(n153), .C(n151), .D(\mem[3][16] ), 
        .Z(n129) );
  HS65_LS_AO22X9 U116 ( .A(wr_data[17]), .B(n153), .C(n151), .D(\mem[3][17] ), 
        .Z(n130) );
  HS65_LS_AO22X9 U117 ( .A(wr_data[18]), .B(n153), .C(n151), .D(\mem[3][18] ), 
        .Z(n131) );
  HS65_LS_AO22X9 U118 ( .A(wr_data[19]), .B(n153), .C(n151), .D(\mem[3][19] ), 
        .Z(n132) );
  HS65_LS_AO22X9 U119 ( .A(wr_data[20]), .B(n153), .C(n12), .D(\mem[3][20] ), 
        .Z(n133) );
  HS65_LS_AO22X9 U120 ( .A(wr_data[21]), .B(n153), .C(n12), .D(\mem[3][21] ), 
        .Z(n134) );
  HS65_LS_AO22X9 U121 ( .A(wr_data[22]), .B(n153), .C(n12), .D(\mem[3][22] ), 
        .Z(n135) );
  HS65_LS_AO22X9 U122 ( .A(wr_data[23]), .B(n153), .C(n12), .D(\mem[3][23] ), 
        .Z(n136) );
  HS65_LS_AO22X9 U123 ( .A(wr_data[24]), .B(n153), .C(n12), .D(\mem[3][24] ), 
        .Z(n137) );
  HS65_LS_AO22X9 U124 ( .A(wr_data[25]), .B(n153), .C(n12), .D(\mem[3][25] ), 
        .Z(n138) );
  HS65_LS_AO22X9 U125 ( .A(wr_data[26]), .B(n153), .C(n12), .D(\mem[3][26] ), 
        .Z(n139) );
  HS65_LS_AO22X9 U126 ( .A(wr_data[27]), .B(n153), .C(n12), .D(\mem[3][27] ), 
        .Z(n140) );
  HS65_LS_AO22X9 U127 ( .A(wr_data[28]), .B(n153), .C(n12), .D(\mem[3][28] ), 
        .Z(n141) );
  HS65_LS_AO22X9 U128 ( .A(wr_data[29]), .B(n153), .C(n12), .D(\mem[3][29] ), 
        .Z(n142) );
  HS65_LS_AO22X9 U129 ( .A(wr_data[30]), .B(n153), .C(n12), .D(\mem[3][30] ), 
        .Z(n143) );
  HS65_LS_AO22X9 U130 ( .A(wr_data[31]), .B(n152), .C(n12), .D(\mem[3][31] ), 
        .Z(n144) );
  HS65_LS_AO22X9 U131 ( .A(wr_data[0]), .B(n164), .C(n161), .D(\mem[1][0] ), 
        .Z(n49) );
  HS65_LS_AO22X9 U132 ( .A(wr_data[1]), .B(n164), .C(n161), .D(\mem[1][1] ), 
        .Z(n50) );
  HS65_LS_AO22X9 U133 ( .A(wr_data[2]), .B(n164), .C(n161), .D(\mem[1][2] ), 
        .Z(n51) );
  HS65_LS_AO22X9 U134 ( .A(wr_data[3]), .B(n164), .C(n161), .D(\mem[1][3] ), 
        .Z(n52) );
  HS65_LS_AO22X9 U135 ( .A(wr_data[4]), .B(n164), .C(n161), .D(\mem[1][4] ), 
        .Z(n53) );
  HS65_LS_AO22X9 U136 ( .A(wr_data[5]), .B(n164), .C(n161), .D(\mem[1][5] ), 
        .Z(n54) );
  HS65_LS_AO22X9 U137 ( .A(wr_data[6]), .B(n164), .C(n161), .D(\mem[1][6] ), 
        .Z(n55) );
  HS65_LS_AO22X9 U138 ( .A(wr_data[7]), .B(n164), .C(n161), .D(\mem[1][7] ), 
        .Z(n56) );
  HS65_LS_AO22X9 U139 ( .A(wr_data[8]), .B(n164), .C(n161), .D(\mem[1][8] ), 
        .Z(n57) );
  HS65_LS_AO22X9 U140 ( .A(wr_data[9]), .B(n164), .C(n161), .D(\mem[1][9] ), 
        .Z(n58) );
  HS65_LS_AO22X9 U141 ( .A(wr_data[10]), .B(n164), .C(n161), .D(\mem[1][10] ), 
        .Z(n59) );
  HS65_LS_AO22X9 U142 ( .A(wr_data[11]), .B(n163), .C(n161), .D(\mem[1][11] ), 
        .Z(n60) );
  HS65_LS_AO22X9 U143 ( .A(wr_data[12]), .B(n163), .C(n161), .D(\mem[1][12] ), 
        .Z(n61) );
  HS65_LS_AO22X9 U144 ( .A(wr_data[13]), .B(n163), .C(n161), .D(\mem[1][13] ), 
        .Z(n62) );
  HS65_LS_AO22X9 U145 ( .A(wr_data[14]), .B(n163), .C(n161), .D(\mem[1][14] ), 
        .Z(n63) );
  HS65_LS_AO22X9 U146 ( .A(wr_data[15]), .B(n163), .C(n161), .D(\mem[1][15] ), 
        .Z(n64) );
  HS65_LS_AO22X9 U147 ( .A(wr_data[16]), .B(n163), .C(n161), .D(\mem[1][16] ), 
        .Z(n65) );
  HS65_LS_AO22X9 U148 ( .A(wr_data[17]), .B(n163), .C(n161), .D(\mem[1][17] ), 
        .Z(n66) );
  HS65_LS_AO22X9 U149 ( .A(wr_data[18]), .B(n163), .C(n161), .D(\mem[1][18] ), 
        .Z(n67) );
  HS65_LS_AO22X9 U150 ( .A(wr_data[19]), .B(n163), .C(n161), .D(\mem[1][19] ), 
        .Z(n68) );
  HS65_LS_AO22X9 U151 ( .A(wr_data[20]), .B(n163), .C(n10), .D(\mem[1][20] ), 
        .Z(n69) );
  HS65_LS_AO22X9 U152 ( .A(wr_data[21]), .B(n163), .C(n10), .D(\mem[1][21] ), 
        .Z(n70) );
  HS65_LS_AO22X9 U153 ( .A(wr_data[22]), .B(n163), .C(n10), .D(\mem[1][22] ), 
        .Z(n71) );
  HS65_LS_AO22X9 U154 ( .A(wr_data[23]), .B(n163), .C(n10), .D(\mem[1][23] ), 
        .Z(n72) );
  HS65_LS_AO22X9 U155 ( .A(wr_data[24]), .B(n163), .C(n10), .D(\mem[1][24] ), 
        .Z(n73) );
  HS65_LS_AO22X9 U156 ( .A(wr_data[25]), .B(n163), .C(n10), .D(\mem[1][25] ), 
        .Z(n74) );
  HS65_LS_AO22X9 U157 ( .A(wr_data[26]), .B(n163), .C(n10), .D(\mem[1][26] ), 
        .Z(n75) );
  HS65_LS_AO22X9 U158 ( .A(wr_data[27]), .B(n163), .C(n10), .D(\mem[1][27] ), 
        .Z(n76) );
  HS65_LS_AO22X9 U159 ( .A(wr_data[28]), .B(n163), .C(n10), .D(\mem[1][28] ), 
        .Z(n77) );
  HS65_LS_AO22X9 U160 ( .A(wr_data[29]), .B(n163), .C(n10), .D(\mem[1][29] ), 
        .Z(n78) );
  HS65_LS_AO22X9 U161 ( .A(wr_data[30]), .B(n163), .C(n10), .D(\mem[1][30] ), 
        .Z(n79) );
  HS65_LS_AO22X9 U162 ( .A(wr_data[31]), .B(n162), .C(n10), .D(\mem[1][31] ), 
        .Z(n80) );
  HS65_LS_AO22X9 U163 ( .A(n170), .B(wr_data[0]), .C(n167), .D(\mem[0][0] ), 
        .Z(n17) );
  HS65_LS_AO22X9 U164 ( .A(n170), .B(wr_data[1]), .C(n166), .D(\mem[0][1] ), 
        .Z(n18) );
  HS65_LS_AO22X9 U165 ( .A(n170), .B(wr_data[2]), .C(n167), .D(\mem[0][2] ), 
        .Z(n19) );
  HS65_LS_AO22X9 U166 ( .A(n170), .B(wr_data[3]), .C(n166), .D(\mem[0][3] ), 
        .Z(n20) );
  HS65_LS_AO22X9 U167 ( .A(n170), .B(wr_data[4]), .C(n167), .D(\mem[0][4] ), 
        .Z(n21) );
  HS65_LS_AO22X9 U168 ( .A(n170), .B(wr_data[5]), .C(n166), .D(\mem[0][5] ), 
        .Z(n22) );
  HS65_LS_AO22X9 U169 ( .A(n170), .B(wr_data[6]), .C(n167), .D(\mem[0][6] ), 
        .Z(n23) );
  HS65_LS_AO22X9 U170 ( .A(n170), .B(wr_data[7]), .C(n167), .D(\mem[0][7] ), 
        .Z(n24) );
  HS65_LS_AO22X9 U171 ( .A(n170), .B(wr_data[8]), .C(n167), .D(\mem[0][8] ), 
        .Z(n25) );
  HS65_LS_AO22X9 U172 ( .A(n170), .B(wr_data[9]), .C(n167), .D(\mem[0][9] ), 
        .Z(n26) );
  HS65_LS_AO22X9 U173 ( .A(n170), .B(wr_data[10]), .C(n167), .D(\mem[0][10] ), 
        .Z(n27) );
  HS65_LS_AO22X9 U174 ( .A(n169), .B(wr_data[11]), .C(n167), .D(\mem[0][11] ), 
        .Z(n28) );
  HS65_LS_AO22X9 U175 ( .A(n169), .B(wr_data[12]), .C(n167), .D(\mem[0][12] ), 
        .Z(n29) );
  HS65_LS_AO22X9 U176 ( .A(n169), .B(wr_data[13]), .C(n167), .D(\mem[0][13] ), 
        .Z(n30) );
  HS65_LS_AO22X9 U177 ( .A(n169), .B(wr_data[14]), .C(n167), .D(\mem[0][14] ), 
        .Z(n31) );
  HS65_LS_AO22X9 U178 ( .A(n169), .B(wr_data[15]), .C(n167), .D(\mem[0][15] ), 
        .Z(n32) );
  HS65_LS_AO22X9 U179 ( .A(n169), .B(wr_data[16]), .C(n167), .D(\mem[0][16] ), 
        .Z(n33) );
  HS65_LS_AO22X9 U180 ( .A(n169), .B(wr_data[17]), .C(n167), .D(\mem[0][17] ), 
        .Z(n34) );
  HS65_LS_AO22X9 U181 ( .A(n169), .B(wr_data[18]), .C(n167), .D(\mem[0][18] ), 
        .Z(n35) );
  HS65_LS_AO22X9 U182 ( .A(n169), .B(wr_data[19]), .C(n166), .D(\mem[0][19] ), 
        .Z(n36) );
  HS65_LS_AO22X9 U183 ( .A(n169), .B(wr_data[20]), .C(n166), .D(\mem[0][20] ), 
        .Z(n37) );
  HS65_LS_AO22X9 U184 ( .A(n169), .B(wr_data[21]), .C(n166), .D(\mem[0][21] ), 
        .Z(n38) );
  HS65_LS_AO22X9 U185 ( .A(n169), .B(wr_data[22]), .C(n166), .D(\mem[0][22] ), 
        .Z(n39) );
  HS65_LS_AO22X9 U186 ( .A(n169), .B(wr_data[23]), .C(n166), .D(\mem[0][23] ), 
        .Z(n40) );
  HS65_LS_AO22X9 U187 ( .A(n169), .B(wr_data[24]), .C(n166), .D(\mem[0][24] ), 
        .Z(n41) );
  HS65_LS_AO22X9 U188 ( .A(n169), .B(wr_data[25]), .C(n166), .D(\mem[0][25] ), 
        .Z(n42) );
  HS65_LS_AO22X9 U189 ( .A(n169), .B(wr_data[26]), .C(n166), .D(\mem[0][26] ), 
        .Z(n43) );
  HS65_LS_AO22X9 U190 ( .A(n169), .B(wr_data[27]), .C(n166), .D(\mem[0][27] ), 
        .Z(n44) );
  HS65_LS_AO22X9 U191 ( .A(n169), .B(wr_data[28]), .C(n166), .D(\mem[0][28] ), 
        .Z(n45) );
  HS65_LS_AO22X9 U192 ( .A(n169), .B(wr_data[29]), .C(n166), .D(\mem[0][29] ), 
        .Z(n46) );
  HS65_LS_AO22X9 U193 ( .A(n169), .B(wr_data[30]), .C(n166), .D(\mem[0][30] ), 
        .Z(n47) );
  HS65_LS_AO22X9 U194 ( .A(n168), .B(wr_data[31]), .C(n166), .D(\mem[0][31] ), 
        .Z(n48) );
  HS65_LS_AO22X9 U195 ( .A(wr_data[0]), .B(n159), .C(n156), .D(\mem[2][0] ), 
        .Z(n81) );
  HS65_LS_AO22X9 U196 ( .A(wr_data[1]), .B(n159), .C(n156), .D(\mem[2][1] ), 
        .Z(n82) );
  HS65_LS_AO22X9 U197 ( .A(wr_data[2]), .B(n159), .C(n156), .D(\mem[2][2] ), 
        .Z(n83) );
  HS65_LS_AO22X9 U198 ( .A(wr_data[3]), .B(n159), .C(n156), .D(\mem[2][3] ), 
        .Z(n84) );
  HS65_LS_AO22X9 U199 ( .A(wr_data[4]), .B(n159), .C(n156), .D(\mem[2][4] ), 
        .Z(n85) );
  HS65_LS_AO22X9 U200 ( .A(wr_data[5]), .B(n159), .C(n156), .D(\mem[2][5] ), 
        .Z(n86) );
  HS65_LS_AO22X9 U201 ( .A(wr_data[6]), .B(n159), .C(n156), .D(\mem[2][6] ), 
        .Z(n87) );
  HS65_LS_AO22X9 U202 ( .A(wr_data[7]), .B(n159), .C(n156), .D(\mem[2][7] ), 
        .Z(n88) );
  HS65_LS_AO22X9 U203 ( .A(wr_data[8]), .B(n159), .C(n156), .D(\mem[2][8] ), 
        .Z(n89) );
  HS65_LS_AO22X9 U204 ( .A(wr_data[9]), .B(n159), .C(n156), .D(\mem[2][9] ), 
        .Z(n90) );
  HS65_LS_AO22X9 U205 ( .A(wr_data[10]), .B(n159), .C(n156), .D(\mem[2][10] ), 
        .Z(n91) );
  HS65_LS_AO22X9 U206 ( .A(wr_data[11]), .B(n158), .C(n156), .D(\mem[2][11] ), 
        .Z(n92) );
  HS65_LS_AO22X9 U207 ( .A(wr_data[12]), .B(n158), .C(n156), .D(\mem[2][12] ), 
        .Z(n93) );
  HS65_LS_AO22X9 U208 ( .A(wr_data[13]), .B(n158), .C(n156), .D(\mem[2][13] ), 
        .Z(n94) );
  HS65_LS_AO22X9 U209 ( .A(wr_data[14]), .B(n158), .C(n156), .D(\mem[2][14] ), 
        .Z(n95) );
  HS65_LS_AO22X9 U210 ( .A(wr_data[15]), .B(n158), .C(n156), .D(\mem[2][15] ), 
        .Z(n96) );
  HS65_LS_AO22X9 U211 ( .A(wr_data[16]), .B(n158), .C(n156), .D(\mem[2][16] ), 
        .Z(n97) );
  HS65_LS_AO22X9 U212 ( .A(wr_data[17]), .B(n158), .C(n156), .D(\mem[2][17] ), 
        .Z(n98) );
  HS65_LS_AO22X9 U213 ( .A(wr_data[18]), .B(n158), .C(n156), .D(\mem[2][18] ), 
        .Z(n99) );
  HS65_LS_AO22X9 U214 ( .A(wr_data[19]), .B(n158), .C(n156), .D(\mem[2][19] ), 
        .Z(n100) );
  HS65_LS_AO22X9 U215 ( .A(wr_data[20]), .B(n158), .C(n11), .D(\mem[2][20] ), 
        .Z(n101) );
  HS65_LS_AO22X9 U216 ( .A(wr_data[21]), .B(n158), .C(n11), .D(\mem[2][21] ), 
        .Z(n102) );
  HS65_LS_AO22X9 U217 ( .A(wr_data[22]), .B(n158), .C(n11), .D(\mem[2][22] ), 
        .Z(n103) );
  HS65_LS_AO22X9 U218 ( .A(wr_data[23]), .B(n158), .C(n11), .D(\mem[2][23] ), 
        .Z(n104) );
  HS65_LS_AO22X9 U219 ( .A(wr_data[24]), .B(n158), .C(n11), .D(\mem[2][24] ), 
        .Z(n105) );
  HS65_LS_AO22X9 U220 ( .A(wr_data[25]), .B(n158), .C(n11), .D(\mem[2][25] ), 
        .Z(n106) );
  HS65_LS_AO22X9 U221 ( .A(wr_data[26]), .B(n158), .C(n11), .D(\mem[2][26] ), 
        .Z(n107) );
  HS65_LS_AO22X9 U222 ( .A(wr_data[27]), .B(n158), .C(n11), .D(\mem[2][27] ), 
        .Z(n108) );
  HS65_LS_AO22X9 U223 ( .A(wr_data[28]), .B(n158), .C(n11), .D(\mem[2][28] ), 
        .Z(n109) );
  HS65_LS_AO22X9 U224 ( .A(wr_data[29]), .B(n158), .C(n11), .D(\mem[2][29] ), 
        .Z(n110) );
  HS65_LS_AO22X9 U225 ( .A(wr_data[30]), .B(n158), .C(n11), .D(\mem[2][30] ), 
        .Z(n111) );
  HS65_LS_AO22X9 U226 ( .A(wr_data[31]), .B(n157), .C(n11), .D(\mem[2][31] ), 
        .Z(n112) );
endmodule


module bram_DATA16_ADDR2_7 ( clk, reset, rd_addr, wr_addr, wr_data, wr_ena, 
        rd_data );
  input [1:0] rd_addr;
  input [1:0] wr_addr;
  input [15:0] wr_data;
  output [15:0] rd_data;
  input clk, reset, wr_ena;
  wire   \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] ,
         \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][15] , \mem[1][14] , \mem[1][13] ,
         \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] , \mem[1][8] ,
         \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] ,
         \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][15] , \mem[0][14] ,
         \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] ,
         \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] ,
         \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, n1,
         n2, n3, n4, n5, n6, n7, n8, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162;

  HS65_LS_DFPRQX9 \mem_reg[3][15]  ( .D(n91), .CP(clk), .RN(n1), .Q(
        \mem[3][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][14]  ( .D(n92), .CP(clk), .RN(n1), .Q(
        \mem[3][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][13]  ( .D(n93), .CP(clk), .RN(n1), .Q(
        \mem[3][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][12]  ( .D(n94), .CP(clk), .RN(n1), .Q(
        \mem[3][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][11]  ( .D(n95), .CP(clk), .RN(n1), .Q(
        \mem[3][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][10]  ( .D(n96), .CP(clk), .RN(n1), .Q(
        \mem[3][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][9]  ( .D(n97), .CP(clk), .RN(n1), .Q(\mem[3][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][8]  ( .D(n98), .CP(clk), .RN(n1), .Q(\mem[3][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][7]  ( .D(n99), .CP(clk), .RN(n1), .Q(\mem[3][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][6]  ( .D(n100), .CP(clk), .RN(n1), .Q(
        \mem[3][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][5]  ( .D(n101), .CP(clk), .RN(n1), .Q(
        \mem[3][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][4]  ( .D(n102), .CP(clk), .RN(n1), .Q(
        \mem[3][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][3]  ( .D(n103), .CP(clk), .RN(n1), .Q(
        \mem[3][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][2]  ( .D(n104), .CP(clk), .RN(n2), .Q(
        \mem[3][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][1]  ( .D(n105), .CP(clk), .RN(n2), .Q(
        \mem[3][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][0]  ( .D(n106), .CP(clk), .RN(n2), .Q(
        \mem[3][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][15]  ( .D(n107), .CP(clk), .RN(n2), .Q(
        \mem[2][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][14]  ( .D(n108), .CP(clk), .RN(n2), .Q(
        \mem[2][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][13]  ( .D(n109), .CP(clk), .RN(n2), .Q(
        \mem[2][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][12]  ( .D(n110), .CP(clk), .RN(n2), .Q(
        \mem[2][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][11]  ( .D(n111), .CP(clk), .RN(n2), .Q(
        \mem[2][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][10]  ( .D(n112), .CP(clk), .RN(n2), .Q(
        \mem[2][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][9]  ( .D(n113), .CP(clk), .RN(n2), .Q(
        \mem[2][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][8]  ( .D(n114), .CP(clk), .RN(n2), .Q(
        \mem[2][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][7]  ( .D(n115), .CP(clk), .RN(n2), .Q(
        \mem[2][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][6]  ( .D(n116), .CP(clk), .RN(n2), .Q(
        \mem[2][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][5]  ( .D(n117), .CP(clk), .RN(n3), .Q(
        \mem[2][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][4]  ( .D(n118), .CP(clk), .RN(n3), .Q(
        \mem[2][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][3]  ( .D(n119), .CP(clk), .RN(n3), .Q(
        \mem[2][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][2]  ( .D(n120), .CP(clk), .RN(n3), .Q(
        \mem[2][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][1]  ( .D(n121), .CP(clk), .RN(n3), .Q(
        \mem[2][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][0]  ( .D(n122), .CP(clk), .RN(n3), .Q(
        \mem[2][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][15]  ( .D(n123), .CP(clk), .RN(n3), .Q(
        \mem[1][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][14]  ( .D(n124), .CP(clk), .RN(n3), .Q(
        \mem[1][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][13]  ( .D(n125), .CP(clk), .RN(n3), .Q(
        \mem[1][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][12]  ( .D(n126), .CP(clk), .RN(n3), .Q(
        \mem[1][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][11]  ( .D(n127), .CP(clk), .RN(n3), .Q(
        \mem[1][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][10]  ( .D(n128), .CP(clk), .RN(n3), .Q(
        \mem[1][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][9]  ( .D(n129), .CP(clk), .RN(n3), .Q(
        \mem[1][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][8]  ( .D(n130), .CP(clk), .RN(n4), .Q(
        \mem[1][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][7]  ( .D(n131), .CP(clk), .RN(n4), .Q(
        \mem[1][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][6]  ( .D(n132), .CP(clk), .RN(n4), .Q(
        \mem[1][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][5]  ( .D(n133), .CP(clk), .RN(n4), .Q(
        \mem[1][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][4]  ( .D(n134), .CP(clk), .RN(n4), .Q(
        \mem[1][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][3]  ( .D(n135), .CP(clk), .RN(n4), .Q(
        \mem[1][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][2]  ( .D(n136), .CP(clk), .RN(n4), .Q(
        \mem[1][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][1]  ( .D(n137), .CP(clk), .RN(n4), .Q(
        \mem[1][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][0]  ( .D(n138), .CP(clk), .RN(n4), .Q(
        \mem[1][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][15]  ( .D(n139), .CP(clk), .RN(n4), .Q(
        \mem[0][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][14]  ( .D(n140), .CP(clk), .RN(n4), .Q(
        \mem[0][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][13]  ( .D(n141), .CP(clk), .RN(n4), .Q(
        \mem[0][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][12]  ( .D(n142), .CP(clk), .RN(n4), .Q(
        \mem[0][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][11]  ( .D(n143), .CP(clk), .RN(n5), .Q(
        \mem[0][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][10]  ( .D(n144), .CP(clk), .RN(n5), .Q(
        \mem[0][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][9]  ( .D(n145), .CP(clk), .RN(n5), .Q(
        \mem[0][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][8]  ( .D(n146), .CP(clk), .RN(n5), .Q(
        \mem[0][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][7]  ( .D(n147), .CP(clk), .RN(n5), .Q(
        \mem[0][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][6]  ( .D(n148), .CP(clk), .RN(n5), .Q(
        \mem[0][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][5]  ( .D(n149), .CP(clk), .RN(n5), .Q(
        \mem[0][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][4]  ( .D(n150), .CP(clk), .RN(n5), .Q(
        \mem[0][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][3]  ( .D(n151), .CP(clk), .RN(n5), .Q(
        \mem[0][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][2]  ( .D(n152), .CP(clk), .RN(n5), .Q(
        \mem[0][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][1]  ( .D(n153), .CP(clk), .RN(n5), .Q(
        \mem[0][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][0]  ( .D(n154), .CP(clk), .RN(n5), .Q(
        \mem[0][0] ) );
  HS65_LS_DFPRQX9 \rd_data_reg[15]  ( .D(N17), .CP(clk), .RN(n5), .Q(
        rd_data[15]) );
  HS65_LS_DFPRQX9 \rd_data_reg[14]  ( .D(N18), .CP(clk), .RN(n6), .Q(
        rd_data[14]) );
  HS65_LS_DFPRQX9 \rd_data_reg[13]  ( .D(N19), .CP(clk), .RN(n6), .Q(
        rd_data[13]) );
  HS65_LS_DFPRQX9 \rd_data_reg[12]  ( .D(N20), .CP(clk), .RN(n6), .Q(
        rd_data[12]) );
  HS65_LS_DFPRQX9 \rd_data_reg[11]  ( .D(N21), .CP(clk), .RN(n6), .Q(
        rd_data[11]) );
  HS65_LS_DFPRQX9 \rd_data_reg[10]  ( .D(N22), .CP(clk), .RN(n6), .Q(
        rd_data[10]) );
  HS65_LS_DFPRQX9 \rd_data_reg[9]  ( .D(N23), .CP(clk), .RN(n6), .Q(rd_data[9]) );
  HS65_LS_DFPRQX9 \rd_data_reg[8]  ( .D(N24), .CP(clk), .RN(n6), .Q(rd_data[8]) );
  HS65_LS_DFPRQX9 \rd_data_reg[7]  ( .D(N25), .CP(clk), .RN(n6), .Q(rd_data[7]) );
  HS65_LS_DFPRQX9 \rd_data_reg[6]  ( .D(N26), .CP(clk), .RN(n6), .Q(rd_data[6]) );
  HS65_LS_DFPRQX9 \rd_data_reg[5]  ( .D(N27), .CP(clk), .RN(n6), .Q(rd_data[5]) );
  HS65_LS_DFPRQX9 \rd_data_reg[4]  ( .D(N28), .CP(clk), .RN(n6), .Q(rd_data[4]) );
  HS65_LS_DFPRQX9 \rd_data_reg[3]  ( .D(N29), .CP(clk), .RN(n6), .Q(rd_data[3]) );
  HS65_LS_DFPRQX9 \rd_data_reg[2]  ( .D(N30), .CP(clk), .RN(n6), .Q(rd_data[2]) );
  HS65_LS_DFPRQX9 \rd_data_reg[1]  ( .D(N31), .CP(clk), .RN(n7), .Q(rd_data[1]) );
  HS65_LS_DFPRQX9 \rd_data_reg[0]  ( .D(N32), .CP(clk), .RN(n7), .Q(rd_data[0]) );
  HS65_LS_BFX9 U3 ( .A(n81), .Z(n4) );
  HS65_LS_BFX9 U4 ( .A(n81), .Z(n3) );
  HS65_LS_BFX9 U5 ( .A(n81), .Z(n2) );
  HS65_LS_BFX9 U6 ( .A(n83), .Z(n81) );
  HS65_LS_BFX9 U7 ( .A(n8), .Z(n6) );
  HS65_LS_BFX9 U8 ( .A(n8), .Z(n5) );
  HS65_LS_BFX9 U9 ( .A(n82), .Z(n1) );
  HS65_LS_BFX9 U10 ( .A(n83), .Z(n82) );
  HS65_LS_BFX9 U11 ( .A(n8), .Z(n7) );
  HS65_LS_BFX9 U12 ( .A(n83), .Z(n8) );
  HS65_LS_IVX9 U13 ( .A(reset), .Z(n83) );
  HS65_LS_IVX9 U14 ( .A(n161), .Z(n85) );
  HS65_LS_IVX9 U15 ( .A(n162), .Z(n84) );
  HS65_LS_NAND3X5 U16 ( .A(wr_ena), .B(n86), .C(wr_addr[0]), .Z(n161) );
  HS65_LS_IVX9 U17 ( .A(wr_addr[0]), .Z(n89) );
  HS65_LS_NAND3X5 U18 ( .A(n89), .B(n86), .C(wr_ena), .Z(n162) );
  HS65_LS_IVX9 U19 ( .A(n160), .Z(n88) );
  HS65_LS_IVX9 U20 ( .A(n159), .Z(n87) );
  HS65_LS_NAND3X5 U21 ( .A(wr_ena), .B(n89), .C(wr_addr[1]), .Z(n160) );
  HS65_LS_NOR2X6 U22 ( .A(n90), .B(rd_addr[1]), .Z(n157) );
  HS65_LS_NOR2X6 U23 ( .A(rd_addr[0]), .B(rd_addr[1]), .Z(n158) );
  HS65_LS_IVX9 U24 ( .A(wr_addr[1]), .Z(n86) );
  HS65_LS_NAND3X5 U25 ( .A(wr_addr[0]), .B(wr_ena), .C(wr_addr[1]), .Z(n159)
         );
  HS65_LS_AND2X4 U26 ( .A(rd_addr[1]), .B(n90), .Z(n156) );
  HS65_LS_AND2X4 U27 ( .A(rd_addr[1]), .B(rd_addr[0]), .Z(n155) );
  HS65_LS_IVX9 U28 ( .A(rd_addr[0]), .Z(n90) );
  HS65_LS_MX41X7 U29 ( .D0(n158), .S0(\mem[0][0] ), .D1(n157), .S1(\mem[1][0] ), .D2(n156), .S2(\mem[2][0] ), .D3(n155), .S3(\mem[3][0] ), .Z(N32) );
  HS65_LS_MX41X7 U30 ( .D0(n158), .S0(\mem[0][1] ), .D1(n157), .S1(\mem[1][1] ), .D2(n156), .S2(\mem[2][1] ), .D3(n155), .S3(\mem[3][1] ), .Z(N31) );
  HS65_LS_MX41X7 U31 ( .D0(n158), .S0(\mem[0][2] ), .D1(n157), .S1(\mem[1][2] ), .D2(n156), .S2(\mem[2][2] ), .D3(n155), .S3(\mem[3][2] ), .Z(N30) );
  HS65_LS_MX41X7 U32 ( .D0(n158), .S0(\mem[0][3] ), .D1(n157), .S1(\mem[1][3] ), .D2(n156), .S2(\mem[2][3] ), .D3(n155), .S3(\mem[3][3] ), .Z(N29) );
  HS65_LS_MX41X7 U33 ( .D0(n158), .S0(\mem[0][4] ), .D1(n157), .S1(\mem[1][4] ), .D2(n156), .S2(\mem[2][4] ), .D3(n155), .S3(\mem[3][4] ), .Z(N28) );
  HS65_LS_MX41X7 U34 ( .D0(n158), .S0(\mem[0][5] ), .D1(n157), .S1(\mem[1][5] ), .D2(n156), .S2(\mem[2][5] ), .D3(n155), .S3(\mem[3][5] ), .Z(N27) );
  HS65_LS_MX41X7 U35 ( .D0(n158), .S0(\mem[0][6] ), .D1(n157), .S1(\mem[1][6] ), .D2(n156), .S2(\mem[2][6] ), .D3(n155), .S3(\mem[3][6] ), .Z(N26) );
  HS65_LS_MX41X7 U36 ( .D0(n158), .S0(\mem[0][7] ), .D1(n157), .S1(\mem[1][7] ), .D2(n156), .S2(\mem[2][7] ), .D3(n155), .S3(\mem[3][7] ), .Z(N25) );
  HS65_LS_MX41X7 U37 ( .D0(n158), .S0(\mem[0][8] ), .D1(n157), .S1(\mem[1][8] ), .D2(n156), .S2(\mem[2][8] ), .D3(n155), .S3(\mem[3][8] ), .Z(N24) );
  HS65_LS_MX41X7 U38 ( .D0(n158), .S0(\mem[0][9] ), .D1(n157), .S1(\mem[1][9] ), .D2(n156), .S2(\mem[2][9] ), .D3(n155), .S3(\mem[3][9] ), .Z(N23) );
  HS65_LS_MX41X7 U39 ( .D0(n158), .S0(\mem[0][10] ), .D1(n157), .S1(
        \mem[1][10] ), .D2(n156), .S2(\mem[2][10] ), .D3(n155), .S3(
        \mem[3][10] ), .Z(N22) );
  HS65_LS_MX41X7 U40 ( .D0(n158), .S0(\mem[0][11] ), .D1(n157), .S1(
        \mem[1][11] ), .D2(n156), .S2(\mem[2][11] ), .D3(n155), .S3(
        \mem[3][11] ), .Z(N21) );
  HS65_LS_MX41X7 U41 ( .D0(n158), .S0(\mem[0][12] ), .D1(n157), .S1(
        \mem[1][12] ), .D2(n156), .S2(\mem[2][12] ), .D3(n155), .S3(
        \mem[3][12] ), .Z(N20) );
  HS65_LS_MX41X7 U42 ( .D0(n158), .S0(\mem[0][13] ), .D1(n157), .S1(
        \mem[1][13] ), .D2(n156), .S2(\mem[2][13] ), .D3(n155), .S3(
        \mem[3][13] ), .Z(N19) );
  HS65_LS_MX41X7 U43 ( .D0(n158), .S0(\mem[0][14] ), .D1(n157), .S1(
        \mem[1][14] ), .D2(n156), .S2(\mem[2][14] ), .D3(n155), .S3(
        \mem[3][14] ), .Z(N18) );
  HS65_LS_MX41X7 U44 ( .D0(n158), .S0(\mem[0][15] ), .D1(n157), .S1(
        \mem[1][15] ), .D2(n156), .S2(\mem[2][15] ), .D3(n155), .S3(
        \mem[3][15] ), .Z(N17) );
  HS65_LS_AO22X9 U45 ( .A(wr_data[0]), .B(n85), .C(n161), .D(\mem[1][0] ), .Z(
        n138) );
  HS65_LS_AO22X9 U46 ( .A(wr_data[1]), .B(n85), .C(n161), .D(\mem[1][1] ), .Z(
        n137) );
  HS65_LS_AO22X9 U47 ( .A(wr_data[2]), .B(n85), .C(n161), .D(\mem[1][2] ), .Z(
        n136) );
  HS65_LS_AO22X9 U48 ( .A(wr_data[3]), .B(n85), .C(n161), .D(\mem[1][3] ), .Z(
        n135) );
  HS65_LS_AO22X9 U49 ( .A(wr_data[4]), .B(n85), .C(n161), .D(\mem[1][4] ), .Z(
        n134) );
  HS65_LS_AO22X9 U50 ( .A(wr_data[5]), .B(n85), .C(n161), .D(\mem[1][5] ), .Z(
        n133) );
  HS65_LS_AO22X9 U51 ( .A(wr_data[6]), .B(n85), .C(n161), .D(\mem[1][6] ), .Z(
        n132) );
  HS65_LS_AO22X9 U52 ( .A(wr_data[7]), .B(n85), .C(n161), .D(\mem[1][7] ), .Z(
        n131) );
  HS65_LS_AO22X9 U53 ( .A(wr_data[8]), .B(n85), .C(n161), .D(\mem[1][8] ), .Z(
        n130) );
  HS65_LS_AO22X9 U54 ( .A(wr_data[9]), .B(n85), .C(n161), .D(\mem[1][9] ), .Z(
        n129) );
  HS65_LS_AO22X9 U55 ( .A(wr_data[10]), .B(n85), .C(n161), .D(\mem[1][10] ), 
        .Z(n128) );
  HS65_LS_AO22X9 U56 ( .A(wr_data[11]), .B(n85), .C(n161), .D(\mem[1][11] ), 
        .Z(n127) );
  HS65_LS_AO22X9 U57 ( .A(wr_data[12]), .B(n85), .C(n161), .D(\mem[1][12] ), 
        .Z(n126) );
  HS65_LS_AO22X9 U58 ( .A(wr_data[13]), .B(n85), .C(n161), .D(\mem[1][13] ), 
        .Z(n125) );
  HS65_LS_AO22X9 U59 ( .A(wr_data[14]), .B(n85), .C(n161), .D(\mem[1][14] ), 
        .Z(n124) );
  HS65_LS_AO22X9 U60 ( .A(wr_data[15]), .B(n85), .C(n161), .D(\mem[1][15] ), 
        .Z(n123) );
  HS65_LS_AO22X9 U61 ( .A(wr_data[0]), .B(n88), .C(n160), .D(\mem[2][0] ), .Z(
        n122) );
  HS65_LS_AO22X9 U62 ( .A(wr_data[1]), .B(n88), .C(n160), .D(\mem[2][1] ), .Z(
        n121) );
  HS65_LS_AO22X9 U63 ( .A(wr_data[2]), .B(n88), .C(n160), .D(\mem[2][2] ), .Z(
        n120) );
  HS65_LS_AO22X9 U64 ( .A(wr_data[3]), .B(n88), .C(n160), .D(\mem[2][3] ), .Z(
        n119) );
  HS65_LS_AO22X9 U65 ( .A(wr_data[4]), .B(n88), .C(n160), .D(\mem[2][4] ), .Z(
        n118) );
  HS65_LS_AO22X9 U66 ( .A(wr_data[5]), .B(n88), .C(n160), .D(\mem[2][5] ), .Z(
        n117) );
  HS65_LS_AO22X9 U67 ( .A(wr_data[6]), .B(n88), .C(n160), .D(\mem[2][6] ), .Z(
        n116) );
  HS65_LS_AO22X9 U68 ( .A(wr_data[7]), .B(n88), .C(n160), .D(\mem[2][7] ), .Z(
        n115) );
  HS65_LS_AO22X9 U69 ( .A(wr_data[8]), .B(n88), .C(n160), .D(\mem[2][8] ), .Z(
        n114) );
  HS65_LS_AO22X9 U70 ( .A(wr_data[9]), .B(n88), .C(n160), .D(\mem[2][9] ), .Z(
        n113) );
  HS65_LS_AO22X9 U71 ( .A(wr_data[10]), .B(n88), .C(n160), .D(\mem[2][10] ), 
        .Z(n112) );
  HS65_LS_AO22X9 U72 ( .A(wr_data[11]), .B(n88), .C(n160), .D(\mem[2][11] ), 
        .Z(n111) );
  HS65_LS_AO22X9 U73 ( .A(wr_data[12]), .B(n88), .C(n160), .D(\mem[2][12] ), 
        .Z(n110) );
  HS65_LS_AO22X9 U74 ( .A(wr_data[13]), .B(n88), .C(n160), .D(\mem[2][13] ), 
        .Z(n109) );
  HS65_LS_AO22X9 U75 ( .A(wr_data[14]), .B(n88), .C(n160), .D(\mem[2][14] ), 
        .Z(n108) );
  HS65_LS_AO22X9 U76 ( .A(wr_data[15]), .B(n88), .C(n160), .D(\mem[2][15] ), 
        .Z(n107) );
  HS65_LS_AO22X9 U77 ( .A(n84), .B(wr_data[0]), .C(n162), .D(\mem[0][0] ), .Z(
        n154) );
  HS65_LS_AO22X9 U78 ( .A(n84), .B(wr_data[1]), .C(n162), .D(\mem[0][1] ), .Z(
        n153) );
  HS65_LS_AO22X9 U79 ( .A(n84), .B(wr_data[2]), .C(n162), .D(\mem[0][2] ), .Z(
        n152) );
  HS65_LS_AO22X9 U80 ( .A(n84), .B(wr_data[3]), .C(n162), .D(\mem[0][3] ), .Z(
        n151) );
  HS65_LS_AO22X9 U81 ( .A(n84), .B(wr_data[4]), .C(n162), .D(\mem[0][4] ), .Z(
        n150) );
  HS65_LS_AO22X9 U82 ( .A(n84), .B(wr_data[5]), .C(n162), .D(\mem[0][5] ), .Z(
        n149) );
  HS65_LS_AO22X9 U83 ( .A(n84), .B(wr_data[6]), .C(n162), .D(\mem[0][6] ), .Z(
        n148) );
  HS65_LS_AO22X9 U84 ( .A(n84), .B(wr_data[7]), .C(n162), .D(\mem[0][7] ), .Z(
        n147) );
  HS65_LS_AO22X9 U85 ( .A(n84), .B(wr_data[8]), .C(n162), .D(\mem[0][8] ), .Z(
        n146) );
  HS65_LS_AO22X9 U86 ( .A(n84), .B(wr_data[9]), .C(n162), .D(\mem[0][9] ), .Z(
        n145) );
  HS65_LS_AO22X9 U87 ( .A(n84), .B(wr_data[10]), .C(n162), .D(\mem[0][10] ), 
        .Z(n144) );
  HS65_LS_AO22X9 U88 ( .A(n84), .B(wr_data[11]), .C(n162), .D(\mem[0][11] ), 
        .Z(n143) );
  HS65_LS_AO22X9 U89 ( .A(n84), .B(wr_data[12]), .C(n162), .D(\mem[0][12] ), 
        .Z(n142) );
  HS65_LS_AO22X9 U90 ( .A(n84), .B(wr_data[13]), .C(n162), .D(\mem[0][13] ), 
        .Z(n141) );
  HS65_LS_AO22X9 U91 ( .A(n84), .B(wr_data[14]), .C(n162), .D(\mem[0][14] ), 
        .Z(n140) );
  HS65_LS_AO22X9 U92 ( .A(n84), .B(wr_data[15]), .C(n162), .D(\mem[0][15] ), 
        .Z(n139) );
  HS65_LS_AO22X9 U93 ( .A(wr_data[0]), .B(n87), .C(n159), .D(\mem[3][0] ), .Z(
        n106) );
  HS65_LS_AO22X9 U94 ( .A(wr_data[1]), .B(n87), .C(n159), .D(\mem[3][1] ), .Z(
        n105) );
  HS65_LS_AO22X9 U95 ( .A(wr_data[2]), .B(n87), .C(n159), .D(\mem[3][2] ), .Z(
        n104) );
  HS65_LS_AO22X9 U96 ( .A(wr_data[3]), .B(n87), .C(n159), .D(\mem[3][3] ), .Z(
        n103) );
  HS65_LS_AO22X9 U97 ( .A(wr_data[4]), .B(n87), .C(n159), .D(\mem[3][4] ), .Z(
        n102) );
  HS65_LS_AO22X9 U98 ( .A(wr_data[5]), .B(n87), .C(n159), .D(\mem[3][5] ), .Z(
        n101) );
  HS65_LS_AO22X9 U99 ( .A(wr_data[6]), .B(n87), .C(n159), .D(\mem[3][6] ), .Z(
        n100) );
  HS65_LS_AO22X9 U100 ( .A(wr_data[7]), .B(n87), .C(n159), .D(\mem[3][7] ), 
        .Z(n99) );
  HS65_LS_AO22X9 U101 ( .A(wr_data[8]), .B(n87), .C(n159), .D(\mem[3][8] ), 
        .Z(n98) );
  HS65_LS_AO22X9 U102 ( .A(wr_data[9]), .B(n87), .C(n159), .D(\mem[3][9] ), 
        .Z(n97) );
  HS65_LS_AO22X9 U103 ( .A(wr_data[10]), .B(n87), .C(n159), .D(\mem[3][10] ), 
        .Z(n96) );
  HS65_LS_AO22X9 U104 ( .A(wr_data[11]), .B(n87), .C(n159), .D(\mem[3][11] ), 
        .Z(n95) );
  HS65_LS_AO22X9 U105 ( .A(wr_data[12]), .B(n87), .C(n159), .D(\mem[3][12] ), 
        .Z(n94) );
  HS65_LS_AO22X9 U106 ( .A(wr_data[13]), .B(n87), .C(n159), .D(\mem[3][13] ), 
        .Z(n93) );
  HS65_LS_AO22X9 U107 ( .A(wr_data[14]), .B(n87), .C(n159), .D(\mem[3][14] ), 
        .Z(n92) );
  HS65_LS_AO22X9 U108 ( .A(wr_data[15]), .B(n87), .C(n159), .D(\mem[3][15] ), 
        .Z(n91) );
endmodule


module dma_sdp_DATA64_ADDR2_0 ( clk, reset, ren, wen, waddr, wdata, raddr, 
        rdata );
  input [2:0] ren;
  input [2:0] wen;
  input [1:0] waddr;
  input [63:0] wdata;
  input [1:0] raddr;
  output [63:0] rdata;
  input clk, reset;
  wire   n37, n38, n39, n40, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n41, n42, n43, n44;
  wire   [2:0] sel_out;
  wire   [15:0] rdata0;
  wire   [31:0] rdata1;
  wire   [15:0] rdata2;

  HS65_LS_DFPRQX9 \sel_out_reg[2]  ( .D(ren[2]), .CP(clk), .RN(n5), .Q(
        sel_out[2]) );
  HS65_LS_DFPRQX9 \sel_out_reg[1]  ( .D(ren[1]), .CP(clk), .RN(n5), .Q(
        sel_out[1]) );
  HS65_LS_DFPRQX9 \sel_out_reg[0]  ( .D(ren[0]), .CP(clk), .RN(n5), .Q(
        sel_out[0]) );
  bram_DATA16_ADDR2_0 dma0 ( .clk(clk), .reset(reset), .rd_addr(raddr), 
        .wr_addr(waddr), .wr_data(wdata[63:48]), .wr_ena(wen[2]), .rd_data(
        rdata0) );
  bram_DATA32_ADDR2_0 dma1 ( .clk(clk), .reset(reset), .rd_addr(raddr), 
        .wr_addr(waddr), .wr_data(wdata[47:16]), .wr_ena(wen[1]), .rd_data(
        rdata1) );
  bram_DATA16_ADDR2_7 dma2 ( .clk(clk), .reset(reset), .rd_addr(raddr), 
        .wr_addr(waddr), .wr_data(wdata[15:0]), .wr_ena(wen[0]), .rd_data(
        rdata2) );
  HS65_LS_NAND3X5 U3 ( .A(sel_out[2]), .B(sel_out[1]), .C(sel_out[0]), .Z(n39)
         );
  HS65_LS_IVX9 U4 ( .A(reset), .Z(n5) );
  HS65_LS_NOR2X6 U5 ( .A(n2), .B(n13), .Z(rdata[40]) );
  HS65_LS_NOR2X6 U6 ( .A(n2), .B(n12), .Z(rdata[41]) );
  HS65_LS_NOR2X6 U7 ( .A(n2), .B(n11), .Z(rdata[42]) );
  HS65_LS_NOR2X6 U8 ( .A(n2), .B(n10), .Z(rdata[43]) );
  HS65_LS_NOR2X6 U9 ( .A(n2), .B(n9), .Z(rdata[44]) );
  HS65_LS_NOR2X6 U10 ( .A(n2), .B(n8), .Z(rdata[45]) );
  HS65_LS_NOR2X6 U11 ( .A(n2), .B(n7), .Z(rdata[46]) );
  HS65_LS_NOR2X6 U12 ( .A(n2), .B(n14), .Z(rdata[39]) );
  HS65_LS_BFX9 U13 ( .A(n39), .Z(n2) );
  HS65_LS_NOR2X6 U14 ( .A(n2), .B(n15), .Z(rdata[38]) );
  HS65_LS_NOR2X6 U15 ( .A(n3), .B(n19), .Z(rdata[34]) );
  HS65_LS_NOR2X6 U16 ( .A(n2), .B(n18), .Z(rdata[35]) );
  HS65_LS_NOR2X6 U17 ( .A(n3), .B(n17), .Z(rdata[36]) );
  HS65_LS_NOR2X6 U18 ( .A(n2), .B(n16), .Z(rdata[37]) );
  HS65_LS_NOR2X6 U19 ( .A(n3), .B(n20), .Z(rdata[33]) );
  HS65_LS_BFX9 U20 ( .A(n39), .Z(n3) );
  HS65_LS_BFX9 U21 ( .A(n39), .Z(n1) );
  HS65_LS_BFX9 U22 ( .A(n39), .Z(n4) );
  HS65_LS_IVX9 U23 ( .A(n40), .Z(n42) );
  HS65_LS_NOR2X6 U24 ( .A(n2), .B(n6), .Z(rdata[47]) );
  HS65_LS_NAND3X5 U25 ( .A(n44), .B(n43), .C(sel_out[1]), .Z(n40) );
  HS65_LS_IVX9 U26 ( .A(sel_out[0]), .Z(n44) );
  HS65_LS_IVX9 U27 ( .A(sel_out[2]), .Z(n43) );
  HS65_LS_OAI22X6 U28 ( .A(n40), .B(n19), .C(n1), .D(n35), .Z(rdata[18]) );
  HS65_LS_IVX9 U29 ( .A(rdata1[2]), .Z(n35) );
  HS65_LS_OAI22X6 U30 ( .A(n40), .B(n18), .C(n1), .D(n34), .Z(rdata[19]) );
  HS65_LS_IVX9 U31 ( .A(rdata1[3]), .Z(n34) );
  HS65_LS_OAI22X6 U32 ( .A(n40), .B(n17), .C(n1), .D(n33), .Z(rdata[20]) );
  HS65_LS_IVX9 U33 ( .A(rdata1[4]), .Z(n33) );
  HS65_LS_OAI22X6 U34 ( .A(n40), .B(n16), .C(n1), .D(n32), .Z(rdata[21]) );
  HS65_LS_IVX9 U35 ( .A(rdata1[5]), .Z(n32) );
  HS65_LS_OAI22X6 U36 ( .A(n40), .B(n15), .C(n31), .D(n3), .Z(rdata[22]) );
  HS65_LS_IVX9 U37 ( .A(rdata1[6]), .Z(n31) );
  HS65_LS_OAI22X6 U38 ( .A(n40), .B(n14), .C(n30), .D(n3), .Z(rdata[23]) );
  HS65_LS_IVX9 U39 ( .A(rdata1[7]), .Z(n30) );
  HS65_LS_OAI22X6 U40 ( .A(n40), .B(n13), .C(n29), .D(n3), .Z(rdata[24]) );
  HS65_LS_IVX9 U41 ( .A(rdata1[8]), .Z(n29) );
  HS65_LS_OAI22X6 U42 ( .A(n40), .B(n12), .C(n28), .D(n3), .Z(rdata[25]) );
  HS65_LS_IVX9 U43 ( .A(rdata1[9]), .Z(n28) );
  HS65_LS_OAI22X6 U44 ( .A(n40), .B(n11), .C(n1), .D(n27), .Z(rdata[26]) );
  HS65_LS_IVX9 U45 ( .A(rdata1[10]), .Z(n27) );
  HS65_LS_OAI22X6 U46 ( .A(n40), .B(n10), .C(n1), .D(n26), .Z(rdata[27]) );
  HS65_LS_IVX9 U47 ( .A(rdata1[11]), .Z(n26) );
  HS65_LS_OAI22X6 U48 ( .A(n40), .B(n20), .C(n1), .D(n36), .Z(rdata[17]) );
  HS65_LS_IVX9 U49 ( .A(rdata1[1]), .Z(n36) );
  HS65_LS_NOR2X6 U50 ( .A(n3), .B(n21), .Z(rdata[32]) );
  HS65_LS_NOR2AX3 U51 ( .A(rdata0[15]), .B(n3), .Z(rdata[63]) );
  HS65_LS_IVX9 U52 ( .A(rdata1[18]), .Z(n19) );
  HS65_LS_IVX9 U53 ( .A(rdata1[19]), .Z(n18) );
  HS65_LS_IVX9 U54 ( .A(rdata1[17]), .Z(n20) );
  HS65_LS_NOR2AX3 U55 ( .A(rdata0[3]), .B(n3), .Z(rdata[51]) );
  HS65_LS_NOR2AX3 U56 ( .A(rdata0[4]), .B(n4), .Z(rdata[52]) );
  HS65_LS_NOR2AX3 U57 ( .A(rdata0[7]), .B(n4), .Z(rdata[55]) );
  HS65_LS_NOR2AX3 U58 ( .A(rdata0[8]), .B(n4), .Z(rdata[56]) );
  HS65_LS_NOR2AX3 U59 ( .A(rdata0[10]), .B(n4), .Z(rdata[58]) );
  HS65_LS_NOR2AX3 U60 ( .A(rdata0[12]), .B(n4), .Z(rdata[60]) );
  HS65_LS_NOR2AX3 U61 ( .A(rdata0[1]), .B(n3), .Z(rdata[49]) );
  HS65_LS_NOR2AX3 U62 ( .A(rdata0[2]), .B(n3), .Z(rdata[50]) );
  HS65_LS_NOR2AX3 U63 ( .A(rdata0[5]), .B(n4), .Z(rdata[53]) );
  HS65_LS_NOR2AX3 U64 ( .A(rdata0[6]), .B(n4), .Z(rdata[54]) );
  HS65_LS_NOR2AX3 U65 ( .A(rdata0[9]), .B(n4), .Z(rdata[57]) );
  HS65_LS_NOR2AX3 U66 ( .A(rdata0[11]), .B(n4), .Z(rdata[59]) );
  HS65_LS_NOR2AX3 U67 ( .A(rdata0[14]), .B(n4), .Z(rdata[62]) );
  HS65_LS_OAI31X5 U68 ( .A(n44), .B(sel_out[2]), .C(sel_out[1]), .D(n2), .Z(
        n38) );
  HS65_LS_NOR3X4 U69 ( .A(sel_out[0]), .B(sel_out[1]), .C(n43), .Z(n37) );
  HS65_LS_OAI22X6 U70 ( .A(n40), .B(n9), .C(n1), .D(n25), .Z(rdata[28]) );
  HS65_LS_IVX9 U71 ( .A(rdata1[12]), .Z(n25) );
  HS65_LS_OAI22X6 U72 ( .A(n40), .B(n8), .C(n1), .D(n24), .Z(rdata[29]) );
  HS65_LS_IVX9 U73 ( .A(rdata1[13]), .Z(n24) );
  HS65_LS_OAI22X6 U74 ( .A(n40), .B(n7), .C(n1), .D(n23), .Z(rdata[30]) );
  HS65_LS_IVX9 U75 ( .A(rdata1[14]), .Z(n23) );
  HS65_LS_OAI22X6 U76 ( .A(n40), .B(n6), .C(n1), .D(n22), .Z(rdata[31]) );
  HS65_LS_IVX9 U77 ( .A(rdata1[15]), .Z(n22) );
  HS65_LS_OAI22X6 U78 ( .A(n40), .B(n21), .C(n1), .D(n41), .Z(rdata[16]) );
  HS65_LS_IVX9 U79 ( .A(rdata1[0]), .Z(n41) );
  HS65_LS_NOR2AX3 U80 ( .A(rdata0[0]), .B(n3), .Z(rdata[48]) );
  HS65_LS_IVX9 U81 ( .A(rdata1[20]), .Z(n17) );
  HS65_LS_IVX9 U82 ( .A(rdata1[21]), .Z(n16) );
  HS65_LS_IVX9 U83 ( .A(rdata1[22]), .Z(n15) );
  HS65_LS_IVX9 U84 ( .A(rdata1[23]), .Z(n14) );
  HS65_LS_IVX9 U85 ( .A(rdata1[24]), .Z(n13) );
  HS65_LS_IVX9 U86 ( .A(rdata1[25]), .Z(n12) );
  HS65_LS_IVX9 U87 ( .A(rdata1[26]), .Z(n11) );
  HS65_LS_IVX9 U88 ( .A(rdata1[27]), .Z(n10) );
  HS65_LS_IVX9 U89 ( .A(rdata1[28]), .Z(n9) );
  HS65_LS_IVX9 U90 ( .A(rdata1[29]), .Z(n8) );
  HS65_LS_IVX9 U91 ( .A(rdata1[30]), .Z(n7) );
  HS65_LS_IVX9 U92 ( .A(rdata1[31]), .Z(n6) );
  HS65_LS_IVX9 U93 ( .A(rdata1[16]), .Z(n21) );
  HS65_LS_AO222X4 U94 ( .A(rdata0[0]), .B(n37), .C(rdata1[0]), .D(n42), .E(
        rdata2[0]), .F(n38), .Z(rdata[0]) );
  HS65_LS_AO222X4 U95 ( .A(rdata0[1]), .B(n37), .C(rdata1[1]), .D(n42), .E(
        rdata2[1]), .F(n38), .Z(rdata[1]) );
  HS65_LS_AO222X4 U96 ( .A(rdata0[2]), .B(n37), .C(rdata1[2]), .D(n42), .E(
        rdata2[2]), .F(n38), .Z(rdata[2]) );
  HS65_LS_AO222X4 U97 ( .A(rdata0[3]), .B(n37), .C(rdata1[3]), .D(n42), .E(
        rdata2[3]), .F(n38), .Z(rdata[3]) );
  HS65_LS_AO222X4 U98 ( .A(rdata0[4]), .B(n37), .C(rdata1[4]), .D(n42), .E(
        rdata2[4]), .F(n38), .Z(rdata[4]) );
  HS65_LS_AO222X4 U99 ( .A(rdata0[5]), .B(n37), .C(rdata1[5]), .D(n42), .E(
        rdata2[5]), .F(n38), .Z(rdata[5]) );
  HS65_LS_AO222X4 U100 ( .A(rdata0[6]), .B(n37), .C(rdata1[6]), .D(n42), .E(
        rdata2[6]), .F(n38), .Z(rdata[6]) );
  HS65_LS_AO222X4 U101 ( .A(rdata0[7]), .B(n37), .C(rdata1[7]), .D(n42), .E(
        rdata2[7]), .F(n38), .Z(rdata[7]) );
  HS65_LS_AO222X4 U102 ( .A(rdata0[8]), .B(n37), .C(rdata1[8]), .D(n42), .E(
        rdata2[8]), .F(n38), .Z(rdata[8]) );
  HS65_LS_AO222X4 U103 ( .A(rdata0[9]), .B(n37), .C(rdata1[9]), .D(n42), .E(
        rdata2[9]), .F(n38), .Z(rdata[9]) );
  HS65_LS_AO222X4 U104 ( .A(rdata0[10]), .B(n37), .C(rdata1[10]), .D(n42), .E(
        rdata2[10]), .F(n38), .Z(rdata[10]) );
  HS65_LS_AO222X4 U105 ( .A(rdata0[11]), .B(n37), .C(rdata1[11]), .D(n42), .E(
        rdata2[11]), .F(n38), .Z(rdata[11]) );
  HS65_LS_AO222X4 U106 ( .A(rdata0[12]), .B(n37), .C(rdata1[12]), .D(n42), .E(
        rdata2[12]), .F(n38), .Z(rdata[12]) );
  HS65_LS_AO222X4 U107 ( .A(rdata0[13]), .B(n37), .C(rdata1[13]), .D(n42), .E(
        rdata2[13]), .F(n38), .Z(rdata[13]) );
  HS65_LS_AO222X4 U108 ( .A(rdata0[14]), .B(n37), .C(rdata1[14]), .D(n42), .E(
        rdata2[14]), .F(n38), .Z(rdata[14]) );
  HS65_LS_AO222X4 U109 ( .A(rdata0[15]), .B(n37), .C(rdata1[15]), .D(n42), .E(
        rdata2[15]), .F(n38), .Z(rdata[15]) );
  HS65_LS_NOR2AX3 U110 ( .A(rdata0[13]), .B(n4), .Z(rdata[61]) );
endmodule


module bram_DATA5_ADDR3_0 ( clk, reset, rd_addr, wr_addr, wr_data, wr_ena, 
        rd_data );
  input [2:0] rd_addr;
  input [2:0] wr_addr;
  input [4:0] wr_data;
  output [4:0] rd_data;
  input clk, reset, wr_ena;
  wire   \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N34,
         N35, N36, N37, N38, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n1, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n117, n118,
         n119, n120;

  HS65_LS_DFPRQX9 \mem_reg[5][4]  ( .D(n106), .CP(clk), .RN(n1), .Q(
        \mem[5][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[5][3]  ( .D(n105), .CP(clk), .RN(n1), .Q(
        \mem[5][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[5][2]  ( .D(n104), .CP(clk), .RN(n1), .Q(
        \mem[5][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[5][1]  ( .D(n103), .CP(clk), .RN(n1), .Q(
        \mem[5][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[5][0]  ( .D(n102), .CP(clk), .RN(n22), .Q(
        \mem[5][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[4][4]  ( .D(n101), .CP(clk), .RN(n22), .Q(
        \mem[4][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[4][3]  ( .D(n100), .CP(clk), .RN(n22), .Q(
        \mem[4][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[4][2]  ( .D(n99), .CP(clk), .RN(n22), .Q(
        \mem[4][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[4][1]  ( .D(n98), .CP(clk), .RN(n22), .Q(
        \mem[4][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[4][0]  ( .D(n97), .CP(clk), .RN(n22), .Q(
        \mem[4][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][4]  ( .D(n86), .CP(clk), .RN(n22), .Q(
        \mem[1][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][3]  ( .D(n85), .CP(clk), .RN(n22), .Q(
        \mem[1][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][2]  ( .D(n84), .CP(clk), .RN(n22), .Q(
        \mem[1][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][1]  ( .D(n83), .CP(clk), .RN(n22), .Q(
        \mem[1][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][0]  ( .D(n82), .CP(clk), .RN(n22), .Q(
        \mem[1][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][4]  ( .D(n81), .CP(clk), .RN(n22), .Q(
        \mem[0][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][3]  ( .D(n80), .CP(clk), .RN(n1), .Q(\mem[0][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][2]  ( .D(n79), .CP(clk), .RN(n1), .Q(\mem[0][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][1]  ( .D(n78), .CP(clk), .RN(n1), .Q(\mem[0][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][0]  ( .D(n77), .CP(clk), .RN(n1), .Q(\mem[0][0] ) );
  HS65_LS_DFPRQX9 \rd_data_reg[4]  ( .D(N34), .CP(clk), .RN(n1), .Q(rd_data[4]) );
  HS65_LS_DFPRQX9 \rd_data_reg[3]  ( .D(N35), .CP(clk), .RN(n1), .Q(rd_data[3]) );
  HS65_LS_DFPRQX9 \rd_data_reg[2]  ( .D(N36), .CP(clk), .RN(n1), .Q(rd_data[2]) );
  HS65_LS_DFPRQX9 \rd_data_reg[1]  ( .D(N37), .CP(clk), .RN(n1), .Q(rd_data[1]) );
  HS65_LS_DFPRQX9 \rd_data_reg[0]  ( .D(N38), .CP(clk), .RN(n1), .Q(rd_data[0]) );
  HS65_LS_DFPRQNX9 \mem_reg[7][4]  ( .D(n116), .CP(clk), .RN(n23), .QN(n2) );
  HS65_LS_DFPRQNX9 \mem_reg[7][3]  ( .D(n115), .CP(clk), .RN(n22), .QN(n3) );
  HS65_LS_DFPRQNX9 \mem_reg[7][2]  ( .D(n114), .CP(clk), .RN(n24), .QN(n4) );
  HS65_LS_DFPRQNX9 \mem_reg[7][1]  ( .D(n113), .CP(clk), .RN(n24), .QN(n5) );
  HS65_LS_DFPRQNX9 \mem_reg[7][0]  ( .D(n112), .CP(clk), .RN(n24), .QN(n6) );
  HS65_LS_DFPRQNX9 \mem_reg[3][4]  ( .D(n96), .CP(clk), .RN(n23), .QN(n12) );
  HS65_LS_DFPRQNX9 \mem_reg[3][3]  ( .D(n95), .CP(clk), .RN(n23), .QN(n13) );
  HS65_LS_DFPRQNX9 \mem_reg[3][2]  ( .D(n94), .CP(clk), .RN(n23), .QN(n14) );
  HS65_LS_DFPRQNX9 \mem_reg[3][1]  ( .D(n93), .CP(clk), .RN(n23), .QN(n15) );
  HS65_LS_DFPRQNX9 \mem_reg[3][0]  ( .D(n92), .CP(clk), .RN(n23), .QN(n16) );
  HS65_LS_DFPRQNX9 \mem_reg[6][4]  ( .D(n111), .CP(clk), .RN(n24), .QN(n7) );
  HS65_LS_DFPRQNX9 \mem_reg[6][3]  ( .D(n110), .CP(clk), .RN(n24), .QN(n8) );
  HS65_LS_DFPRQNX9 \mem_reg[6][2]  ( .D(n109), .CP(clk), .RN(n23), .QN(n9) );
  HS65_LS_DFPRQNX9 \mem_reg[6][1]  ( .D(n108), .CP(clk), .RN(n23), .QN(n10) );
  HS65_LS_DFPRQNX9 \mem_reg[6][0]  ( .D(n107), .CP(clk), .RN(n23), .QN(n11) );
  HS65_LS_DFPRQNX9 \mem_reg[2][4]  ( .D(n91), .CP(clk), .RN(n23), .QN(n17) );
  HS65_LS_DFPRQNX9 \mem_reg[2][3]  ( .D(n90), .CP(clk), .RN(n23), .QN(n18) );
  HS65_LS_DFPRQNX9 \mem_reg[2][2]  ( .D(n89), .CP(clk), .RN(n23), .QN(n19) );
  HS65_LS_DFPRQNX9 \mem_reg[2][1]  ( .D(n88), .CP(clk), .RN(n23), .QN(n20) );
  HS65_LS_DFPRQNX9 \mem_reg[2][0]  ( .D(n87), .CP(clk), .RN(n23), .QN(n21) );
  HS65_LS_BFX9 U3 ( .A(n25), .Z(n1) );
  HS65_LS_BFX9 U4 ( .A(n25), .Z(n22) );
  HS65_LS_BFX9 U5 ( .A(n25), .Z(n23) );
  HS65_LS_BFX9 U6 ( .A(n25), .Z(n24) );
  HS65_LS_IVX9 U7 ( .A(reset), .Z(n25) );
  HS65_LS_IVX9 U8 ( .A(n39), .Z(n35) );
  HS65_LS_IVX9 U9 ( .A(n44), .Z(n31) );
  HS65_LS_IVX9 U10 ( .A(n43), .Z(n32) );
  HS65_LS_IVX9 U11 ( .A(n47), .Z(n29) );
  HS65_LS_IVX9 U12 ( .A(n48), .Z(n28) );
  HS65_LS_IVX9 U13 ( .A(n42), .Z(n33) );
  HS65_LS_NAND3X5 U14 ( .A(n37), .B(n36), .C(n40), .Z(n39) );
  HS65_LS_NAND3X5 U15 ( .A(n37), .B(n36), .C(n45), .Z(n44) );
  HS65_LS_IVX9 U16 ( .A(n46), .Z(n30) );
  HS65_LS_IVX9 U17 ( .A(n41), .Z(n34) );
  HS65_LS_NOR3X4 U18 ( .A(n26), .B(rd_addr[1]), .C(n27), .Z(n51) );
  HS65_LS_NOR3X4 U19 ( .A(rd_addr[1]), .B(rd_addr[2]), .C(n26), .Z(n56) );
  HS65_LS_NOR3X4 U20 ( .A(rd_addr[1]), .B(rd_addr[2]), .C(rd_addr[0]), .Z(n57)
         );
  HS65_LS_NOR3X4 U21 ( .A(rd_addr[0]), .B(rd_addr[1]), .C(n27), .Z(n52) );
  HS65_LS_NAND3X5 U22 ( .A(n26), .B(n27), .C(rd_addr[1]), .Z(n59) );
  HS65_LS_NAND3X5 U23 ( .A(rd_addr[0]), .B(n27), .C(rd_addr[1]), .Z(n60) );
  HS65_LS_NAND3X5 U24 ( .A(rd_addr[1]), .B(n26), .C(rd_addr[2]), .Z(n54) );
  HS65_LS_NAND3X5 U25 ( .A(rd_addr[1]), .B(rd_addr[0]), .C(rd_addr[2]), .Z(n55) );
  HS65_LS_OAI22X6 U26 ( .A(n21), .B(n59), .C(n16), .D(n60), .Z(n58) );
  HS65_LS_OAI22X6 U27 ( .A(n20), .B(n59), .C(n15), .D(n60), .Z(n64) );
  HS65_LS_OAI22X6 U28 ( .A(n19), .B(n59), .C(n14), .D(n60), .Z(n68) );
  HS65_LS_OAI22X6 U29 ( .A(n18), .B(n59), .C(n13), .D(n60), .Z(n72) );
  HS65_LS_OAI22X6 U30 ( .A(n17), .B(n59), .C(n12), .D(n60), .Z(n76) );
  HS65_LS_IVX9 U31 ( .A(rd_addr[0]), .Z(n26) );
  HS65_LS_IVX9 U32 ( .A(rd_addr[2]), .Z(n27) );
  HS65_LS_OAI22X6 U33 ( .A(n120), .B(n43), .C(n32), .D(n16), .Z(n92) );
  HS65_LS_OAI22X6 U34 ( .A(n119), .B(n43), .C(n32), .D(n15), .Z(n93) );
  HS65_LS_OAI22X6 U35 ( .A(n118), .B(n43), .C(n32), .D(n14), .Z(n94) );
  HS65_LS_OAI22X6 U36 ( .A(n117), .B(n43), .C(n32), .D(n13), .Z(n95) );
  HS65_LS_OAI22X6 U37 ( .A(n38), .B(n43), .C(n32), .D(n12), .Z(n96) );
  HS65_LS_OAI22X6 U38 ( .A(n120), .B(n47), .C(n29), .D(n11), .Z(n107) );
  HS65_LS_OAI22X6 U39 ( .A(n119), .B(n47), .C(n29), .D(n10), .Z(n108) );
  HS65_LS_OAI22X6 U40 ( .A(n118), .B(n47), .C(n29), .D(n9), .Z(n109) );
  HS65_LS_OAI22X6 U41 ( .A(n117), .B(n47), .C(n29), .D(n8), .Z(n110) );
  HS65_LS_OAI22X6 U42 ( .A(n38), .B(n47), .C(n29), .D(n7), .Z(n111) );
  HS65_LS_OAI22X6 U43 ( .A(n120), .B(n48), .C(n28), .D(n6), .Z(n112) );
  HS65_LS_OAI22X6 U44 ( .A(n119), .B(n48), .C(n28), .D(n5), .Z(n113) );
  HS65_LS_OAI22X6 U45 ( .A(n118), .B(n48), .C(n28), .D(n4), .Z(n114) );
  HS65_LS_OAI22X6 U46 ( .A(n117), .B(n48), .C(n28), .D(n3), .Z(n115) );
  HS65_LS_OAI22X6 U47 ( .A(n38), .B(n48), .C(n28), .D(n2), .Z(n116) );
  HS65_LS_OAI22X6 U48 ( .A(n120), .B(n42), .C(n33), .D(n21), .Z(n87) );
  HS65_LS_OAI22X6 U49 ( .A(n119), .B(n42), .C(n33), .D(n20), .Z(n88) );
  HS65_LS_OAI22X6 U50 ( .A(n118), .B(n42), .C(n33), .D(n19), .Z(n89) );
  HS65_LS_OAI22X6 U51 ( .A(n117), .B(n42), .C(n33), .D(n18), .Z(n90) );
  HS65_LS_OAI22X6 U52 ( .A(n38), .B(n42), .C(n33), .D(n17), .Z(n91) );
  HS65_LS_NAND2X7 U53 ( .A(n49), .B(n50), .Z(N38) );
  HS65_LS_AOI212X4 U54 ( .A(n51), .B(\mem[5][0] ), .C(n52), .D(\mem[4][0] ), 
        .E(n53), .Z(n50) );
  HS65_LS_AOI212X4 U55 ( .A(n56), .B(\mem[1][0] ), .C(n57), .D(\mem[0][0] ), 
        .E(n58), .Z(n49) );
  HS65_LS_OAI22X6 U56 ( .A(n11), .B(n54), .C(n6), .D(n55), .Z(n53) );
  HS65_LS_NAND2X7 U57 ( .A(n61), .B(n62), .Z(N37) );
  HS65_LS_AOI212X4 U58 ( .A(n51), .B(\mem[5][1] ), .C(n52), .D(\mem[4][1] ), 
        .E(n63), .Z(n62) );
  HS65_LS_AOI212X4 U59 ( .A(n56), .B(\mem[1][1] ), .C(n57), .D(\mem[0][1] ), 
        .E(n64), .Z(n61) );
  HS65_LS_OAI22X6 U60 ( .A(n10), .B(n54), .C(n5), .D(n55), .Z(n63) );
  HS65_LS_NAND2X7 U61 ( .A(n65), .B(n66), .Z(N36) );
  HS65_LS_AOI212X4 U62 ( .A(n51), .B(\mem[5][2] ), .C(n52), .D(\mem[4][2] ), 
        .E(n67), .Z(n66) );
  HS65_LS_AOI212X4 U63 ( .A(n56), .B(\mem[1][2] ), .C(n57), .D(\mem[0][2] ), 
        .E(n68), .Z(n65) );
  HS65_LS_OAI22X6 U64 ( .A(n9), .B(n54), .C(n4), .D(n55), .Z(n67) );
  HS65_LS_NAND2X7 U65 ( .A(n69), .B(n70), .Z(N35) );
  HS65_LS_AOI212X4 U66 ( .A(n51), .B(\mem[5][3] ), .C(n52), .D(\mem[4][3] ), 
        .E(n71), .Z(n70) );
  HS65_LS_AOI212X4 U67 ( .A(n56), .B(\mem[1][3] ), .C(n57), .D(\mem[0][3] ), 
        .E(n72), .Z(n69) );
  HS65_LS_OAI22X6 U68 ( .A(n8), .B(n54), .C(n3), .D(n55), .Z(n71) );
  HS65_LS_NAND2X7 U69 ( .A(n73), .B(n74), .Z(N34) );
  HS65_LS_AOI212X4 U70 ( .A(n51), .B(\mem[5][4] ), .C(n52), .D(\mem[4][4] ), 
        .E(n75), .Z(n74) );
  HS65_LS_AOI212X4 U71 ( .A(n56), .B(\mem[1][4] ), .C(n57), .D(\mem[0][4] ), 
        .E(n76), .Z(n73) );
  HS65_LS_OAI22X6 U72 ( .A(n7), .B(n54), .C(n2), .D(n55), .Z(n75) );
  HS65_LS_AO22X9 U73 ( .A(n35), .B(wr_data[0]), .C(n39), .D(\mem[0][0] ), .Z(
        n77) );
  HS65_LS_AO22X9 U74 ( .A(n35), .B(wr_data[1]), .C(n39), .D(\mem[0][1] ), .Z(
        n78) );
  HS65_LS_AO22X9 U75 ( .A(n35), .B(wr_data[2]), .C(n39), .D(\mem[0][2] ), .Z(
        n79) );
  HS65_LS_AO22X9 U76 ( .A(n35), .B(wr_data[3]), .C(n39), .D(\mem[0][3] ), .Z(
        n80) );
  HS65_LS_AO22X9 U77 ( .A(n35), .B(wr_data[4]), .C(n39), .D(\mem[0][4] ), .Z(
        n81) );
  HS65_LS_AO22X9 U78 ( .A(wr_data[0]), .B(n31), .C(n44), .D(\mem[4][0] ), .Z(
        n97) );
  HS65_LS_AO22X9 U79 ( .A(wr_data[1]), .B(n31), .C(n44), .D(\mem[4][1] ), .Z(
        n98) );
  HS65_LS_AO22X9 U80 ( .A(wr_data[2]), .B(n31), .C(n44), .D(\mem[4][2] ), .Z(
        n99) );
  HS65_LS_AO22X9 U81 ( .A(wr_data[3]), .B(n31), .C(n44), .D(\mem[4][3] ), .Z(
        n100) );
  HS65_LS_AO22X9 U82 ( .A(wr_data[4]), .B(n31), .C(n44), .D(\mem[4][4] ), .Z(
        n101) );
  HS65_LS_AO22X9 U83 ( .A(wr_data[0]), .B(n30), .C(n46), .D(\mem[5][0] ), .Z(
        n102) );
  HS65_LS_AO22X9 U84 ( .A(wr_data[1]), .B(n30), .C(n46), .D(\mem[5][1] ), .Z(
        n103) );
  HS65_LS_AO22X9 U85 ( .A(wr_data[2]), .B(n30), .C(n46), .D(\mem[5][2] ), .Z(
        n104) );
  HS65_LS_AO22X9 U86 ( .A(wr_data[3]), .B(n30), .C(n46), .D(\mem[5][3] ), .Z(
        n105) );
  HS65_LS_AO22X9 U87 ( .A(wr_data[4]), .B(n30), .C(n46), .D(\mem[5][4] ), .Z(
        n106) );
  HS65_LS_AO22X9 U88 ( .A(wr_data[0]), .B(n34), .C(n41), .D(\mem[1][0] ), .Z(
        n82) );
  HS65_LS_AO22X9 U89 ( .A(wr_data[1]), .B(n34), .C(n41), .D(\mem[1][1] ), .Z(
        n83) );
  HS65_LS_AO22X9 U90 ( .A(wr_data[2]), .B(n34), .C(n41), .D(\mem[1][2] ), .Z(
        n84) );
  HS65_LS_AO22X9 U91 ( .A(wr_data[3]), .B(n34), .C(n41), .D(\mem[1][3] ), .Z(
        n85) );
  HS65_LS_AO22X9 U92 ( .A(wr_data[4]), .B(n34), .C(n41), .D(\mem[1][4] ), .Z(
        n86) );
  HS65_LS_NAND3X5 U93 ( .A(wr_addr[0]), .B(n40), .C(wr_addr[1]), .Z(n43) );
  HS65_LS_NAND3X5 U94 ( .A(wr_addr[1]), .B(n37), .C(n45), .Z(n47) );
  HS65_LS_NAND3X5 U95 ( .A(wr_addr[1]), .B(wr_addr[0]), .C(n45), .Z(n48) );
  HS65_LS_NAND3X5 U96 ( .A(n40), .B(n37), .C(wr_addr[1]), .Z(n42) );
  HS65_LS_NOR2AX3 U97 ( .A(wr_ena), .B(wr_addr[2]), .Z(n40) );
  HS65_LS_NAND3X5 U98 ( .A(wr_addr[0]), .B(n36), .C(n45), .Z(n46) );
  HS65_LS_NAND3X5 U99 ( .A(n40), .B(n36), .C(wr_addr[0]), .Z(n41) );
  HS65_LS_IVX9 U100 ( .A(wr_addr[0]), .Z(n37) );
  HS65_LS_IVX9 U101 ( .A(wr_data[0]), .Z(n120) );
  HS65_LS_IVX9 U102 ( .A(wr_data[1]), .Z(n119) );
  HS65_LS_IVX9 U103 ( .A(wr_data[2]), .Z(n118) );
  HS65_LS_IVX9 U104 ( .A(wr_data[3]), .Z(n117) );
  HS65_LS_IVX9 U105 ( .A(wr_data[4]), .Z(n38) );
  HS65_LS_IVX9 U106 ( .A(wr_addr[1]), .Z(n36) );
  HS65_LS_AND2X4 U107 ( .A(wr_addr[2]), .B(wr_ena), .Z(n45) );
endmodule


module nAdapter_0 ( na_clk, na_reset, .proc_in({\proc_in[MCMD][1] , 
        \proc_in[MCMD][0] , \proc_in[MADDR][31] , \proc_in[MADDR][30] , 
        \proc_in[MADDR][29] , \proc_in[MADDR][28] , \proc_in[MADDR][27] , 
        \proc_in[MADDR][26] , \proc_in[MADDR][25] , \proc_in[MADDR][24] , 
        \proc_in[MADDR][23] , \proc_in[MADDR][22] , \proc_in[MADDR][21] , 
        \proc_in[MADDR][20] , \proc_in[MADDR][19] , \proc_in[MADDR][18] , 
        \proc_in[MADDR][17] , \proc_in[MADDR][16] , \proc_in[MADDR][15] , 
        \proc_in[MADDR][14] , \proc_in[MADDR][13] , \proc_in[MADDR][12] , 
        \proc_in[MADDR][11] , \proc_in[MADDR][10] , \proc_in[MADDR][9] , 
        \proc_in[MADDR][8] , \proc_in[MADDR][7] , \proc_in[MADDR][6] , 
        \proc_in[MADDR][5] , \proc_in[MADDR][4] , \proc_in[MADDR][3] , 
        \proc_in[MADDR][2] , \proc_in[MADDR][1] , \proc_in[MADDR][0] , 
        \proc_in[MDATA][31] , \proc_in[MDATA][30] , \proc_in[MDATA][29] , 
        \proc_in[MDATA][28] , \proc_in[MDATA][27] , \proc_in[MDATA][26] , 
        \proc_in[MDATA][25] , \proc_in[MDATA][24] , \proc_in[MDATA][23] , 
        \proc_in[MDATA][22] , \proc_in[MDATA][21] , \proc_in[MDATA][20] , 
        \proc_in[MDATA][19] , \proc_in[MDATA][18] , \proc_in[MDATA][17] , 
        \proc_in[MDATA][16] , \proc_in[MDATA][15] , \proc_in[MDATA][14] , 
        \proc_in[MDATA][13] , \proc_in[MDATA][12] , \proc_in[MDATA][11] , 
        \proc_in[MDATA][10] , \proc_in[MDATA][9] , \proc_in[MDATA][8] , 
        \proc_in[MDATA][7] , \proc_in[MDATA][6] , \proc_in[MDATA][5] , 
        \proc_in[MDATA][4] , \proc_in[MDATA][3] , \proc_in[MDATA][2] , 
        \proc_in[MDATA][1] , \proc_in[MDATA][0] }), .proc_out({
        \proc_out[SCMDACCEPT] , \proc_out[SRESP] , \proc_out[SDATA][31] , 
        \proc_out[SDATA][30] , \proc_out[SDATA][29] , \proc_out[SDATA][28] , 
        \proc_out[SDATA][27] , \proc_out[SDATA][26] , \proc_out[SDATA][25] , 
        \proc_out[SDATA][24] , \proc_out[SDATA][23] , \proc_out[SDATA][22] , 
        \proc_out[SDATA][21] , \proc_out[SDATA][20] , \proc_out[SDATA][19] , 
        \proc_out[SDATA][18] , \proc_out[SDATA][17] , \proc_out[SDATA][16] , 
        \proc_out[SDATA][15] , \proc_out[SDATA][14] , \proc_out[SDATA][13] , 
        \proc_out[SDATA][12] , \proc_out[SDATA][11] , \proc_out[SDATA][10] , 
        \proc_out[SDATA][9] , \proc_out[SDATA][8] , \proc_out[SDATA][7] , 
        \proc_out[SDATA][6] , \proc_out[SDATA][5] , \proc_out[SDATA][4] , 
        \proc_out[SDATA][3] , \proc_out[SDATA][2] , \proc_out[SDATA][1] , 
        \proc_out[SDATA][0] }), .spm_in({\spm_in[SCMDACCEPT] , \spm_in[SRESP] , 
        \spm_in[SDATA][63] , \spm_in[SDATA][62] , \spm_in[SDATA][61] , 
        \spm_in[SDATA][60] , \spm_in[SDATA][59] , \spm_in[SDATA][58] , 
        \spm_in[SDATA][57] , \spm_in[SDATA][56] , \spm_in[SDATA][55] , 
        \spm_in[SDATA][54] , \spm_in[SDATA][53] , \spm_in[SDATA][52] , 
        \spm_in[SDATA][51] , \spm_in[SDATA][50] , \spm_in[SDATA][49] , 
        \spm_in[SDATA][48] , \spm_in[SDATA][47] , \spm_in[SDATA][46] , 
        \spm_in[SDATA][45] , \spm_in[SDATA][44] , \spm_in[SDATA][43] , 
        \spm_in[SDATA][42] , \spm_in[SDATA][41] , \spm_in[SDATA][40] , 
        \spm_in[SDATA][39] , \spm_in[SDATA][38] , \spm_in[SDATA][37] , 
        \spm_in[SDATA][36] , \spm_in[SDATA][35] , \spm_in[SDATA][34] , 
        \spm_in[SDATA][33] , \spm_in[SDATA][32] , \spm_in[SDATA][31] , 
        \spm_in[SDATA][30] , \spm_in[SDATA][29] , \spm_in[SDATA][28] , 
        \spm_in[SDATA][27] , \spm_in[SDATA][26] , \spm_in[SDATA][25] , 
        \spm_in[SDATA][24] , \spm_in[SDATA][23] , \spm_in[SDATA][22] , 
        \spm_in[SDATA][21] , \spm_in[SDATA][20] , \spm_in[SDATA][19] , 
        \spm_in[SDATA][18] , \spm_in[SDATA][17] , \spm_in[SDATA][16] , 
        \spm_in[SDATA][15] , \spm_in[SDATA][14] , \spm_in[SDATA][13] , 
        \spm_in[SDATA][12] , \spm_in[SDATA][11] , \spm_in[SDATA][10] , 
        \spm_in[SDATA][9] , \spm_in[SDATA][8] , \spm_in[SDATA][7] , 
        \spm_in[SDATA][6] , \spm_in[SDATA][5] , \spm_in[SDATA][4] , 
        \spm_in[SDATA][3] , \spm_in[SDATA][2] , \spm_in[SDATA][1] , 
        \spm_in[SDATA][0] }), .spm_out({\spm_out[MCMD][1] , \spm_out[MCMD][0] , 
        \spm_out[MADDR][31] , \spm_out[MADDR][30] , \spm_out[MADDR][29] , 
        \spm_out[MADDR][28] , \spm_out[MADDR][27] , \spm_out[MADDR][26] , 
        \spm_out[MADDR][25] , \spm_out[MADDR][24] , \spm_out[MADDR][23] , 
        \spm_out[MADDR][22] , \spm_out[MADDR][21] , \spm_out[MADDR][20] , 
        \spm_out[MADDR][19] , \spm_out[MADDR][18] , \spm_out[MADDR][17] , 
        \spm_out[MADDR][16] , \spm_out[MADDR][15] , \spm_out[MADDR][14] , 
        \spm_out[MADDR][13] , \spm_out[MADDR][12] , \spm_out[MADDR][11] , 
        \spm_out[MADDR][10] , \spm_out[MADDR][9] , \spm_out[MADDR][8] , 
        \spm_out[MADDR][7] , \spm_out[MADDR][6] , \spm_out[MADDR][5] , 
        \spm_out[MADDR][4] , \spm_out[MADDR][3] , \spm_out[MADDR][2] , 
        \spm_out[MADDR][1] , \spm_out[MADDR][0] , \spm_out[MDATA][63] , 
        \spm_out[MDATA][62] , \spm_out[MDATA][61] , \spm_out[MDATA][60] , 
        \spm_out[MDATA][59] , \spm_out[MDATA][58] , \spm_out[MDATA][57] , 
        \spm_out[MDATA][56] , \spm_out[MDATA][55] , \spm_out[MDATA][54] , 
        \spm_out[MDATA][53] , \spm_out[MDATA][52] , \spm_out[MDATA][51] , 
        \spm_out[MDATA][50] , \spm_out[MDATA][49] , \spm_out[MDATA][48] , 
        \spm_out[MDATA][47] , \spm_out[MDATA][46] , \spm_out[MDATA][45] , 
        \spm_out[MDATA][44] , \spm_out[MDATA][43] , \spm_out[MDATA][42] , 
        \spm_out[MDATA][41] , \spm_out[MDATA][40] , \spm_out[MDATA][39] , 
        \spm_out[MDATA][38] , \spm_out[MDATA][37] , \spm_out[MDATA][36] , 
        \spm_out[MDATA][35] , \spm_out[MDATA][34] , \spm_out[MDATA][33] , 
        \spm_out[MDATA][32] , \spm_out[MDATA][31] , \spm_out[MDATA][30] , 
        \spm_out[MDATA][29] , \spm_out[MDATA][28] , \spm_out[MDATA][27] , 
        \spm_out[MDATA][26] , \spm_out[MDATA][25] , \spm_out[MDATA][24] , 
        \spm_out[MDATA][23] , \spm_out[MDATA][22] , \spm_out[MDATA][21] , 
        \spm_out[MDATA][20] , \spm_out[MDATA][19] , \spm_out[MDATA][18] , 
        \spm_out[MDATA][17] , \spm_out[MDATA][16] , \spm_out[MDATA][15] , 
        \spm_out[MDATA][14] , \spm_out[MDATA][13] , \spm_out[MDATA][12] , 
        \spm_out[MDATA][11] , \spm_out[MDATA][10] , \spm_out[MDATA][9] , 
        \spm_out[MDATA][8] , \spm_out[MDATA][7] , \spm_out[MDATA][6] , 
        \spm_out[MDATA][5] , \spm_out[MDATA][4] , \spm_out[MDATA][3] , 
        \spm_out[MDATA][2] , \spm_out[MDATA][1] , \spm_out[MDATA][0] }), 
        pkt_in, pkt_out );
  input [34:0] pkt_in;
  output [34:0] pkt_out;
  input na_clk, na_reset, \proc_in[MCMD][1] , \proc_in[MCMD][0] ,
         \proc_in[MADDR][31] , \proc_in[MADDR][30] , \proc_in[MADDR][29] ,
         \proc_in[MADDR][28] , \proc_in[MADDR][27] , \proc_in[MADDR][26] ,
         \proc_in[MADDR][25] , \proc_in[MADDR][24] , \proc_in[MADDR][23] ,
         \proc_in[MADDR][22] , \proc_in[MADDR][21] , \proc_in[MADDR][20] ,
         \proc_in[MADDR][19] , \proc_in[MADDR][18] , \proc_in[MADDR][17] ,
         \proc_in[MADDR][16] , \proc_in[MADDR][15] , \proc_in[MADDR][14] ,
         \proc_in[MADDR][13] , \proc_in[MADDR][12] , \proc_in[MADDR][11] ,
         \proc_in[MADDR][10] , \proc_in[MADDR][9] , \proc_in[MADDR][8] ,
         \proc_in[MADDR][7] , \proc_in[MADDR][6] , \proc_in[MADDR][5] ,
         \proc_in[MADDR][4] , \proc_in[MADDR][3] , \proc_in[MADDR][2] ,
         \proc_in[MADDR][1] , \proc_in[MADDR][0] , \proc_in[MDATA][31] ,
         \proc_in[MDATA][30] , \proc_in[MDATA][29] , \proc_in[MDATA][28] ,
         \proc_in[MDATA][27] , \proc_in[MDATA][26] , \proc_in[MDATA][25] ,
         \proc_in[MDATA][24] , \proc_in[MDATA][23] , \proc_in[MDATA][22] ,
         \proc_in[MDATA][21] , \proc_in[MDATA][20] , \proc_in[MDATA][19] ,
         \proc_in[MDATA][18] , \proc_in[MDATA][17] , \proc_in[MDATA][16] ,
         \proc_in[MDATA][15] , \proc_in[MDATA][14] , \proc_in[MDATA][13] ,
         \proc_in[MDATA][12] , \proc_in[MDATA][11] , \proc_in[MDATA][10] ,
         \proc_in[MDATA][9] , \proc_in[MDATA][8] , \proc_in[MDATA][7] ,
         \proc_in[MDATA][6] , \proc_in[MDATA][5] , \proc_in[MDATA][4] ,
         \proc_in[MDATA][3] , \proc_in[MDATA][2] , \proc_in[MDATA][1] ,
         \proc_in[MDATA][0] , \spm_in[SCMDACCEPT] , \spm_in[SRESP] ,
         \spm_in[SDATA][63] , \spm_in[SDATA][62] , \spm_in[SDATA][61] ,
         \spm_in[SDATA][60] , \spm_in[SDATA][59] , \spm_in[SDATA][58] ,
         \spm_in[SDATA][57] , \spm_in[SDATA][56] , \spm_in[SDATA][55] ,
         \spm_in[SDATA][54] , \spm_in[SDATA][53] , \spm_in[SDATA][52] ,
         \spm_in[SDATA][51] , \spm_in[SDATA][50] , \spm_in[SDATA][49] ,
         \spm_in[SDATA][48] , \spm_in[SDATA][47] , \spm_in[SDATA][46] ,
         \spm_in[SDATA][45] , \spm_in[SDATA][44] , \spm_in[SDATA][43] ,
         \spm_in[SDATA][42] , \spm_in[SDATA][41] , \spm_in[SDATA][40] ,
         \spm_in[SDATA][39] , \spm_in[SDATA][38] , \spm_in[SDATA][37] ,
         \spm_in[SDATA][36] , \spm_in[SDATA][35] , \spm_in[SDATA][34] ,
         \spm_in[SDATA][33] , \spm_in[SDATA][32] , \spm_in[SDATA][31] ,
         \spm_in[SDATA][30] , \spm_in[SDATA][29] , \spm_in[SDATA][28] ,
         \spm_in[SDATA][27] , \spm_in[SDATA][26] , \spm_in[SDATA][25] ,
         \spm_in[SDATA][24] , \spm_in[SDATA][23] , \spm_in[SDATA][22] ,
         \spm_in[SDATA][21] , \spm_in[SDATA][20] , \spm_in[SDATA][19] ,
         \spm_in[SDATA][18] , \spm_in[SDATA][17] , \spm_in[SDATA][16] ,
         \spm_in[SDATA][15] , \spm_in[SDATA][14] , \spm_in[SDATA][13] ,
         \spm_in[SDATA][12] , \spm_in[SDATA][11] , \spm_in[SDATA][10] ,
         \spm_in[SDATA][9] , \spm_in[SDATA][8] , \spm_in[SDATA][7] ,
         \spm_in[SDATA][6] , \spm_in[SDATA][5] , \spm_in[SDATA][4] ,
         \spm_in[SDATA][3] , \spm_in[SDATA][2] , \spm_in[SDATA][1] ,
         \spm_in[SDATA][0] ;
  output \proc_out[SCMDACCEPT] , \proc_out[SRESP] , \proc_out[SDATA][31] ,
         \proc_out[SDATA][30] , \proc_out[SDATA][29] , \proc_out[SDATA][28] ,
         \proc_out[SDATA][27] , \proc_out[SDATA][26] , \proc_out[SDATA][25] ,
         \proc_out[SDATA][24] , \proc_out[SDATA][23] , \proc_out[SDATA][22] ,
         \proc_out[SDATA][21] , \proc_out[SDATA][20] , \proc_out[SDATA][19] ,
         \proc_out[SDATA][18] , \proc_out[SDATA][17] , \proc_out[SDATA][16] ,
         \proc_out[SDATA][15] , \proc_out[SDATA][14] , \proc_out[SDATA][13] ,
         \proc_out[SDATA][12] , \proc_out[SDATA][11] , \proc_out[SDATA][10] ,
         \proc_out[SDATA][9] , \proc_out[SDATA][8] , \proc_out[SDATA][7] ,
         \proc_out[SDATA][6] , \proc_out[SDATA][5] , \proc_out[SDATA][4] ,
         \proc_out[SDATA][3] , \proc_out[SDATA][2] , \proc_out[SDATA][1] ,
         \proc_out[SDATA][0] , \spm_out[MCMD][1] , \spm_out[MCMD][0] ,
         \spm_out[MADDR][31] , \spm_out[MADDR][30] , \spm_out[MADDR][29] ,
         \spm_out[MADDR][28] , \spm_out[MADDR][27] , \spm_out[MADDR][26] ,
         \spm_out[MADDR][25] , \spm_out[MADDR][24] , \spm_out[MADDR][23] ,
         \spm_out[MADDR][22] , \spm_out[MADDR][21] , \spm_out[MADDR][20] ,
         \spm_out[MADDR][19] , \spm_out[MADDR][18] , \spm_out[MADDR][17] ,
         \spm_out[MADDR][16] , \spm_out[MADDR][15] , \spm_out[MADDR][14] ,
         \spm_out[MADDR][13] , \spm_out[MADDR][12] , \spm_out[MADDR][11] ,
         \spm_out[MADDR][10] , \spm_out[MADDR][9] , \spm_out[MADDR][8] ,
         \spm_out[MADDR][7] , \spm_out[MADDR][6] , \spm_out[MADDR][5] ,
         \spm_out[MADDR][4] , \spm_out[MADDR][3] , \spm_out[MADDR][2] ,
         \spm_out[MADDR][1] , \spm_out[MADDR][0] , \spm_out[MDATA][63] ,
         \spm_out[MDATA][62] , \spm_out[MDATA][61] , \spm_out[MDATA][60] ,
         \spm_out[MDATA][59] , \spm_out[MDATA][58] , \spm_out[MDATA][57] ,
         \spm_out[MDATA][56] , \spm_out[MDATA][55] , \spm_out[MDATA][54] ,
         \spm_out[MDATA][53] , \spm_out[MDATA][52] , \spm_out[MDATA][51] ,
         \spm_out[MDATA][50] , \spm_out[MDATA][49] , \spm_out[MDATA][48] ,
         \spm_out[MDATA][47] , \spm_out[MDATA][46] , \spm_out[MDATA][45] ,
         \spm_out[MDATA][44] , \spm_out[MDATA][43] , \spm_out[MDATA][42] ,
         \spm_out[MDATA][41] , \spm_out[MDATA][40] , \spm_out[MDATA][39] ,
         \spm_out[MDATA][38] , \spm_out[MDATA][37] , \spm_out[MDATA][36] ,
         \spm_out[MDATA][35] , \spm_out[MDATA][34] , \spm_out[MDATA][33] ,
         \spm_out[MDATA][32] , \spm_out[MDATA][31] , \spm_out[MDATA][30] ,
         \spm_out[MDATA][29] , \spm_out[MDATA][28] , \spm_out[MDATA][27] ,
         \spm_out[MDATA][26] , \spm_out[MDATA][25] , \spm_out[MDATA][24] ,
         \spm_out[MDATA][23] , \spm_out[MDATA][22] , \spm_out[MDATA][21] ,
         \spm_out[MDATA][20] , \spm_out[MDATA][19] , \spm_out[MDATA][18] ,
         \spm_out[MDATA][17] , \spm_out[MDATA][16] , \spm_out[MDATA][15] ,
         \spm_out[MDATA][14] , \spm_out[MDATA][13] , \spm_out[MDATA][12] ,
         \spm_out[MDATA][11] , \spm_out[MDATA][10] , \spm_out[MDATA][9] ,
         \spm_out[MDATA][8] , \spm_out[MDATA][7] , \spm_out[MDATA][6] ,
         \spm_out[MDATA][5] , \spm_out[MDATA][4] , \spm_out[MDATA][3] ,
         \spm_out[MDATA][2] , \spm_out[MDATA][1] , \spm_out[MDATA][0] ;
  wire   \spm_out[MCMD][0] , \phase_prev[0] , \phase_next[1] , vld_pkt, n7, n8,
         n9, n10, n11, n12, n13, n14, n16, n33, n36, n38, n40, n60, n61, n63,
         n65, n66, n67, n68, n69, n70, n71, n76, n81, n82, n83, n85, n86, n92,
         n96, n97, n98, n99, n100, n107, n110, n115, n119, n121, n123, n126,
         n131, n135, n141, n143, n145, n146, n147, n148, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n307, n308, n309,
         n315, n316, n317, n318, n319, n320, n321, n322, \add_545/A[8] ,
         \add_545/A[9] , \add_545/A[10] , \add_545/A[11] , \add_545/A[12] ,
         \add_545/A[13] , \add_545/A[14] , \add_545/A[15] , \sub_544/A[1] ,
         \sub_544/A[2] , \sub_544/A[3] , \sub_544/A[4] , \sub_544/A[5] ,
         \sub_544/A[6] , \sub_544/A[7] , \sub_544/A[8] , \sub_544/A[9] ,
         \sub_544/A[10] , \sub_544/A[11] , \sub_544/A[12] , n1, n2, n3, n4, n5,
         n6, n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n34, n35, n37, n39, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n62,
         n64, n72, n73, n74, n75, n77, n78, n79, n80, n84, n87, n88, n89, n90,
         n91, n93, n94, n95, n101, n102, n103, n104, n105, n106, n108, n109,
         n111, n112, n113, n114, n116, n117, n118, n120, n122, n124, n125,
         n127, n128, n129, n130, n132, n133, n134, n136, n137, n138, n139,
         n140, n142, n144, n149, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n310, n311, n312, n313,
         n314, n323, n324, n325, n326, n327, n328, n329, n330, n331, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672;
  wire   [2:0] slt_index;
  wire   [2:0] dma_ren;
  wire   [2:0] dma_wen;
  wire   [1:0] dma_waddr;
  wire   [63:0] dma_wdata;
  wire   [1:0] dma_raddr;
  wire   [63:0] dma_rdata;
  wire   [4:0] slt_entry;
  wire   [1:0] state_cnt;
  wire   [4:0] config_reg;
  wire   [70:64] flit_buf;
  wire   [34:0] phitIn;
  wire   [31:0] mux_out;
  wire   [31:0] dOut_l;
  wire   [34:32] phit_togo;
  wire   [34:0] phitOut0;
  wire   [34:0] phitOut1;
  wire   [34:0] phitOut2;
  wire   [13:0] dma_cnt_new;
  wire   [15:0] dma_rp_new;
  wire   [15:0] dma_wp_new;
  wire   [6:0] address;
  wire   [31:0] dIn_h;
  assign \spm_out[MADDR][15]  = 1'b0;
  assign \spm_out[MADDR][16]  = 1'b0;
  assign \spm_out[MADDR][17]  = 1'b0;
  assign \spm_out[MADDR][18]  = 1'b0;
  assign \spm_out[MADDR][19]  = 1'b0;
  assign \spm_out[MADDR][20]  = 1'b0;
  assign \spm_out[MADDR][21]  = 1'b0;
  assign \spm_out[MADDR][22]  = 1'b0;
  assign \spm_out[MADDR][23]  = 1'b0;
  assign \spm_out[MADDR][24]  = 1'b0;
  assign \spm_out[MADDR][25]  = 1'b0;
  assign \spm_out[MADDR][26]  = 1'b0;
  assign \spm_out[MADDR][27]  = 1'b0;
  assign \spm_out[MADDR][28]  = 1'b0;
  assign \spm_out[MADDR][29]  = 1'b0;
  assign \spm_out[MADDR][30]  = 1'b0;
  assign \spm_out[MADDR][31]  = 1'b0;
  assign \spm_out[MCMD][1]  = \spm_out[MCMD][0] ;

  HS65_LS_DFPRQX9 \state_cnt_reg[0]  ( .D(n136), .CP(na_clk), .RN(n336), .Q(
        state_cnt[0]) );
  HS65_LS_DFPRQX9 \state_cnt_reg[1]  ( .D(n595), .CP(na_clk), .RN(n337), .Q(
        state_cnt[1]) );
  HS65_LS_DFPRQX9 \phase_next_reg[1]  ( .D(n321), .CP(na_clk), .RN(n339), .Q(
        \phase_next[1] ) );
  HS65_LS_DFPRQX9 \dOut_l_reg[31]  ( .D(n292), .CP(na_clk), .RN(n349), .Q(
        dOut_l[31]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[30]  ( .D(n291), .CP(na_clk), .RN(n337), .Q(
        dOut_l[30]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[29]  ( .D(n290), .CP(na_clk), .RN(n341), .Q(
        dOut_l[29]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[28]  ( .D(n289), .CP(na_clk), .RN(n348), .Q(
        dOut_l[28]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[27]  ( .D(n288), .CP(na_clk), .RN(n340), .Q(
        dOut_l[27]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[26]  ( .D(n287), .CP(na_clk), .RN(n338), .Q(
        dOut_l[26]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[25]  ( .D(n286), .CP(na_clk), .RN(n339), .Q(
        dOut_l[25]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[24]  ( .D(n285), .CP(na_clk), .RN(n344), .Q(
        dOut_l[24]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[23]  ( .D(n284), .CP(na_clk), .RN(n350), .Q(
        dOut_l[23]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[22]  ( .D(n283), .CP(na_clk), .RN(n338), .Q(
        dOut_l[22]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[21]  ( .D(n282), .CP(na_clk), .RN(n336), .Q(
        dOut_l[21]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[20]  ( .D(n281), .CP(na_clk), .RN(n340), .Q(
        dOut_l[20]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[19]  ( .D(n280), .CP(na_clk), .RN(n337), .Q(
        dOut_l[19]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[18]  ( .D(n279), .CP(na_clk), .RN(n342), .Q(
        dOut_l[18]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[17]  ( .D(n278), .CP(na_clk), .RN(n347), .Q(
        dOut_l[17]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[16]  ( .D(n277), .CP(na_clk), .RN(n337), .Q(
        dOut_l[16]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[15]  ( .D(n276), .CP(na_clk), .RN(n336), .Q(
        dOut_l[15]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[14]  ( .D(n275), .CP(na_clk), .RN(n340), .Q(
        dOut_l[14]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[13]  ( .D(n274), .CP(na_clk), .RN(n342), .Q(
        dOut_l[13]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[12]  ( .D(n273), .CP(na_clk), .RN(n346), .Q(
        dOut_l[12]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[11]  ( .D(n272), .CP(na_clk), .RN(n350), .Q(
        dOut_l[11]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[10]  ( .D(n271), .CP(na_clk), .RN(n341), .Q(
        dOut_l[10]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[9]  ( .D(n270), .CP(na_clk), .RN(n345), .Q(
        dOut_l[9]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[8]  ( .D(n269), .CP(na_clk), .RN(n343), .Q(
        dOut_l[8]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[7]  ( .D(n268), .CP(na_clk), .RN(n348), .Q(
        dOut_l[7]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[6]  ( .D(n267), .CP(na_clk), .RN(n349), .Q(
        dOut_l[6]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[5]  ( .D(n266), .CP(na_clk), .RN(n339), .Q(
        dOut_l[5]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[4]  ( .D(n265), .CP(na_clk), .RN(n344), .Q(
        dOut_l[4]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[3]  ( .D(n264), .CP(na_clk), .RN(n338), .Q(
        dOut_l[3]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[2]  ( .D(n263), .CP(na_clk), .RN(n345), .Q(
        dOut_l[2]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[1]  ( .D(n262), .CP(na_clk), .RN(n345), .Q(
        dOut_l[1]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[0]  ( .D(n261), .CP(na_clk), .RN(n345), .Q(
        dOut_l[0]) );
  HS65_LS_DFPRQX9 \phitIn_reg[34]  ( .D(pkt_in[34]), .CP(na_clk), .RN(n345), 
        .Q(phitIn[34]) );
  HS65_LS_DFPRQX9 \phitIn_reg[33]  ( .D(pkt_in[33]), .CP(na_clk), .RN(n345), 
        .Q(phitIn[33]) );
  HS65_LS_DFPRQX9 vld_pkt_reg ( .D(n318), .CP(na_clk), .RN(n345), .Q(vld_pkt)
         );
  HS65_LS_DFPRQX9 \phitIn_reg[32]  ( .D(pkt_in[32]), .CP(na_clk), .RN(n345), 
        .Q(phitIn[32]) );
  HS65_LS_DFPRQX9 \phitIn_reg[31]  ( .D(pkt_in[31]), .CP(na_clk), .RN(n345), 
        .Q(phitIn[31]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[31]  ( .D(n260), .CP(na_clk), .RN(n345), .Q(
        dIn_h[31]) );
  HS65_LS_DFPRQX9 \phitIn_reg[30]  ( .D(pkt_in[30]), .CP(na_clk), .RN(n345), 
        .Q(phitIn[30]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[30]  ( .D(n259), .CP(na_clk), .RN(n345), .Q(
        dIn_h[30]) );
  HS65_LS_DFPRQX9 \phitIn_reg[29]  ( .D(pkt_in[29]), .CP(na_clk), .RN(n345), 
        .Q(phitIn[29]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[29]  ( .D(n258), .CP(na_clk), .RN(n345), .Q(
        dIn_h[29]) );
  HS65_LS_DFPRQX9 \phitIn_reg[28]  ( .D(pkt_in[28]), .CP(na_clk), .RN(n345), 
        .Q(phitIn[28]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[28]  ( .D(n257), .CP(na_clk), .RN(n345), .Q(
        dIn_h[28]) );
  HS65_LS_DFPRQX9 \phitIn_reg[27]  ( .D(pkt_in[27]), .CP(na_clk), .RN(n346), 
        .Q(phitIn[27]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[27]  ( .D(n256), .CP(na_clk), .RN(n346), .Q(
        dIn_h[27]) );
  HS65_LS_DFPRQX9 \phitIn_reg[26]  ( .D(pkt_in[26]), .CP(na_clk), .RN(n346), 
        .Q(phitIn[26]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[26]  ( .D(n255), .CP(na_clk), .RN(n346), .Q(
        dIn_h[26]) );
  HS65_LS_DFPRQX9 \phitIn_reg[25]  ( .D(pkt_in[25]), .CP(na_clk), .RN(n346), 
        .Q(phitIn[25]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[25]  ( .D(n254), .CP(na_clk), .RN(n346), .Q(
        dIn_h[25]) );
  HS65_LS_DFPRQX9 \phitIn_reg[24]  ( .D(pkt_in[24]), .CP(na_clk), .RN(n346), 
        .Q(phitIn[24]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[24]  ( .D(n253), .CP(na_clk), .RN(n346), .Q(
        dIn_h[24]) );
  HS65_LS_DFPRQX9 \phitIn_reg[23]  ( .D(pkt_in[23]), .CP(na_clk), .RN(n346), 
        .Q(phitIn[23]) );
  HS65_LS_DFPRQX9 \address_reg[6]  ( .D(n252), .CP(na_clk), .RN(n346), .Q(
        address[6]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[23]  ( .D(n251), .CP(na_clk), .RN(n346), .Q(
        dIn_h[23]) );
  HS65_LS_DFPRQX9 \phitIn_reg[22]  ( .D(pkt_in[22]), .CP(na_clk), .RN(n346), 
        .Q(phitIn[22]) );
  HS65_LS_DFPRQX9 \address_reg[5]  ( .D(n250), .CP(na_clk), .RN(n346), .Q(
        address[5]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[22]  ( .D(n249), .CP(na_clk), .RN(n346), .Q(
        dIn_h[22]) );
  HS65_LS_DFPRQX9 \phitIn_reg[21]  ( .D(pkt_in[21]), .CP(na_clk), .RN(n346), 
        .Q(phitIn[21]) );
  HS65_LS_DFPRQX9 \address_reg[4]  ( .D(n248), .CP(na_clk), .RN(n339), .Q(
        address[4]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[21]  ( .D(n247), .CP(na_clk), .RN(n338), .Q(
        dIn_h[21]) );
  HS65_LS_DFPRQX9 \phitIn_reg[20]  ( .D(pkt_in[20]), .CP(na_clk), .RN(n341), 
        .Q(phitIn[20]) );
  HS65_LS_DFPRQX9 \address_reg[3]  ( .D(n246), .CP(na_clk), .RN(n336), .Q(
        address[3]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[20]  ( .D(n245), .CP(na_clk), .RN(n342), .Q(
        dIn_h[20]) );
  HS65_LS_DFPRQX9 \phitIn_reg[19]  ( .D(pkt_in[19]), .CP(na_clk), .RN(n344), 
        .Q(phitIn[19]) );
  HS65_LS_DFPRQX9 \address_reg[2]  ( .D(n244), .CP(na_clk), .RN(n349), .Q(
        address[2]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[19]  ( .D(n243), .CP(na_clk), .RN(n348), .Q(
        dIn_h[19]) );
  HS65_LS_DFPRQX9 \phitIn_reg[18]  ( .D(pkt_in[18]), .CP(na_clk), .RN(n341), 
        .Q(phitIn[18]) );
  HS65_LS_DFPRQX9 \address_reg[1]  ( .D(n242), .CP(na_clk), .RN(n345), .Q(
        address[1]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[18]  ( .D(n241), .CP(na_clk), .RN(n343), .Q(
        dIn_h[18]) );
  HS65_LS_DFPRQX9 \phitIn_reg[17]  ( .D(pkt_in[17]), .CP(na_clk), .RN(n346), 
        .Q(phitIn[17]) );
  HS65_LS_DFPRQX9 \address_reg[0]  ( .D(n240), .CP(na_clk), .RN(n343), .Q(
        address[0]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[17]  ( .D(n239), .CP(na_clk), .RN(n347), .Q(
        dIn_h[17]) );
  HS65_LS_DFPRQX9 \phitIn_reg[16]  ( .D(pkt_in[16]), .CP(na_clk), .RN(n347), 
        .Q(phitIn[16]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[16]  ( .D(n238), .CP(na_clk), .RN(n347), .Q(
        dIn_h[16]) );
  HS65_LS_DFPRQX9 \phitIn_reg[15]  ( .D(pkt_in[15]), .CP(na_clk), .RN(n347), 
        .Q(phitIn[15]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[15]  ( .D(n237), .CP(na_clk), .RN(n347), .Q(
        dIn_h[15]) );
  HS65_LS_DFPRQX9 \phitIn_reg[14]  ( .D(pkt_in[14]), .CP(na_clk), .RN(n347), 
        .Q(phitIn[14]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[14]  ( .D(n236), .CP(na_clk), .RN(n347), .Q(
        dIn_h[14]) );
  HS65_LS_DFPRQX9 \phitIn_reg[13]  ( .D(pkt_in[13]), .CP(na_clk), .RN(n347), 
        .Q(phitIn[13]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[13]  ( .D(n235), .CP(na_clk), .RN(n347), .Q(
        dIn_h[13]) );
  HS65_LS_DFPRQX9 \phitIn_reg[12]  ( .D(pkt_in[12]), .CP(na_clk), .RN(n347), 
        .Q(phitIn[12]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[12]  ( .D(n234), .CP(na_clk), .RN(n347), .Q(
        dIn_h[12]) );
  HS65_LS_DFPRQX9 \phitIn_reg[11]  ( .D(pkt_in[11]), .CP(na_clk), .RN(n347), 
        .Q(phitIn[11]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[11]  ( .D(n233), .CP(na_clk), .RN(n347), .Q(
        dIn_h[11]) );
  HS65_LS_DFPRQX9 \phitIn_reg[10]  ( .D(pkt_in[10]), .CP(na_clk), .RN(n347), 
        .Q(phitIn[10]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[10]  ( .D(n232), .CP(na_clk), .RN(n347), .Q(
        dIn_h[10]) );
  HS65_LS_DFPRQX9 \phitIn_reg[9]  ( .D(pkt_in[9]), .CP(na_clk), .RN(n347), .Q(
        phitIn[9]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[9]  ( .D(n231), .CP(na_clk), .RN(n348), .Q(
        dIn_h[9]) );
  HS65_LS_DFPRQX9 \phitIn_reg[8]  ( .D(pkt_in[8]), .CP(na_clk), .RN(n348), .Q(
        phitIn[8]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[8]  ( .D(n230), .CP(na_clk), .RN(n348), .Q(
        dIn_h[8]) );
  HS65_LS_DFPRQX9 \phitIn_reg[7]  ( .D(pkt_in[7]), .CP(na_clk), .RN(n348), .Q(
        phitIn[7]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[7]  ( .D(n229), .CP(na_clk), .RN(n348), .Q(
        dIn_h[7]) );
  HS65_LS_DFPRQX9 \phitIn_reg[6]  ( .D(pkt_in[6]), .CP(na_clk), .RN(n348), .Q(
        phitIn[6]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[6]  ( .D(n228), .CP(na_clk), .RN(n348), .Q(
        dIn_h[6]) );
  HS65_LS_DFPRQX9 \phitIn_reg[5]  ( .D(pkt_in[5]), .CP(na_clk), .RN(n348), .Q(
        phitIn[5]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[5]  ( .D(n227), .CP(na_clk), .RN(n348), .Q(
        dIn_h[5]) );
  HS65_LS_DFPRQX9 \phitIn_reg[4]  ( .D(pkt_in[4]), .CP(na_clk), .RN(n348), .Q(
        phitIn[4]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[4]  ( .D(n226), .CP(na_clk), .RN(n348), .Q(
        dIn_h[4]) );
  HS65_LS_DFPRQX9 \phitIn_reg[3]  ( .D(pkt_in[3]), .CP(na_clk), .RN(n348), .Q(
        phitIn[3]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[3]  ( .D(n225), .CP(na_clk), .RN(n348), .Q(
        dIn_h[3]) );
  HS65_LS_DFPRQX9 \phitIn_reg[2]  ( .D(pkt_in[2]), .CP(na_clk), .RN(n348), .Q(
        phitIn[2]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[2]  ( .D(n224), .CP(na_clk), .RN(n348), .Q(
        dIn_h[2]) );
  HS65_LS_DFPRQX9 \phitIn_reg[1]  ( .D(pkt_in[1]), .CP(na_clk), .RN(n349), .Q(
        phitIn[1]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[1]  ( .D(n223), .CP(na_clk), .RN(n349), .Q(
        dIn_h[1]) );
  HS65_LS_DFPRQX9 \phitIn_reg[0]  ( .D(pkt_in[0]), .CP(na_clk), .RN(n349), .Q(
        phitIn[0]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[0]  ( .D(n222), .CP(na_clk), .RN(n349), .Q(
        dIn_h[0]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[34]  ( .D(phit_togo[34]), .CP(na_clk), .RN(
        n349), .Q(phitOut0[34]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[33]  ( .D(n328), .CP(na_clk), .RN(n349), .Q(
        phitOut0[33]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[32]  ( .D(phit_togo[32]), .CP(na_clk), .RN(
        n349), .Q(phitOut0[32]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[31]  ( .D(mux_out[31]), .CP(na_clk), .RN(n349), 
        .Q(phitOut0[31]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[30]  ( .D(mux_out[30]), .CP(na_clk), .RN(n349), 
        .Q(phitOut0[30]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[29]  ( .D(mux_out[29]), .CP(na_clk), .RN(n349), 
        .Q(phitOut0[29]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[28]  ( .D(mux_out[28]), .CP(na_clk), .RN(n349), 
        .Q(phitOut0[28]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[27]  ( .D(mux_out[27]), .CP(na_clk), .RN(n349), 
        .Q(phitOut0[27]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[26]  ( .D(mux_out[26]), .CP(na_clk), .RN(n349), 
        .Q(phitOut0[26]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[25]  ( .D(mux_out[25]), .CP(na_clk), .RN(n349), 
        .Q(phitOut0[25]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[24]  ( .D(mux_out[24]), .CP(na_clk), .RN(n349), 
        .Q(phitOut0[24]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[23]  ( .D(mux_out[23]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[23]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[22]  ( .D(mux_out[22]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[22]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[21]  ( .D(mux_out[21]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[21]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[20]  ( .D(mux_out[20]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[20]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[19]  ( .D(mux_out[19]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[19]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[18]  ( .D(mux_out[18]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[18]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[17]  ( .D(mux_out[17]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[17]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[16]  ( .D(mux_out[16]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[16]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[15]  ( .D(mux_out[15]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[15]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[14]  ( .D(mux_out[14]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[14]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[13]  ( .D(mux_out[13]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[13]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[12]  ( .D(mux_out[12]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[12]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[11]  ( .D(mux_out[11]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[11]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[10]  ( .D(mux_out[10]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[10]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[9]  ( .D(mux_out[9]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[9]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[8]  ( .D(mux_out[8]), .CP(na_clk), .RN(n342), 
        .Q(phitOut0[8]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[7]  ( .D(mux_out[7]), .CP(na_clk), .RN(n341), 
        .Q(phitOut0[7]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[6]  ( .D(mux_out[6]), .CP(na_clk), .RN(n339), 
        .Q(phitOut0[6]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[5]  ( .D(mux_out[5]), .CP(na_clk), .RN(n338), 
        .Q(phitOut0[5]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[4]  ( .D(mux_out[4]), .CP(na_clk), .RN(n337), 
        .Q(phitOut0[4]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[3]  ( .D(mux_out[3]), .CP(na_clk), .RN(n340), 
        .Q(phitOut0[3]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[2]  ( .D(mux_out[2]), .CP(na_clk), .RN(n336), 
        .Q(phitOut0[2]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[1]  ( .D(mux_out[1]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[1]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[0]  ( .D(mux_out[0]), .CP(na_clk), .RN(n343), 
        .Q(phitOut0[0]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[34]  ( .D(phitOut0[34]), .CP(na_clk), .RN(n340), .Q(phitOut1[34]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[33]  ( .D(phitOut0[33]), .CP(na_clk), .RN(n336), .Q(phitOut1[33]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[32]  ( .D(phitOut0[32]), .CP(na_clk), .RN(n336), .Q(phitOut1[32]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[31]  ( .D(phitOut0[31]), .CP(na_clk), .RN(n336), .Q(phitOut1[31]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[30]  ( .D(phitOut0[30]), .CP(na_clk), .RN(n336), .Q(phitOut1[30]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[29]  ( .D(phitOut0[29]), .CP(na_clk), .RN(n336), .Q(phitOut1[29]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[28]  ( .D(phitOut0[28]), .CP(na_clk), .RN(n336), .Q(phitOut1[28]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[27]  ( .D(phitOut0[27]), .CP(na_clk), .RN(n336), .Q(phitOut1[27]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[26]  ( .D(phitOut0[26]), .CP(na_clk), .RN(n336), .Q(phitOut1[26]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[25]  ( .D(phitOut0[25]), .CP(na_clk), .RN(n336), .Q(phitOut1[25]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[24]  ( .D(phitOut0[24]), .CP(na_clk), .RN(n336), .Q(phitOut1[24]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[23]  ( .D(phitOut0[23]), .CP(na_clk), .RN(n336), .Q(phitOut1[23]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[22]  ( .D(phitOut0[22]), .CP(na_clk), .RN(n336), .Q(phitOut1[22]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[21]  ( .D(phitOut0[21]), .CP(na_clk), .RN(n336), .Q(phitOut1[21]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[20]  ( .D(phitOut0[20]), .CP(na_clk), .RN(n343), .Q(phitOut1[20]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[19]  ( .D(phitOut0[19]), .CP(na_clk), .RN(n347), .Q(phitOut1[19]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[18]  ( .D(phitOut0[18]), .CP(na_clk), .RN(n342), .Q(phitOut1[18]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[17]  ( .D(phitOut0[17]), .CP(na_clk), .RN(n345), .Q(phitOut1[17]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[16]  ( .D(phitOut0[16]), .CP(na_clk), .RN(n346), .Q(phitOut1[16]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[15]  ( .D(phitOut0[15]), .CP(na_clk), .RN(n350), .Q(phitOut1[15]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[14]  ( .D(phitOut0[14]), .CP(na_clk), .RN(n340), .Q(phitOut1[14]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[13]  ( .D(phitOut0[13]), .CP(na_clk), .RN(n347), .Q(phitOut1[13]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[12]  ( .D(phitOut0[12]), .CP(na_clk), .RN(n346), .Q(phitOut1[12]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[11]  ( .D(phitOut0[11]), .CP(na_clk), .RN(n345), .Q(phitOut1[11]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[10]  ( .D(phitOut0[10]), .CP(na_clk), .RN(n350), .Q(phitOut1[10]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[9]  ( .D(phitOut0[9]), .CP(na_clk), .RN(n344), 
        .Q(phitOut1[9]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[8]  ( .D(phitOut0[8]), .CP(na_clk), .RN(n349), 
        .Q(phitOut1[8]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[7]  ( .D(phitOut0[7]), .CP(na_clk), .RN(n348), 
        .Q(phitOut1[7]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[6]  ( .D(phitOut0[6]), .CP(na_clk), .RN(n337), 
        .Q(phitOut1[6]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[5]  ( .D(phitOut0[5]), .CP(na_clk), .RN(n337), 
        .Q(phitOut1[5]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[4]  ( .D(phitOut0[4]), .CP(na_clk), .RN(n337), 
        .Q(phitOut1[4]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[3]  ( .D(phitOut0[3]), .CP(na_clk), .RN(n337), 
        .Q(phitOut1[3]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[2]  ( .D(phitOut0[2]), .CP(na_clk), .RN(n337), 
        .Q(phitOut1[2]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[1]  ( .D(phitOut0[1]), .CP(na_clk), .RN(n337), 
        .Q(phitOut1[1]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[0]  ( .D(phitOut0[0]), .CP(na_clk), .RN(n337), 
        .Q(phitOut1[0]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[34]  ( .D(phitOut1[34]), .CP(na_clk), .RN(n337), .Q(phitOut2[34]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[33]  ( .D(phitOut1[33]), .CP(na_clk), .RN(n337), .Q(phitOut2[33]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[32]  ( .D(phitOut1[32]), .CP(na_clk), .RN(n337), .Q(phitOut2[32]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[31]  ( .D(phitOut1[31]), .CP(na_clk), .RN(n337), .Q(phitOut2[31]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[30]  ( .D(phitOut1[30]), .CP(na_clk), .RN(n337), .Q(phitOut2[30]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[29]  ( .D(phitOut1[29]), .CP(na_clk), .RN(n337), .Q(phitOut2[29]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[28]  ( .D(phitOut1[28]), .CP(na_clk), .RN(n337), .Q(phitOut2[28]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[27]  ( .D(phitOut1[27]), .CP(na_clk), .RN(n337), .Q(phitOut2[27]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[26]  ( .D(phitOut1[26]), .CP(na_clk), .RN(n338), .Q(phitOut2[26]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[25]  ( .D(phitOut1[25]), .CP(na_clk), .RN(n338), .Q(phitOut2[25]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[24]  ( .D(phitOut1[24]), .CP(na_clk), .RN(n338), .Q(phitOut2[24]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[23]  ( .D(phitOut1[23]), .CP(na_clk), .RN(n338), .Q(phitOut2[23]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[22]  ( .D(phitOut1[22]), .CP(na_clk), .RN(n338), .Q(phitOut2[22]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[21]  ( .D(phitOut1[21]), .CP(na_clk), .RN(n338), .Q(phitOut2[21]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[20]  ( .D(phitOut1[20]), .CP(na_clk), .RN(n338), .Q(phitOut2[20]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[19]  ( .D(phitOut1[19]), .CP(na_clk), .RN(n338), .Q(phitOut2[19]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[18]  ( .D(phitOut1[18]), .CP(na_clk), .RN(n338), .Q(phitOut2[18]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[17]  ( .D(phitOut1[17]), .CP(na_clk), .RN(n338), .Q(phitOut2[17]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[16]  ( .D(phitOut1[16]), .CP(na_clk), .RN(n338), .Q(phitOut2[16]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[15]  ( .D(phitOut1[15]), .CP(na_clk), .RN(n338), .Q(phitOut2[15]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[14]  ( .D(phitOut1[14]), .CP(na_clk), .RN(n338), .Q(phitOut2[14]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[13]  ( .D(phitOut1[13]), .CP(na_clk), .RN(n338), .Q(phitOut2[13]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[12]  ( .D(phitOut1[12]), .CP(na_clk), .RN(n338), .Q(phitOut2[12]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[11]  ( .D(phitOut1[11]), .CP(na_clk), .RN(n339), .Q(phitOut2[11]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[10]  ( .D(phitOut1[10]), .CP(na_clk), .RN(n339), .Q(phitOut2[10]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[9]  ( .D(phitOut1[9]), .CP(na_clk), .RN(n339), 
        .Q(phitOut2[9]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[8]  ( .D(phitOut1[8]), .CP(na_clk), .RN(n339), 
        .Q(phitOut2[8]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[7]  ( .D(phitOut1[7]), .CP(na_clk), .RN(n339), 
        .Q(phitOut2[7]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[6]  ( .D(phitOut1[6]), .CP(na_clk), .RN(n339), 
        .Q(phitOut2[6]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[5]  ( .D(phitOut1[5]), .CP(na_clk), .RN(n339), 
        .Q(phitOut2[5]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[4]  ( .D(phitOut1[4]), .CP(na_clk), .RN(n339), 
        .Q(phitOut2[4]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[3]  ( .D(phitOut1[3]), .CP(na_clk), .RN(n339), 
        .Q(phitOut2[3]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[2]  ( .D(phitOut1[2]), .CP(na_clk), .RN(n339), 
        .Q(phitOut2[2]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[1]  ( .D(phitOut1[1]), .CP(na_clk), .RN(n339), 
        .Q(phitOut2[1]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[0]  ( .D(phitOut1[0]), .CP(na_clk), .RN(n339), 
        .Q(phitOut2[0]) );
  HS65_LS_DFPRQX9 \config_reg_reg[4]  ( .D(\proc_in[MCMD][1] ), .CP(na_clk), 
        .RN(n339), .Q(config_reg[4]) );
  HS65_LS_DFPRQX9 \config_reg_reg[3]  ( .D(n322), .CP(na_clk), .RN(n339), .Q(
        config_reg[3]) );
  HS65_LS_DFPRQX9 \config_reg_reg[2]  ( .D(n650), .CP(na_clk), .RN(n339), .Q(
        config_reg[2]) );
  HS65_LS_DFPRQX9 \config_reg_reg[1]  ( .D(n651), .CP(na_clk), .RN(n340), .Q(
        config_reg[1]) );
  HS65_LS_DFPRQX9 \config_reg_reg[0]  ( .D(n649), .CP(na_clk), .RN(n340), .Q(
        config_reg[0]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[70]  ( .D(n221), .CP(na_clk), .RN(n340), .Q(
        flit_buf[70]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[69]  ( .D(n220), .CP(na_clk), .RN(n340), .Q(
        flit_buf[69]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[68]  ( .D(n219), .CP(na_clk), .RN(n340), .Q(
        flit_buf[68]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[67]  ( .D(n218), .CP(na_clk), .RN(n340), .Q(
        flit_buf[67]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[66]  ( .D(n217), .CP(na_clk), .RN(n340), .Q(
        flit_buf[66]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[65]  ( .D(n216), .CP(na_clk), .RN(n340), .Q(
        flit_buf[65]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[64]  ( .D(n215), .CP(na_clk), .RN(n340), .Q(
        flit_buf[64]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[63]  ( .D(n214), .CP(na_clk), .RN(n340), .Q(
        \spm_out[MDATA][63] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[62]  ( .D(n213), .CP(na_clk), .RN(n340), .Q(
        \spm_out[MDATA][62] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[61]  ( .D(n212), .CP(na_clk), .RN(n340), .Q(
        \spm_out[MDATA][61] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[60]  ( .D(n211), .CP(na_clk), .RN(n340), .Q(
        \spm_out[MDATA][60] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[59]  ( .D(n210), .CP(na_clk), .RN(n340), .Q(
        \spm_out[MDATA][59] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[58]  ( .D(n209), .CP(na_clk), .RN(n341), .Q(
        \spm_out[MDATA][58] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[57]  ( .D(n208), .CP(na_clk), .RN(n341), .Q(
        \spm_out[MDATA][57] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[56]  ( .D(n207), .CP(na_clk), .RN(n341), .Q(
        \spm_out[MDATA][56] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[55]  ( .D(n206), .CP(na_clk), .RN(n341), .Q(
        \spm_out[MDATA][55] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[54]  ( .D(n205), .CP(na_clk), .RN(n341), .Q(
        \spm_out[MDATA][54] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[53]  ( .D(n204), .CP(na_clk), .RN(n341), .Q(
        \spm_out[MDATA][53] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[52]  ( .D(n203), .CP(na_clk), .RN(n341), .Q(
        \spm_out[MDATA][52] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[51]  ( .D(n202), .CP(na_clk), .RN(n341), .Q(
        \spm_out[MDATA][51] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[50]  ( .D(n201), .CP(na_clk), .RN(n341), .Q(
        \spm_out[MDATA][50] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[49]  ( .D(n200), .CP(na_clk), .RN(n341), .Q(
        \spm_out[MDATA][49] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[48]  ( .D(n199), .CP(na_clk), .RN(n341), .Q(
        \spm_out[MDATA][48] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[47]  ( .D(n198), .CP(na_clk), .RN(n341), .Q(
        \spm_out[MDATA][47] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[46]  ( .D(n197), .CP(na_clk), .RN(n341), .Q(
        \spm_out[MDATA][46] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[45]  ( .D(n196), .CP(na_clk), .RN(n341), .Q(
        \spm_out[MDATA][45] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[44]  ( .D(n195), .CP(na_clk), .RN(n341), .Q(
        \spm_out[MDATA][44] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[43]  ( .D(n194), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][43] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[42]  ( .D(n193), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][42] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[41]  ( .D(n192), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][41] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[40]  ( .D(n191), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][40] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[39]  ( .D(n190), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][39] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[38]  ( .D(n189), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][38] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[37]  ( .D(n188), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][37] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[36]  ( .D(n187), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][36] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[35]  ( .D(n186), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][35] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[34]  ( .D(n185), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][34] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[33]  ( .D(n184), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][33] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[32]  ( .D(n183), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][32] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[31]  ( .D(n182), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][31] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[30]  ( .D(n181), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][30] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[29]  ( .D(n180), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][29] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[28]  ( .D(n179), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][28] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[27]  ( .D(n178), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][27] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[26]  ( .D(n177), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][26] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[25]  ( .D(n176), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][25] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[24]  ( .D(n175), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][24] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[23]  ( .D(n174), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][23] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[22]  ( .D(n173), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][22] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[21]  ( .D(n172), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][21] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[20]  ( .D(n171), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][20] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[19]  ( .D(n170), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][19] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[18]  ( .D(n169), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][18] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[17]  ( .D(n168), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][17] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[16]  ( .D(n167), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][16] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[15]  ( .D(n166), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][15] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[14]  ( .D(n165), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][14] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[13]  ( .D(n164), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][13] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[12]  ( .D(n163), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][12] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[11]  ( .D(n162), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][11] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[10]  ( .D(n161), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][10] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[9]  ( .D(n160), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][9] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[8]  ( .D(n159), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][8] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[7]  ( .D(n158), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][7] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[6]  ( .D(n157), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][6] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[5]  ( .D(n156), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][5] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[4]  ( .D(n155), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][4] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[3]  ( .D(n154), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][3] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[2]  ( .D(n153), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][2] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[1]  ( .D(n152), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][1] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[0]  ( .D(n151), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][0] ) );
  HS65_LS_DFPRQX9 \phase_prev_reg[0]  ( .D(n315), .CP(na_clk), .RN(n344), .Q(
        \phase_prev[0] ) );
  counter_WIDTH3_0 slt_cnt ( .clk(na_clk), .reset(n351), .enable(n645), .cnt(
        slt_index) );
  dma_sdp_DATA64_ADDR2_0 dma_table ( .clk(na_clk), .reset(n352), .ren(dma_ren), 
        .wen(dma_wen), .waddr(dma_waddr), .wdata(dma_wdata), .raddr(dma_raddr), 
        .rdata(dma_rdata) );
  bram_DATA5_ADDR3_0 slt_table ( .clk(na_clk), .reset(n351), .rd_addr(
        slt_index), .wr_addr({\proc_in[MADDR][2] , \proc_in[MADDR][1] , 
        \proc_in[MADDR][0] }), .wr_data({\proc_in[MDATA][4] , 
        \proc_in[MDATA][3] , \proc_in[MDATA][2] , \proc_in[MDATA][1] , 
        \proc_in[MDATA][0] }), .wr_ena(n648), .rd_data(slt_entry) );
  HS65_LS_DFPRQNX9 vld_buf_reg ( .D(n317), .CP(na_clk), .RN(n344), .QN(n309)
         );
  HS65_LS_DFPRQNX9 dma_ctrl_reg_reg ( .D(n319), .CP(na_clk), .RN(n348), .QN(
        n308) );
  HS65_LS_DFPRQNX9 \phase_next_reg[0]  ( .D(n320), .CP(na_clk), .RN(n349), 
        .QN(n307) );
  HS65_LS_DFPRQX9 \phase_prev_reg[1]  ( .D(n316), .CP(na_clk), .RN(n336), .Q(
        n20) );
  HS65_LS_IVX27 U3 ( .A(n25), .Z(n112) );
  HS65_LS_IVX4 U4 ( .A(n570), .Z(n1) );
  HS65_LS_IVX9 U5 ( .A(n444), .Z(n2) );
  HS65_LS_IVX18 U6 ( .A(n17), .Z(n3) );
  HS65_LS_IVX18 U7 ( .A(n17), .Z(n18) );
  HS65_LS_NAND2X5 U8 ( .A(phitOut2[33]), .B(n471), .Z(n567) );
  HS65_LS_NAND2X5 U9 ( .A(phitOut2[28]), .B(n471), .Z(n552) );
  HS65_LS_NAND2X7 U10 ( .A(phitOut2[1]), .B(n471), .Z(n468) );
  HS65_LS_NAND2X5 U11 ( .A(phitOut2[2]), .B(n471), .Z(n472) );
  HS65_LS_NAND2X5 U12 ( .A(phitOut2[10]), .B(n471), .Z(n497) );
  HS65_LS_NAND2X5 U13 ( .A(phitOut2[16]), .B(n471), .Z(n515) );
  HS65_LS_NAND2X5 U14 ( .A(n19), .B(n460), .Z(n445) );
  HS65_LS_NAND2X5 U15 ( .A(phitOut2[15]), .B(n28), .Z(n512) );
  HS65_LS_NAND2X5 U16 ( .A(phitOut2[6]), .B(n28), .Z(n485) );
  HS65_LS_NAND2X5 U17 ( .A(phitOut2[9]), .B(n28), .Z(n494) );
  HS65_LS_NAND2X5 U18 ( .A(phitOut2[8]), .B(n28), .Z(n491) );
  HS65_LS_NAND2X5 U19 ( .A(phitOut2[11]), .B(n28), .Z(n500) );
  HS65_LS_NAND2X5 U20 ( .A(phitOut2[18]), .B(n28), .Z(n521) );
  HS65_LS_NAND2X5 U21 ( .A(phitOut2[20]), .B(n28), .Z(n528) );
  HS65_LS_NAND2X5 U22 ( .A(phitOut2[25]), .B(n28), .Z(n543) );
  HS65_LS_IVX53 U23 ( .A(n25), .Z(n113) );
  HS65_LS_OR2X9 U24 ( .A(n526), .B(n466), .Z(n41) );
  HS65_LS_IVX9 U25 ( .A(n526), .Z(n17) );
  HS65_LS_NAND2X14 U26 ( .A(n570), .B(n105), .Z(n526) );
  HS65_LH_OAI12X2 U27 ( .A(n308), .B(n645), .C(n314), .Z(n319) );
  HS65_LH_OAI12X2 U28 ( .A(n645), .B(n132), .C(n355), .Z(n357) );
  HS65_LH_IVX2 U29 ( .A(n645), .Z(n29) );
  HS65_LS_NAND2X14 U30 ( .A(slt_entry[4]), .B(n645), .Z(n85) );
  HS65_LS_IVX9 U31 ( .A(n463), .Z(n30) );
  HS65_LS_NAND2X5 U32 ( .A(phitOut2[29]), .B(n471), .Z(n555) );
  HS65_LS_IVX18 U33 ( .A(n462), .Z(n31) );
  HS65_LS_CBI4I1X11 U34 ( .A(n453), .B(n24), .C(n307), .D(n23), .Z(n462) );
  HS65_LS_OAI222X2 U35 ( .A(n656), .B(n86), .C(n644), .D(n29), .E(n655), .F(
        n83), .Z(dma_waddr[0]) );
  HS65_LS_OAI222X2 U36 ( .A(n655), .B(n86), .C(n643), .D(n29), .E(n654), .F(
        n83), .Z(dma_waddr[1]) );
  HS65_LS_IVX9 U37 ( .A(n85), .Z(n618) );
  HS65_LS_IVX9 U38 ( .A(state_cnt[0]), .Z(n443) );
  HS65_LS_AO222X4 U39 ( .A(\add_545/A[15] ), .B(n314), .C(\proc_in[MDATA][31] ), .D(n149), .E(dma_rp_new[15]), .F(n328), .Z(dma_wdata[47]) );
  HS65_LS_AND2X4 U40 ( .A(\proc_in[MCMD][0] ), .B(n590), .Z(n4) );
  HS65_LS_AND2X4 U41 ( .A(n609), .B(n53), .Z(n5) );
  HS65_LS_AND2X4 U42 ( .A(\add_545/A[14] ), .B(n73), .Z(n6) );
  HS65_LS_AND2X4 U43 ( .A(n132), .B(n410), .Z(n15) );
  HS65_LS_IVX18 U44 ( .A(n22), .Z(n116) );
  HS65_LS_IVX9 U45 ( .A(n573), .Z(n22) );
  HS65_LS_NAND3X13 U46 ( .A(n41), .B(n39), .C(n465), .Z(pkt_out[0]) );
  HS65_LS_NAND2X5 U47 ( .A(phitOut2[5]), .B(n471), .Z(n482) );
  HS65_LS_IVX9 U48 ( .A(n22), .Z(n114) );
  HS65_LS_NAND2X7 U49 ( .A(n105), .B(n461), .Z(n464) );
  HS65_LS_NOR2X13 U50 ( .A(n462), .B(n463), .Z(n105) );
  HS65_LS_AND2X27 U51 ( .A(n105), .B(n461), .Z(n28) );
  HS65_LS_NAND2X4 U52 ( .A(n448), .B(n459), .Z(n455) );
  HS65_LS_IVX2 U53 ( .A(n21), .Z(n120) );
  HS65_LS_OAI21X6 U54 ( .A(n572), .B(n113), .C(n571), .Z(pkt_out[34]) );
  HS65_LS_NAND2X4 U55 ( .A(state_cnt[0]), .B(state_cnt[1]), .Z(n456) );
  HS65_LS_NAND2X2 U56 ( .A(state_cnt[1]), .B(n443), .Z(n446) );
  HS65_LS_IVX18 U57 ( .A(n448), .Z(n34) );
  HS65_LS_NAND2X5 U58 ( .A(phitOut2[3]), .B(n28), .Z(n476) );
  HS65_LS_NAND2X5 U59 ( .A(phitOut2[13]), .B(n28), .Z(n506) );
  HS65_LS_NAND2X5 U60 ( .A(phitOut2[7]), .B(n28), .Z(n488) );
  HS65_LS_BFX53 U61 ( .A(n526), .Z(n27) );
  HS65_LS_OAI212X5 U62 ( .A(n112), .B(n502), .C(n501), .D(n27), .E(n500), .Z(
        pkt_out[11]) );
  HS65_LS_IVX2 U63 ( .A(n443), .Z(n26) );
  HS65_LS_IVX4 U64 ( .A(n34), .Z(n19) );
  HS65_LS_NAND2X4 U65 ( .A(phitOut2[4]), .B(n28), .Z(n479) );
  HS65_LS_NAND3X6 U66 ( .A(n118), .B(n449), .C(n450), .Z(n451) );
  HS65_LS_NAND2X4 U67 ( .A(phitOut2[19]), .B(n28), .Z(n524) );
  HS65_LS_AND2X18 U68 ( .A(n447), .B(n460), .Z(n24) );
  HS65_LS_IVX18 U69 ( .A(n20), .Z(n21) );
  HS65_LS_NAND2X21 U70 ( .A(n570), .B(n32), .Z(n573) );
  HS65_LS_IVX27 U71 ( .A(n573), .Z(n25) );
  HS65_LH_IVX2 U72 ( .A(n457), .Z(n23) );
  HS65_LS_IVX4 U73 ( .A(n460), .Z(n450) );
  HS65_LS_NAND2X14 U74 ( .A(n31), .B(n30), .Z(n32) );
  HS65_LS_IVX4 U75 ( .A(n455), .Z(n458) );
  HS65_LS_NAND2X4 U76 ( .A(phitOut2[0]), .B(n471), .Z(n465) );
  HS65_LS_NAND2X4 U77 ( .A(phitOut2[27]), .B(n28), .Z(n549) );
  HS65_LS_NAND2X4 U78 ( .A(phitOut2[30]), .B(n28), .Z(n558) );
  HS65_LS_NAND2X4 U79 ( .A(phitOut2[32]), .B(n28), .Z(n564) );
  HS65_LS_IVX9 U80 ( .A(n22), .Z(n117) );
  HS65_LS_OAI212X5 U81 ( .A(n113), .B(n523), .C(n27), .D(n522), .E(n521), .Z(
        pkt_out[18]) );
  HS65_LS_OAI212X5 U82 ( .A(n113), .B(n545), .C(n544), .D(n18), .E(n543), .Z(
        pkt_out[25]) );
  HS65_LS_IVX27 U83 ( .A(n461), .Z(n570) );
  HS65_LS_OAI212X3 U84 ( .A(n112), .B(n490), .C(n27), .D(n489), .E(n488), .Z(
        pkt_out[7]) );
  HS65_LS_OAI212X5 U85 ( .A(n112), .B(n527), .C(n27), .D(n525), .E(n524), .Z(
        pkt_out[19]) );
  HS65_LS_NAND2X7 U86 ( .A(state_cnt[0]), .B(n455), .Z(n453) );
  HS65_LS_AO33X9 U87 ( .A(n34), .B(n460), .C(n118), .D(\phase_next[1] ), .E(
        n446), .F(n445), .Z(n463) );
  HS65_LS_OAI212X5 U88 ( .A(n551), .B(n117), .C(n550), .D(n18), .E(n549), .Z(
        pkt_out[27]) );
  HS65_LS_OAI212X5 U89 ( .A(n113), .B(n470), .C(n27), .D(n469), .E(n468), .Z(
        pkt_out[1]) );
  HS65_LS_OAI212X5 U90 ( .A(n116), .B(n499), .C(n27), .D(n498), .E(n497), .Z(
        pkt_out[10]) );
  HS65_LS_NAND2X21 U91 ( .A(n35), .B(n37), .Z(n460) );
  HS65_LS_AOI33X2 U92 ( .A(n1), .B(n105), .C(phitOut2[34]), .D(n105), .E(
        phitOut0[34]), .F(n570), .Z(n571) );
  HS65_LH_MUX21I1X3 U93 ( .D0(n19), .D1(n449), .S0(n645), .Z(n315) );
  HS65_LS_OAI212X3 U94 ( .A(n112), .B(n508), .C(n27), .D(n507), .E(n506), .Z(
        pkt_out[13]) );
  HS65_LS_OR2X18 U95 ( .A(n112), .B(n467), .Z(n39) );
  HS65_LS_IVX18 U96 ( .A(n21), .Z(n459) );
  HS65_LS_IVX18 U97 ( .A(n454), .Z(n475) );
  HS65_LS_CBI4I1X11 U98 ( .A(n453), .B(n24), .C(n452), .D(n451), .Z(n454) );
  HS65_LS_IVX27 U99 ( .A(n464), .Z(n471) );
  HS65_LH_OAI212X3 U100 ( .A(n129), .B(n428), .C(n323), .D(n380), .E(n379), 
        .Z(mux_out[17]) );
  HS65_LS_OAI212X3 U101 ( .A(n129), .B(n429), .C(n323), .D(n382), .E(n381), 
        .Z(mux_out[18]) );
  HS65_LS_OAI212X5 U102 ( .A(n117), .B(n474), .C(n473), .D(n27), .E(n472), .Z(
        pkt_out[2]) );
  HS65_LH_IVX2 U103 ( .A(n446), .Z(n645) );
  HS65_LS_OAI212X3 U104 ( .A(n112), .B(n478), .C(n27), .D(n477), .E(n476), .Z(
        pkt_out[3]) );
  HS65_LS_NAND2X14 U105 ( .A(n448), .B(n459), .Z(n35) );
  HS65_LS_NAND2X14 U106 ( .A(n21), .B(n34), .Z(n37) );
  HS65_LS_NAND2X14 U107 ( .A(n475), .B(n109), .Z(n461) );
  HS65_LS_IVX9 U108 ( .A(state_cnt[1]), .Z(n447) );
  HS65_LS_BFX9 U109 ( .A(n330), .Z(n326) );
  HS65_LS_BFX9 U110 ( .A(n330), .Z(n325) );
  HS65_LS_BFX9 U111 ( .A(n311), .Z(n302) );
  HS65_LS_BFX9 U112 ( .A(n311), .Z(n303) );
  HS65_LS_BFX9 U113 ( .A(n293), .Z(n296) );
  HS65_LS_BFX9 U114 ( .A(n335), .Z(n353) );
  HS65_LS_BFX9 U115 ( .A(n334), .Z(n352) );
  HS65_LS_BFX9 U116 ( .A(n334), .Z(n351) );
  HS65_LH_MUXI21X2 U117 ( .D0(n452), .D1(n108), .S0(n645), .Z(n321) );
  HS65_LS_IVX9 U118 ( .A(n326), .Z(n312) );
  HS65_LS_IVX9 U119 ( .A(n326), .Z(n313) );
  HS65_LS_IVX9 U120 ( .A(n325), .Z(n314) );
  HS65_LS_IVX9 U121 ( .A(n325), .Z(n323) );
  HS65_LS_IVX9 U122 ( .A(n325), .Z(n324) );
  HS65_LS_AND2X4 U123 ( .A(n612), .B(n611), .Z(n42) );
  HS65_LS_AND2X4 U124 ( .A(n598), .B(n74), .Z(n43) );
  HS65_LS_AND2X4 U125 ( .A(n599), .B(n43), .Z(n44) );
  HS65_LS_AND2X4 U126 ( .A(n600), .B(n44), .Z(n45) );
  HS65_LS_AND2X4 U127 ( .A(n601), .B(n45), .Z(n46) );
  HS65_LS_AND2X4 U128 ( .A(n602), .B(n46), .Z(n47) );
  HS65_LS_AND2X4 U129 ( .A(n603), .B(n47), .Z(n48) );
  HS65_LS_AND2X4 U130 ( .A(n604), .B(n48), .Z(n49) );
  HS65_LS_AND2X4 U131 ( .A(n605), .B(n49), .Z(n50) );
  HS65_LS_AND2X4 U132 ( .A(n606), .B(n50), .Z(n51) );
  HS65_LS_AND2X4 U133 ( .A(n607), .B(n51), .Z(n52) );
  HS65_LS_AND2X4 U134 ( .A(n608), .B(n52), .Z(n53) );
  HS65_LS_AND2X4 U135 ( .A(n617), .B(n75), .Z(n54) );
  HS65_LS_AND2X4 U136 ( .A(n613), .B(n42), .Z(n55) );
  HS65_LS_AND2X4 U137 ( .A(n614), .B(n55), .Z(n56) );
  HS65_LS_AND2X4 U138 ( .A(n615), .B(n56), .Z(n57) );
  HS65_LS_AND2X4 U139 ( .A(\add_545/A[8] ), .B(n54), .Z(n58) );
  HS65_LS_AND2X4 U140 ( .A(\add_545/A[9] ), .B(n58), .Z(n59) );
  HS65_LS_AND2X4 U141 ( .A(\add_545/A[10] ), .B(n59), .Z(n62) );
  HS65_LS_AND2X4 U142 ( .A(\add_545/A[11] ), .B(n62), .Z(n64) );
  HS65_LS_AND2X4 U143 ( .A(\add_545/A[12] ), .B(n64), .Z(n72) );
  HS65_LS_AND2X4 U144 ( .A(\add_545/A[13] ), .B(n72), .Z(n73) );
  HS65_LS_AND2X4 U145 ( .A(n597), .B(n596), .Z(n74) );
  HS65_LS_AND2X4 U146 ( .A(n616), .B(n57), .Z(n75) );
  HS65_LS_BFX9 U147 ( .A(n329), .Z(n327) );
  HS65_LS_BFX9 U148 ( .A(n329), .Z(n328) );
  HS65_LS_IVX9 U149 ( .A(n302), .Z(n301) );
  HS65_LS_IVX9 U150 ( .A(n303), .Z(n300) );
  HS65_LS_IVX9 U151 ( .A(n303), .Z(n299) );
  HS65_LS_OAI21X3 U152 ( .A(n40), .B(n81), .C(n312), .Z(dma_wen[2]) );
  HS65_LS_NOR2AX3 U153 ( .A(n83), .B(n594), .Z(n40) );
  HS65_LS_IVX9 U154 ( .A(n86), .Z(n594) );
  HS65_LSS_XNOR2X6 U155 ( .A(n94), .B(\sub_544/A[10] ), .Z(dma_cnt_new[10]) );
  HS65_LSS_XNOR2X6 U156 ( .A(n88), .B(\sub_544/A[5] ), .Z(dma_cnt_new[5]) );
  HS65_LSS_XNOR2X6 U157 ( .A(n93), .B(\sub_544/A[9] ), .Z(dma_cnt_new[9]) );
  HS65_LSS_XNOR2X6 U158 ( .A(n87), .B(\sub_544/A[4] ), .Z(dma_cnt_new[4]) );
  HS65_LSS_XNOR2X6 U159 ( .A(n91), .B(\sub_544/A[8] ), .Z(dma_cnt_new[8]) );
  HS65_LS_NOR4ABX2 U160 ( .A(n102), .B(n103), .C(n65), .D(dma_cnt_new[13]), 
        .Z(n100) );
  HS65_LSS_XOR2X6 U161 ( .A(n90), .B(\sub_544/A[7] ), .Z(n77) );
  HS65_LSS_XOR2X6 U162 ( .A(n84), .B(\sub_544/A[3] ), .Z(n78) );
  HS65_LSS_XOR2X6 U163 ( .A(n89), .B(\sub_544/A[6] ), .Z(n79) );
  HS65_LS_IVX9 U164 ( .A(n9), .Z(\add_545/A[8] ) );
  HS65_LS_IVX9 U165 ( .A(n8), .Z(\add_545/A[9] ) );
  HS65_LS_IVX9 U166 ( .A(n7), .Z(\add_545/A[10] ) );
  HS65_LS_IVX9 U167 ( .A(n14), .Z(\add_545/A[11] ) );
  HS65_LS_IVX9 U168 ( .A(n13), .Z(\add_545/A[12] ) );
  HS65_LS_IVX9 U169 ( .A(n12), .Z(\add_545/A[13] ) );
  HS65_LS_IVX9 U170 ( .A(n11), .Z(\add_545/A[14] ) );
  HS65_LS_BFX9 U171 ( .A(n104), .Z(n329) );
  HS65_LS_BFX9 U172 ( .A(n104), .Z(n330) );
  HS65_LSS_XOR2X6 U173 ( .A(\sub_544/A[1] ), .B(\sub_544/A[2] ), .Z(n80) );
  HS65_LS_OR2X9 U174 ( .A(\sub_544/A[2] ), .B(\sub_544/A[1] ), .Z(n84) );
  HS65_LS_OR2X9 U175 ( .A(\sub_544/A[3] ), .B(n84), .Z(n87) );
  HS65_LS_OR2X9 U176 ( .A(\sub_544/A[4] ), .B(n87), .Z(n88) );
  HS65_LS_OR2X9 U177 ( .A(\sub_544/A[5] ), .B(n88), .Z(n89) );
  HS65_LS_OR2X9 U178 ( .A(\sub_544/A[6] ), .B(n89), .Z(n90) );
  HS65_LS_OR2X9 U179 ( .A(\sub_544/A[7] ), .B(n90), .Z(n91) );
  HS65_LS_OR2X9 U180 ( .A(\sub_544/A[8] ), .B(n91), .Z(n93) );
  HS65_LS_OR2X9 U181 ( .A(\sub_544/A[9] ), .B(n93), .Z(n94) );
  HS65_LS_OR2X9 U182 ( .A(\sub_544/A[10] ), .B(n94), .Z(n95) );
  HS65_LS_OR2X9 U183 ( .A(\sub_544/A[11] ), .B(n95), .Z(n101) );
  HS65_LSS_XOR2X6 U184 ( .A(n95), .B(\sub_544/A[11] ), .Z(n102) );
  HS65_LSS_XOR2X6 U185 ( .A(n101), .B(\sub_544/A[12] ), .Z(n103) );
  HS65_LS_BFX9 U186 ( .A(n137), .Z(n138) );
  HS65_LS_BFX9 U187 ( .A(n137), .Z(n139) );
  HS65_LS_BFX9 U188 ( .A(n140), .Z(n144) );
  HS65_LS_BFX9 U189 ( .A(n140), .Z(n142) );
  HS65_LS_BFX9 U190 ( .A(n140), .Z(n149) );
  HS65_LS_IVX9 U191 ( .A(n296), .Z(n294) );
  HS65_LS_IVX9 U192 ( .A(n296), .Z(n295) );
  HS65_LS_BFX9 U193 ( .A(n311), .Z(n304) );
  HS65_LS_BFX9 U194 ( .A(n311), .Z(n306) );
  HS65_LS_BFX9 U195 ( .A(n311), .Z(n305) );
  HS65_LS_BFX9 U196 ( .A(n311), .Z(n310) );
  HS65_LS_BFX9 U197 ( .A(n127), .Z(n128) );
  HS65_LS_BFX9 U198 ( .A(n127), .Z(n129) );
  HS65_LS_BFX9 U199 ( .A(n15), .Z(n122) );
  HS65_LS_BFX9 U200 ( .A(n15), .Z(n124) );
  HS65_LS_BFX9 U201 ( .A(n127), .Z(n130) );
  HS65_LS_BFX9 U202 ( .A(n15), .Z(n125) );
  HS65_LS_IVX9 U203 ( .A(n81), .Z(n650) );
  HS65_LS_IVX9 U204 ( .A(\proc_out[SRESP] ), .Z(n331) );
  HS65_LS_IVX9 U205 ( .A(n353), .Z(n344) );
  HS65_LS_IVX9 U206 ( .A(n353), .Z(n343) );
  HS65_LS_IVX9 U207 ( .A(n353), .Z(n347) );
  HS65_LS_IVX9 U208 ( .A(n353), .Z(n346) );
  HS65_LS_IVX9 U209 ( .A(n353), .Z(n345) );
  HS65_LS_IVX9 U210 ( .A(n352), .Z(n342) );
  HS65_LS_IVX9 U211 ( .A(n352), .Z(n341) );
  HS65_LS_IVX9 U212 ( .A(n352), .Z(n339) );
  HS65_LS_IVX9 U213 ( .A(n352), .Z(n338) );
  HS65_LS_IVX9 U214 ( .A(n352), .Z(n337) );
  HS65_LS_IVX9 U215 ( .A(n352), .Z(n340) );
  HS65_LS_IVX9 U216 ( .A(n354), .Z(n350) );
  HS65_LS_IVX9 U217 ( .A(n354), .Z(n349) );
  HS65_LS_IVX9 U218 ( .A(n354), .Z(n348) );
  HS65_LS_IVX9 U219 ( .A(n351), .Z(n336) );
  HS65_LS_NOR2X6 U220 ( .A(n354), .B(n9), .Z(\spm_out[MADDR][7] ) );
  HS65_LS_NOR2X6 U221 ( .A(n354), .B(n8), .Z(\spm_out[MADDR][8] ) );
  HS65_LS_NOR2X6 U222 ( .A(n354), .B(n7), .Z(\spm_out[MADDR][9] ) );
  HS65_LS_NOR2X6 U223 ( .A(n354), .B(n14), .Z(\spm_out[MADDR][10] ) );
  HS65_LS_NOR2X6 U224 ( .A(n354), .B(n13), .Z(\spm_out[MADDR][11] ) );
  HS65_LS_NOR2X6 U225 ( .A(n354), .B(n12), .Z(\spm_out[MADDR][12] ) );
  HS65_LS_NOR2X6 U226 ( .A(n354), .B(n11), .Z(\spm_out[MADDR][13] ) );
  HS65_LS_NOR2X6 U227 ( .A(n354), .B(n10), .Z(\spm_out[MADDR][14] ) );
  HS65_LS_NOR2X6 U228 ( .A(n331), .B(n640), .Z(\proc_out[SDATA][0] ) );
  HS65_LS_NOR2X6 U229 ( .A(n331), .B(n639), .Z(\proc_out[SDATA][1] ) );
  HS65_LS_NOR2X6 U230 ( .A(n331), .B(n638), .Z(\proc_out[SDATA][2] ) );
  HS65_LS_NOR2X6 U231 ( .A(n16), .B(n637), .Z(\proc_out[SDATA][3] ) );
  HS65_LS_NOR2X6 U232 ( .A(n331), .B(n636), .Z(\proc_out[SDATA][4] ) );
  HS65_LS_NOR2X6 U233 ( .A(n16), .B(n635), .Z(\proc_out[SDATA][5] ) );
  HS65_LS_NOR2X6 U234 ( .A(n16), .B(n634), .Z(\proc_out[SDATA][6] ) );
  HS65_LS_NOR2X6 U235 ( .A(n16), .B(n633), .Z(\proc_out[SDATA][7] ) );
  HS65_LS_NOR2X6 U236 ( .A(n331), .B(n632), .Z(\proc_out[SDATA][8] ) );
  HS65_LS_NOR2X6 U237 ( .A(n331), .B(n631), .Z(\proc_out[SDATA][9] ) );
  HS65_LS_NOR2X6 U238 ( .A(n331), .B(n630), .Z(\proc_out[SDATA][10] ) );
  HS65_LS_NOR2X6 U239 ( .A(n331), .B(n629), .Z(\proc_out[SDATA][11] ) );
  HS65_LS_NOR2X6 U240 ( .A(n331), .B(n628), .Z(\proc_out[SDATA][12] ) );
  HS65_LS_NOR2X6 U241 ( .A(n331), .B(n627), .Z(\proc_out[SDATA][13] ) );
  HS65_LS_NOR2X6 U242 ( .A(n331), .B(n626), .Z(\proc_out[SDATA][14] ) );
  HS65_LS_NOR2X6 U243 ( .A(n331), .B(n625), .Z(\proc_out[SDATA][15] ) );
  HS65_LS_AND3X9 U244 ( .A(dma_rdata[63]), .B(n642), .C(n139), .Z(n104) );
  HS65_LS_OAI222X2 U245 ( .A(n326), .B(n131), .C(n92), .D(n672), .E(n312), .F(
        n131), .Z(dma_wdata[48]) );
  HS65_LS_NOR2X6 U246 ( .A(n40), .B(n82), .Z(dma_wen[0]) );
  HS65_LS_OAI222X2 U247 ( .A(n326), .B(n126), .C(n92), .D(n669), .E(n312), .F(
        n78), .Z(dma_wdata[51]) );
  HS65_LS_OAI222X2 U248 ( .A(n326), .B(n123), .C(n92), .D(n668), .E(n312), .F(
        n624), .Z(dma_wdata[52]) );
  HS65_LS_IVX9 U249 ( .A(dma_cnt_new[4]), .Z(n624) );
  HS65_LS_OAI222X2 U250 ( .A(n326), .B(n121), .C(n665), .D(n92), .E(n312), .F(
        n77), .Z(dma_wdata[55]) );
  HS65_LS_OAI222X2 U251 ( .A(n326), .B(n119), .C(n664), .D(n92), .E(n312), .F(
        n622), .Z(dma_wdata[56]) );
  HS65_LS_IVX9 U252 ( .A(dma_cnt_new[8]), .Z(n622) );
  HS65_LS_OAI222X2 U253 ( .A(n326), .B(n115), .C(n92), .D(n662), .E(n313), .F(
        n620), .Z(dma_wdata[58]) );
  HS65_LS_IVX9 U254 ( .A(dma_cnt_new[10]), .Z(n620) );
  HS65_LS_OAI222X2 U255 ( .A(n325), .B(n110), .C(n92), .D(n660), .E(n313), .F(
        n103), .Z(dma_wdata[60]) );
  HS65_LS_OAI222X2 U256 ( .A(n326), .B(n107), .C(n92), .D(n659), .E(n312), .F(
        n619), .Z(dma_wdata[61]) );
  HS65_LS_IVX9 U257 ( .A(dma_cnt_new[13]), .Z(n619) );
  HS65_LS_OAI222X2 U258 ( .A(n326), .B(n65), .C(n92), .D(n671), .E(n312), .F(
        \sub_544/A[1] ), .Z(dma_wdata[49]) );
  HS65_LS_OAI222X2 U259 ( .A(n326), .B(n66), .C(n92), .D(n670), .E(n312), .F(
        n80), .Z(dma_wdata[50]) );
  HS65_LS_OAI222X2 U260 ( .A(n326), .B(n67), .C(n92), .D(n667), .E(n312), .F(
        n623), .Z(dma_wdata[53]) );
  HS65_LS_IVX9 U261 ( .A(dma_cnt_new[5]), .Z(n623) );
  HS65_LS_OAI222X2 U262 ( .A(n326), .B(n68), .C(n666), .D(n92), .E(n312), .F(
        n79), .Z(dma_wdata[54]) );
  HS65_LS_OAI222X2 U263 ( .A(n326), .B(n69), .C(n663), .D(n92), .E(n312), .F(
        n621), .Z(dma_wdata[57]) );
  HS65_LS_IVX9 U264 ( .A(dma_cnt_new[9]), .Z(n621) );
  HS65_LS_OAI222X2 U265 ( .A(n326), .B(n70), .C(n92), .D(n661), .E(n312), .F(
        n102), .Z(dma_wdata[59]) );
  HS65_LS_OAI212X5 U266 ( .A(n92), .B(n658), .C(n85), .D(n642), .E(n96), .Z(
        dma_wdata[62]) );
  HS65_LS_NAND4ABX3 U267 ( .A(n97), .B(n98), .C(n99), .D(n100), .Z(n96) );
  HS65_LS_NAND4ABX3 U268 ( .A(dma_cnt_new[5]), .B(dma_cnt_new[4]), .C(n80), 
        .D(n78), .Z(n98) );
  HS65_LS_NAND4ABX3 U269 ( .A(dma_cnt_new[9]), .B(dma_cnt_new[8]), .C(n79), 
        .D(n77), .Z(n97) );
  HS65_LS_NAND2X7 U270 ( .A(n649), .B(n4), .Z(n86) );
  HS65_LS_OAI21X3 U271 ( .A(n40), .B(n71), .C(n312), .Z(dma_wen[1]) );
  HS65_LH_NAND2X2 U272 ( .A(n360), .B(n444), .Z(n590) );
  HS65_LSS_XNOR2X6 U273 ( .A(n107), .B(n111), .Z(dma_cnt_new[13]) );
  HS65_LS_NOR2X6 U274 ( .A(\sub_544/A[12] ), .B(n101), .Z(n111) );
  HS65_LS_NOR3X4 U275 ( .A(n312), .B(dma_cnt_new[10]), .C(dma_cnt_new[0]), .Z(
        n99) );
  HS65_LS_IVX9 U276 ( .A(n131), .Z(dma_cnt_new[0]) );
  HS65_LS_IVX9 U277 ( .A(n65), .Z(\sub_544/A[1] ) );
  HS65_LS_NAND2X7 U278 ( .A(dma_rdata[40]), .B(n139), .Z(n9) );
  HS65_LS_NAND2X7 U279 ( .A(dma_rdata[41]), .B(n139), .Z(n8) );
  HS65_LS_NAND2X7 U280 ( .A(dma_rdata[42]), .B(n138), .Z(n7) );
  HS65_LS_NAND2X7 U281 ( .A(dma_rdata[43]), .B(n139), .Z(n14) );
  HS65_LS_NAND2X7 U282 ( .A(dma_rdata[44]), .B(n138), .Z(n13) );
  HS65_LS_NAND2X7 U283 ( .A(dma_rdata[45]), .B(n139), .Z(n12) );
  HS65_LS_NAND2X7 U284 ( .A(dma_rdata[46]), .B(n139), .Z(n11) );
  HS65_LS_IVX9 U285 ( .A(n126), .Z(\sub_544/A[3] ) );
  HS65_LS_IVX9 U286 ( .A(n123), .Z(\sub_544/A[4] ) );
  HS65_LS_IVX9 U287 ( .A(n121), .Z(\sub_544/A[7] ) );
  HS65_LS_IVX9 U288 ( .A(n119), .Z(\sub_544/A[8] ) );
  HS65_LS_IVX9 U289 ( .A(n115), .Z(\sub_544/A[10] ) );
  HS65_LS_IVX9 U290 ( .A(n110), .Z(\sub_544/A[12] ) );
  HS65_LS_IVX9 U291 ( .A(n66), .Z(\sub_544/A[2] ) );
  HS65_LS_IVX9 U292 ( .A(n67), .Z(\sub_544/A[5] ) );
  HS65_LS_IVX9 U293 ( .A(n68), .Z(\sub_544/A[6] ) );
  HS65_LS_IVX9 U294 ( .A(n69), .Z(\sub_544/A[9] ) );
  HS65_LS_IVX9 U295 ( .A(n70), .Z(\sub_544/A[11] ) );
  HS65_LS_BFX9 U296 ( .A(n618), .Z(n137) );
  HS65_LS_BFX9 U297 ( .A(n135), .Z(n140) );
  HS65_LS_NOR2AX3 U298 ( .A(n4), .B(n71), .Z(n135) );
  HS65_LS_BFX9 U299 ( .A(n409), .Z(n127) );
  HS65_LS_OAI22X6 U300 ( .A(n85), .B(n640), .C(n86), .D(n672), .Z(dma_wdata[0]) );
  HS65_LS_OAI22X6 U301 ( .A(n85), .B(n639), .C(n86), .D(n671), .Z(dma_wdata[1]) );
  HS65_LS_OAI22X6 U302 ( .A(n85), .B(n638), .C(n86), .D(n670), .Z(dma_wdata[2]) );
  HS65_LS_OAI22X6 U303 ( .A(n85), .B(n637), .C(n86), .D(n669), .Z(dma_wdata[3]) );
  HS65_LS_OAI22X6 U304 ( .A(n85), .B(n636), .C(n86), .D(n668), .Z(dma_wdata[4]) );
  HS65_LS_OAI22X6 U305 ( .A(n85), .B(n635), .C(n86), .D(n667), .Z(dma_wdata[5]) );
  HS65_LS_OAI22X6 U306 ( .A(n85), .B(n634), .C(n86), .D(n666), .Z(dma_wdata[6]) );
  HS65_LS_OAI22X6 U307 ( .A(n85), .B(n633), .C(n86), .D(n665), .Z(dma_wdata[7]) );
  HS65_LS_OAI22X6 U308 ( .A(n85), .B(n632), .C(n86), .D(n664), .Z(dma_wdata[8]) );
  HS65_LS_OAI22X6 U309 ( .A(n85), .B(n631), .C(n86), .D(n663), .Z(dma_wdata[9]) );
  HS65_LS_OAI22X6 U310 ( .A(n85), .B(n630), .C(n86), .D(n662), .Z(
        dma_wdata[10]) );
  HS65_LS_OAI22X6 U311 ( .A(n85), .B(n629), .C(n86), .D(n661), .Z(
        dma_wdata[11]) );
  HS65_LS_OAI22X6 U312 ( .A(n85), .B(n628), .C(n86), .D(n660), .Z(
        dma_wdata[12]) );
  HS65_LS_OAI22X6 U313 ( .A(n85), .B(n627), .C(n86), .D(n659), .Z(
        dma_wdata[13]) );
  HS65_LS_OAI22X6 U314 ( .A(n85), .B(n626), .C(n86), .D(n658), .Z(
        dma_wdata[14]) );
  HS65_LS_OAI22X6 U315 ( .A(n85), .B(n625), .C(n86), .D(n657), .Z(
        dma_wdata[15]) );
  HS65_LS_OAI22X6 U316 ( .A(n85), .B(n641), .C(n92), .D(n657), .Z(
        dma_wdata[63]) );
  HS65_LS_IVX9 U317 ( .A(dma_rdata[63]), .Z(n641) );
  HS65_LS_OAI21X3 U318 ( .A(n649), .B(n141), .C(n356), .Z(n591) );
  HS65_LH_OAI21X2 U319 ( .A(n82), .B(n591), .C(n360), .Z(dma_ren[0]) );
  HS65_LH_OAI21X2 U320 ( .A(n71), .B(n591), .C(n360), .Z(dma_ren[1]) );
  HS65_LH_OAI21X2 U321 ( .A(n81), .B(n591), .C(n360), .Z(dma_ren[2]) );
  HS65_LS_NAND2X7 U322 ( .A(n650), .B(n4), .Z(n92) );
  HS65_LS_IVX9 U323 ( .A(n63), .Z(n646) );
  HS65_LS_NAND2X7 U324 ( .A(dma_rdata[47]), .B(n139), .Z(n10) );
  HS65_LS_IVX9 U325 ( .A(dma_rdata[0]), .Z(n640) );
  HS65_LS_IVX9 U326 ( .A(dma_rdata[1]), .Z(n639) );
  HS65_LS_IVX9 U327 ( .A(dma_rdata[2]), .Z(n638) );
  HS65_LS_IVX9 U328 ( .A(dma_rdata[3]), .Z(n637) );
  HS65_LS_IVX9 U329 ( .A(dma_rdata[4]), .Z(n636) );
  HS65_LS_IVX9 U330 ( .A(dma_rdata[5]), .Z(n635) );
  HS65_LS_IVX9 U331 ( .A(dma_rdata[6]), .Z(n634) );
  HS65_LS_IVX9 U332 ( .A(dma_rdata[7]), .Z(n633) );
  HS65_LS_IVX9 U333 ( .A(dma_rdata[8]), .Z(n632) );
  HS65_LS_IVX9 U334 ( .A(dma_rdata[9]), .Z(n631) );
  HS65_LS_IVX9 U335 ( .A(dma_rdata[10]), .Z(n630) );
  HS65_LS_IVX9 U336 ( .A(dma_rdata[11]), .Z(n629) );
  HS65_LS_IVX9 U337 ( .A(dma_rdata[12]), .Z(n628) );
  HS65_LS_IVX9 U338 ( .A(dma_rdata[13]), .Z(n627) );
  HS65_LS_IVX9 U339 ( .A(dma_rdata[14]), .Z(n626) );
  HS65_LS_IVX9 U340 ( .A(dma_rdata[15]), .Z(n625) );
  HS65_LS_BFX9 U341 ( .A(n293), .Z(n297) );
  HS65_LS_IVX9 U342 ( .A(n60), .Z(n311) );
  HS65_LS_BFX9 U343 ( .A(n293), .Z(n298) );
  HS65_LS_NAND3X5 U344 ( .A(n136), .B(n574), .C(n336), .Z(n589) );
  HS65_LS_IVX9 U345 ( .A(n82), .Z(n649) );
  HS65_LS_NAND2X7 U346 ( .A(n81), .B(n71), .Z(n141) );
  HS65_LS_NAND2X7 U347 ( .A(n146), .B(n656), .Z(n81) );
  HS65_LS_BFX9 U348 ( .A(n333), .Z(\proc_out[SRESP] ) );
  HS65_LS_IVX9 U349 ( .A(n16), .Z(n333) );
  HS65_LS_BFX9 U350 ( .A(n335), .Z(n354) );
  HS65_LS_IVX9 U351 ( .A(n38), .Z(n648) );
  HS65_LS_NOR2AX3 U352 ( .A(dma_rdata[16]), .B(n16), .Z(\proc_out[SDATA][16] )
         );
  HS65_LS_NOR2AX3 U353 ( .A(dma_rdata[17]), .B(n16), .Z(\proc_out[SDATA][17] )
         );
  HS65_LS_NOR2AX3 U354 ( .A(dma_rdata[18]), .B(n16), .Z(\proc_out[SDATA][18] )
         );
  HS65_LS_NOR2AX3 U355 ( .A(dma_rdata[19]), .B(n16), .Z(\proc_out[SDATA][19] )
         );
  HS65_LS_NOR2AX3 U356 ( .A(dma_rdata[20]), .B(n16), .Z(\proc_out[SDATA][20] )
         );
  HS65_LS_NOR2AX3 U357 ( .A(dma_rdata[21]), .B(n16), .Z(\proc_out[SDATA][21] )
         );
  HS65_LS_NOR2AX3 U358 ( .A(dma_rdata[22]), .B(n16), .Z(\proc_out[SDATA][22] )
         );
  HS65_LS_NOR2AX3 U359 ( .A(dma_rdata[23]), .B(n16), .Z(\proc_out[SDATA][23] )
         );
  HS65_LS_NOR2AX3 U360 ( .A(dma_rdata[24]), .B(n16), .Z(\proc_out[SDATA][24] )
         );
  HS65_LS_NOR2AX3 U361 ( .A(dma_rdata[25]), .B(n16), .Z(\proc_out[SDATA][25] )
         );
  HS65_LS_NOR2AX3 U362 ( .A(dma_rdata[26]), .B(n331), .Z(\proc_out[SDATA][26] ) );
  HS65_LS_NOR2AX3 U363 ( .A(dma_rdata[27]), .B(n16), .Z(\proc_out[SDATA][27] )
         );
  HS65_LS_NOR2AX3 U364 ( .A(dma_rdata[28]), .B(n16), .Z(\proc_out[SDATA][28] )
         );
  HS65_LS_NOR2AX3 U365 ( .A(dma_rdata[29]), .B(n331), .Z(\proc_out[SDATA][29] ) );
  HS65_LS_NOR2AX3 U366 ( .A(dma_rdata[30]), .B(n16), .Z(\proc_out[SDATA][30] )
         );
  HS65_LS_NOR2AX3 U367 ( .A(dma_rdata[31]), .B(n16), .Z(\proc_out[SDATA][31] )
         );
  HS65_LS_IVX9 U368 ( .A(n71), .Z(n651) );
  HS65_LS_AOI22X6 U369 ( .A(\proc_in[MADDR][1] ), .B(n649), .C(
        \proc_in[MADDR][2] ), .D(n141), .Z(n143) );
  HS65_LS_AOI22X6 U370 ( .A(\proc_in[MADDR][0] ), .B(n649), .C(
        \proc_in[MADDR][1] ), .D(n141), .Z(n145) );
  HS65_LS_IVX9 U371 ( .A(\proc_in[MADDR][2] ), .Z(n654) );
  HS65_LS_OAI212X5 U372 ( .A(n113), .B(n539), .C(n3), .D(n538), .E(n537), .Z(
        pkt_out[23]) );
  HS65_LS_OAI212X5 U373 ( .A(n113), .B(n542), .C(n3), .D(n541), .E(n540), .Z(
        pkt_out[24]) );
  HS65_LH_MUXI21X2 U374 ( .D0(n307), .D1(n106), .S0(n645), .Z(n320) );
  HS65_LS_NOR2X6 U375 ( .A(slt_entry[0]), .B(n314), .Z(n106) );
  HS65_LS_NOR2X6 U376 ( .A(slt_entry[1]), .B(n314), .Z(n108) );
  HS65_LS_MX41X7 U377 ( .D0(n593), .S0(n327), .D1(n593), .S1(n313), .D2(
        \proc_in[MDATA][16] ), .S2(n594), .D3(n142), .S3(\proc_in[MDATA][0] ), 
        .Z(dma_wdata[16]) );
  HS65_LS_MX41X7 U378 ( .D0(n380), .S0(n326), .D1(n596), .S1(n313), .D2(
        \proc_in[MDATA][17] ), .S2(n594), .D3(n142), .S3(\proc_in[MDATA][1] ), 
        .Z(dma_wdata[17]) );
  HS65_LS_MX41X7 U379 ( .D0(dma_wp_new[2]), .S0(n326), .D1(n597), .S1(n313), 
        .D2(\proc_in[MDATA][18] ), .S2(n594), .D3(n142), .S3(
        \proc_in[MDATA][2] ), .Z(dma_wdata[18]) );
  HS65_LSS_XOR2X6 U380 ( .A(n596), .B(n597), .Z(dma_wp_new[2]) );
  HS65_LS_MX41X7 U381 ( .D0(dma_wp_new[3]), .S0(n326), .D1(n598), .S1(n313), 
        .D2(\proc_in[MDATA][19] ), .S2(n594), .D3(n142), .S3(
        \proc_in[MDATA][3] ), .Z(dma_wdata[19]) );
  HS65_LSS_XOR2X6 U382 ( .A(n74), .B(n598), .Z(dma_wp_new[3]) );
  HS65_LS_MX41X7 U383 ( .D0(dma_wp_new[4]), .S0(n326), .D1(n599), .S1(n313), 
        .D2(\proc_in[MDATA][20] ), .S2(n594), .D3(n142), .S3(
        \proc_in[MDATA][4] ), .Z(dma_wdata[20]) );
  HS65_LSS_XOR2X6 U384 ( .A(n43), .B(n599), .Z(dma_wp_new[4]) );
  HS65_LS_MX41X7 U385 ( .D0(dma_wp_new[5]), .S0(n326), .D1(n600), .S1(n313), 
        .D2(\proc_in[MDATA][21] ), .S2(n594), .D3(n142), .S3(
        \proc_in[MDATA][5] ), .Z(dma_wdata[21]) );
  HS65_LSS_XOR2X6 U386 ( .A(n44), .B(n600), .Z(dma_wp_new[5]) );
  HS65_LS_MX41X7 U387 ( .D0(dma_wp_new[6]), .S0(n327), .D1(n601), .S1(n313), 
        .D2(\proc_in[MDATA][22] ), .S2(n594), .D3(n142), .S3(
        \proc_in[MDATA][6] ), .Z(dma_wdata[22]) );
  HS65_LSS_XOR2X6 U388 ( .A(n45), .B(n601), .Z(dma_wp_new[6]) );
  HS65_LS_MX41X7 U389 ( .D0(dma_wp_new[7]), .S0(n327), .D1(n602), .S1(n313), 
        .D2(\proc_in[MDATA][23] ), .S2(n594), .D3(n142), .S3(
        \proc_in[MDATA][7] ), .Z(dma_wdata[23]) );
  HS65_LSS_XOR2X6 U390 ( .A(n46), .B(n602), .Z(dma_wp_new[7]) );
  HS65_LS_MX41X7 U391 ( .D0(dma_wp_new[8]), .S0(n327), .D1(n603), .S1(n313), 
        .D2(\proc_in[MDATA][24] ), .S2(n594), .D3(n142), .S3(
        \proc_in[MDATA][8] ), .Z(dma_wdata[24]) );
  HS65_LSS_XOR2X6 U392 ( .A(n47), .B(n603), .Z(dma_wp_new[8]) );
  HS65_LS_MX41X7 U393 ( .D0(dma_wp_new[9]), .S0(n327), .D1(n604), .S1(n313), 
        .D2(\proc_in[MDATA][25] ), .S2(n594), .D3(n142), .S3(
        \proc_in[MDATA][9] ), .Z(dma_wdata[25]) );
  HS65_LSS_XOR2X6 U394 ( .A(n48), .B(n604), .Z(dma_wp_new[9]) );
  HS65_LS_MX41X7 U395 ( .D0(dma_wp_new[10]), .S0(n327), .D1(n605), .S1(n313), 
        .D2(\proc_in[MDATA][26] ), .S2(n594), .D3(n142), .S3(
        \proc_in[MDATA][10] ), .Z(dma_wdata[26]) );
  HS65_LSS_XOR2X6 U396 ( .A(n49), .B(n605), .Z(dma_wp_new[10]) );
  HS65_LS_MX41X7 U397 ( .D0(dma_wp_new[11]), .S0(n327), .D1(n606), .S1(n313), 
        .D2(\proc_in[MDATA][27] ), .S2(n594), .D3(n142), .S3(
        \proc_in[MDATA][11] ), .Z(dma_wdata[27]) );
  HS65_LSS_XOR2X6 U398 ( .A(n50), .B(n606), .Z(dma_wp_new[11]) );
  HS65_LS_MX41X7 U399 ( .D0(dma_wp_new[12]), .S0(n327), .D1(n607), .S1(n313), 
        .D2(\proc_in[MDATA][28] ), .S2(n594), .D3(n144), .S3(
        \proc_in[MDATA][12] ), .Z(dma_wdata[28]) );
  HS65_LSS_XOR2X6 U400 ( .A(n51), .B(n607), .Z(dma_wp_new[12]) );
  HS65_LS_MX41X7 U401 ( .D0(dma_wp_new[13]), .S0(n327), .D1(n608), .S1(n313), 
        .D2(\proc_in[MDATA][29] ), .S2(n594), .D3(n144), .S3(
        \proc_in[MDATA][13] ), .Z(dma_wdata[29]) );
  HS65_LSS_XOR2X6 U402 ( .A(n52), .B(n608), .Z(dma_wp_new[13]) );
  HS65_LS_MX41X7 U403 ( .D0(dma_wp_new[14]), .S0(n327), .D1(n609), .S1(n313), 
        .D2(\proc_in[MDATA][30] ), .S2(n594), .D3(n144), .S3(
        \proc_in[MDATA][14] ), .Z(dma_wdata[30]) );
  HS65_LSS_XOR2X6 U404 ( .A(n53), .B(n609), .Z(dma_wp_new[14]) );
  HS65_LS_MX41X7 U405 ( .D0(dma_wp_new[15]), .S0(n327), .D1(n610), .S1(n313), 
        .D2(\proc_in[MDATA][31] ), .S2(n594), .D3(n144), .S3(
        \proc_in[MDATA][15] ), .Z(dma_wdata[31]) );
  HS65_LSS_XOR2X6 U406 ( .A(n610), .B(n5), .Z(dma_wp_new[15]) );
  HS65_LS_AO222X4 U407 ( .A(n611), .B(n314), .C(\proc_in[MDATA][17] ), .D(n144), .E(n576), .F(n327), .Z(dma_wdata[33]) );
  HS65_LS_AO222X4 U408 ( .A(n612), .B(n314), .C(\proc_in[MDATA][18] ), .D(n144), .E(dma_rp_new[2]), .F(n327), .Z(dma_wdata[34]) );
  HS65_LSS_XOR2X6 U409 ( .A(n611), .B(n612), .Z(dma_rp_new[2]) );
  HS65_LS_AO222X4 U410 ( .A(n613), .B(n314), .C(\proc_in[MDATA][19] ), .D(n144), .E(dma_rp_new[3]), .F(n327), .Z(dma_wdata[35]) );
  HS65_LSS_XOR2X6 U411 ( .A(n42), .B(n613), .Z(dma_rp_new[3]) );
  HS65_LS_AO222X4 U412 ( .A(n614), .B(n313), .C(\proc_in[MDATA][20] ), .D(n144), .E(dma_rp_new[4]), .F(n327), .Z(dma_wdata[36]) );
  HS65_LSS_XOR2X6 U413 ( .A(n55), .B(n614), .Z(dma_rp_new[4]) );
  HS65_LS_AO222X4 U414 ( .A(n615), .B(n314), .C(\proc_in[MDATA][21] ), .D(n144), .E(dma_rp_new[5]), .F(n327), .Z(dma_wdata[37]) );
  HS65_LSS_XOR2X6 U415 ( .A(n56), .B(n615), .Z(dma_rp_new[5]) );
  HS65_LS_AO222X4 U416 ( .A(n616), .B(n314), .C(\proc_in[MDATA][22] ), .D(n144), .E(dma_rp_new[6]), .F(n327), .Z(dma_wdata[38]) );
  HS65_LSS_XOR2X6 U417 ( .A(n57), .B(n616), .Z(dma_rp_new[6]) );
  HS65_LS_AO222X4 U418 ( .A(n617), .B(n314), .C(\proc_in[MDATA][23] ), .D(n144), .E(dma_rp_new[7]), .F(n327), .Z(dma_wdata[39]) );
  HS65_LSS_XOR2X6 U419 ( .A(n75), .B(n617), .Z(dma_rp_new[7]) );
  HS65_LS_AO222X4 U420 ( .A(\add_545/A[8] ), .B(n314), .C(\proc_in[MDATA][24] ), .D(n144), .E(dma_rp_new[8]), .F(n327), .Z(dma_wdata[40]) );
  HS65_LSS_XOR2X6 U421 ( .A(n54), .B(\add_545/A[8] ), .Z(dma_rp_new[8]) );
  HS65_LS_AO222X4 U422 ( .A(\add_545/A[9] ), .B(n314), .C(\proc_in[MDATA][25] ), .D(n149), .E(dma_rp_new[9]), .F(n328), .Z(dma_wdata[41]) );
  HS65_LSS_XOR2X6 U423 ( .A(n58), .B(\add_545/A[9] ), .Z(dma_rp_new[9]) );
  HS65_LS_AO222X4 U424 ( .A(\add_545/A[10] ), .B(n314), .C(
        \proc_in[MDATA][26] ), .D(n149), .E(dma_rp_new[10]), .F(n328), .Z(
        dma_wdata[42]) );
  HS65_LSS_XOR2X6 U425 ( .A(n59), .B(\add_545/A[10] ), .Z(dma_rp_new[10]) );
  HS65_LS_AO222X4 U426 ( .A(\add_545/A[11] ), .B(n314), .C(
        \proc_in[MDATA][27] ), .D(n149), .E(dma_rp_new[11]), .F(n328), .Z(
        dma_wdata[43]) );
  HS65_LSS_XOR2X6 U427 ( .A(n62), .B(\add_545/A[11] ), .Z(dma_rp_new[11]) );
  HS65_LS_AO222X4 U428 ( .A(\add_545/A[12] ), .B(n314), .C(
        \proc_in[MDATA][28] ), .D(n149), .E(dma_rp_new[12]), .F(n328), .Z(
        dma_wdata[44]) );
  HS65_LSS_XOR2X6 U429 ( .A(n64), .B(\add_545/A[12] ), .Z(dma_rp_new[12]) );
  HS65_LS_AO222X4 U430 ( .A(\add_545/A[13] ), .B(n314), .C(
        \proc_in[MDATA][29] ), .D(n149), .E(dma_rp_new[13]), .F(n328), .Z(
        dma_wdata[45]) );
  HS65_LSS_XOR2X6 U431 ( .A(n72), .B(\add_545/A[13] ), .Z(dma_rp_new[13]) );
  HS65_LS_AO222X4 U432 ( .A(\add_545/A[14] ), .B(n313), .C(
        \proc_in[MDATA][30] ), .D(n149), .E(dma_rp_new[14]), .F(n328), .Z(
        dma_wdata[46]) );
  HS65_LSS_XOR2X6 U433 ( .A(n73), .B(\add_545/A[14] ), .Z(dma_rp_new[14]) );
  HS65_LS_AO222X4 U434 ( .A(dma_rp_new[0]), .B(n314), .C(\proc_in[MDATA][16] ), 
        .D(n144), .E(dma_rp_new[0]), .F(n327), .Z(dma_wdata[32]) );
  HS65_LS_NOR2AX3 U435 ( .A(dma_rdata[32]), .B(n85), .Z(dma_rp_new[0]) );
  HS65_LSS_XOR2X6 U436 ( .A(\add_545/A[15] ), .B(n6), .Z(dma_rp_new[15]) );
  HS65_LS_IVX9 U437 ( .A(n10), .Z(\add_545/A[15] ) );
  HS65_LH_OAI12X2 U438 ( .A(state_cnt[1]), .B(n308), .C(n312), .Z(
        phit_togo[34]) );
  HS65_LS_NAND2X7 U439 ( .A(dma_rdata[51]), .B(n138), .Z(n126) );
  HS65_LS_NAND2X7 U440 ( .A(dma_rdata[52]), .B(n138), .Z(n123) );
  HS65_LS_NAND2X7 U441 ( .A(dma_rdata[55]), .B(n139), .Z(n121) );
  HS65_LS_NAND2X7 U442 ( .A(dma_rdata[56]), .B(n138), .Z(n119) );
  HS65_LS_NAND2X7 U443 ( .A(dma_rdata[58]), .B(n138), .Z(n115) );
  HS65_LS_NAND2X7 U444 ( .A(dma_rdata[60]), .B(n138), .Z(n110) );
  HS65_LS_NAND2X7 U445 ( .A(dma_rdata[49]), .B(n139), .Z(n65) );
  HS65_LS_NAND2X7 U446 ( .A(dma_rdata[50]), .B(n139), .Z(n66) );
  HS65_LS_NAND2X7 U447 ( .A(dma_rdata[53]), .B(n138), .Z(n67) );
  HS65_LS_NAND2X7 U448 ( .A(dma_rdata[54]), .B(n138), .Z(n68) );
  HS65_LS_NAND2X7 U449 ( .A(dma_rdata[57]), .B(n139), .Z(n69) );
  HS65_LS_NAND2X7 U450 ( .A(dma_rdata[59]), .B(n138), .Z(n70) );
  HS65_LS_AOI312X4 U451 ( .A(n120), .B(n118), .C(n460), .D(n458), .E(n26), .F(
        n457), .Z(n109) );
  HS65_LS_IVX9 U452 ( .A(dma_rdata[62]), .Z(n642) );
  HS65_LH_MUX21X4 U453 ( .D0(n120), .D1(\phase_next[1] ), .S0(n645), .Z(n316)
         );
  HS65_LS_NAND3AX6 U454 ( .A(phitIn[33]), .B(phitIn[32]), .C(phitIn[34]), .Z(
        n60) );
  HS65_LS_NAND2X7 U455 ( .A(phitIn[33]), .B(phitIn[34]), .Z(n63) );
  HS65_LS_NAND3X5 U456 ( .A(n444), .B(n574), .C(n301), .Z(n358) );
  HS65_LS_NAND2X7 U457 ( .A(dma_rdata[48]), .B(n138), .Z(n131) );
  HS65_LS_NAND2X7 U458 ( .A(dma_rdata[61]), .B(n138), .Z(n107) );
  HS65_LS_BFX9 U459 ( .A(n61), .Z(n293) );
  HS65_LS_NOR3AX2 U460 ( .A(phitIn[34]), .B(phitIn[32]), .C(phitIn[33]), .Z(
        n61) );
  HS65_LS_AO22X9 U461 ( .A(n63), .B(address[0]), .C(phitIn[17]), .D(n646), .Z(
        n240) );
  HS65_LS_AO22X9 U462 ( .A(n63), .B(address[1]), .C(phitIn[18]), .D(n646), .Z(
        n242) );
  HS65_LS_AO22X9 U463 ( .A(n63), .B(address[2]), .C(phitIn[19]), .D(n646), .Z(
        n244) );
  HS65_LS_AO22X9 U464 ( .A(n63), .B(address[3]), .C(phitIn[20]), .D(n646), .Z(
        n246) );
  HS65_LS_AO22X9 U465 ( .A(n63), .B(address[4]), .C(phitIn[21]), .D(n646), .Z(
        n248) );
  HS65_LS_AO22X9 U466 ( .A(n63), .B(address[5]), .C(phitIn[22]), .D(n646), .Z(
        n250) );
  HS65_LS_AO22X9 U467 ( .A(n63), .B(address[6]), .C(phitIn[23]), .D(n646), .Z(
        n252) );
  HS65_LS_IVX9 U468 ( .A(slt_entry[2]), .Z(n644) );
  HS65_LS_IVX9 U469 ( .A(slt_entry[3]), .Z(n643) );
  HS65_LS_AO22X9 U470 ( .A(phitIn[0]), .B(n304), .C(\spm_out[MDATA][0] ), .D(
        n301), .Z(n151) );
  HS65_LS_AO22X9 U471 ( .A(phitIn[1]), .B(n310), .C(\spm_out[MDATA][1] ), .D(
        n301), .Z(n152) );
  HS65_LS_AO22X9 U472 ( .A(phitIn[2]), .B(n310), .C(\spm_out[MDATA][2] ), .D(
        n301), .Z(n153) );
  HS65_LS_AO22X9 U473 ( .A(phitIn[3]), .B(n310), .C(\spm_out[MDATA][3] ), .D(
        n301), .Z(n154) );
  HS65_LS_AO22X9 U474 ( .A(phitIn[4]), .B(n310), .C(\spm_out[MDATA][4] ), .D(
        n300), .Z(n155) );
  HS65_LS_AO22X9 U475 ( .A(phitIn[5]), .B(n310), .C(\spm_out[MDATA][5] ), .D(
        n60), .Z(n156) );
  HS65_LS_AO22X9 U476 ( .A(phitIn[6]), .B(n310), .C(\spm_out[MDATA][6] ), .D(
        n299), .Z(n157) );
  HS65_LS_AO22X9 U477 ( .A(phitIn[7]), .B(n310), .C(\spm_out[MDATA][7] ), .D(
        n60), .Z(n158) );
  HS65_LS_AO22X9 U478 ( .A(phitIn[8]), .B(n310), .C(\spm_out[MDATA][8] ), .D(
        n60), .Z(n159) );
  HS65_LS_AO22X9 U479 ( .A(phitIn[9]), .B(n310), .C(\spm_out[MDATA][9] ), .D(
        n60), .Z(n160) );
  HS65_LS_AO22X9 U480 ( .A(phitIn[10]), .B(n306), .C(\spm_out[MDATA][10] ), 
        .D(n60), .Z(n161) );
  HS65_LS_AO22X9 U481 ( .A(phitIn[11]), .B(n306), .C(\spm_out[MDATA][11] ), 
        .D(n60), .Z(n162) );
  HS65_LS_AO22X9 U482 ( .A(phitIn[12]), .B(n306), .C(\spm_out[MDATA][12] ), 
        .D(n60), .Z(n163) );
  HS65_LS_AO22X9 U483 ( .A(phitIn[13]), .B(n306), .C(\spm_out[MDATA][13] ), 
        .D(n60), .Z(n164) );
  HS65_LS_AO22X9 U484 ( .A(phitIn[14]), .B(n306), .C(\spm_out[MDATA][14] ), 
        .D(n60), .Z(n165) );
  HS65_LS_AO22X9 U485 ( .A(phitIn[15]), .B(n306), .C(\spm_out[MDATA][15] ), 
        .D(n60), .Z(n166) );
  HS65_LS_AO22X9 U486 ( .A(phitIn[16]), .B(n306), .C(\spm_out[MDATA][16] ), 
        .D(n60), .Z(n167) );
  HS65_LS_AO22X9 U487 ( .A(phitIn[17]), .B(n306), .C(\spm_out[MDATA][17] ), 
        .D(n60), .Z(n168) );
  HS65_LS_AO22X9 U488 ( .A(phitIn[18]), .B(n306), .C(\spm_out[MDATA][18] ), 
        .D(n60), .Z(n169) );
  HS65_LS_AO22X9 U489 ( .A(phitIn[19]), .B(n306), .C(\spm_out[MDATA][19] ), 
        .D(n301), .Z(n170) );
  HS65_LS_AO22X9 U490 ( .A(phitIn[20]), .B(n306), .C(\spm_out[MDATA][20] ), 
        .D(n301), .Z(n171) );
  HS65_LS_AO22X9 U491 ( .A(phitIn[21]), .B(n306), .C(\spm_out[MDATA][21] ), 
        .D(n301), .Z(n172) );
  HS65_LS_AO22X9 U492 ( .A(phitIn[22]), .B(n306), .C(\spm_out[MDATA][22] ), 
        .D(n301), .Z(n173) );
  HS65_LS_AO22X9 U493 ( .A(phitIn[23]), .B(n306), .C(\spm_out[MDATA][23] ), 
        .D(n301), .Z(n174) );
  HS65_LS_AO22X9 U494 ( .A(phitIn[24]), .B(n306), .C(\spm_out[MDATA][24] ), 
        .D(n301), .Z(n175) );
  HS65_LS_AO22X9 U495 ( .A(phitIn[25]), .B(n306), .C(\spm_out[MDATA][25] ), 
        .D(n301), .Z(n176) );
  HS65_LS_AO22X9 U496 ( .A(phitIn[26]), .B(n306), .C(\spm_out[MDATA][26] ), 
        .D(n301), .Z(n177) );
  HS65_LS_AO22X9 U497 ( .A(phitIn[27]), .B(n306), .C(\spm_out[MDATA][27] ), 
        .D(n301), .Z(n178) );
  HS65_LS_AO22X9 U498 ( .A(phitIn[28]), .B(n306), .C(\spm_out[MDATA][28] ), 
        .D(n301), .Z(n179) );
  HS65_LS_AO22X9 U499 ( .A(phitIn[29]), .B(n306), .C(\spm_out[MDATA][29] ), 
        .D(n301), .Z(n180) );
  HS65_LS_AO22X9 U500 ( .A(phitIn[30]), .B(n305), .C(\spm_out[MDATA][30] ), 
        .D(n301), .Z(n181) );
  HS65_LS_AO22X9 U501 ( .A(phitIn[31]), .B(n305), .C(\spm_out[MDATA][31] ), 
        .D(n301), .Z(n182) );
  HS65_LS_AO22X9 U502 ( .A(dIn_h[0]), .B(n305), .C(\spm_out[MDATA][32] ), .D(
        n300), .Z(n183) );
  HS65_LS_AO22X9 U503 ( .A(dIn_h[1]), .B(n305), .C(\spm_out[MDATA][33] ), .D(
        n300), .Z(n184) );
  HS65_LS_AO22X9 U504 ( .A(dIn_h[2]), .B(n305), .C(\spm_out[MDATA][34] ), .D(
        n300), .Z(n185) );
  HS65_LS_AO22X9 U505 ( .A(dIn_h[3]), .B(n305), .C(\spm_out[MDATA][35] ), .D(
        n300), .Z(n186) );
  HS65_LS_AO22X9 U506 ( .A(dIn_h[4]), .B(n305), .C(\spm_out[MDATA][36] ), .D(
        n300), .Z(n187) );
  HS65_LS_AO22X9 U507 ( .A(dIn_h[5]), .B(n305), .C(\spm_out[MDATA][37] ), .D(
        n300), .Z(n188) );
  HS65_LS_AO22X9 U508 ( .A(dIn_h[6]), .B(n305), .C(\spm_out[MDATA][38] ), .D(
        n300), .Z(n189) );
  HS65_LS_AO22X9 U509 ( .A(dIn_h[7]), .B(n305), .C(\spm_out[MDATA][39] ), .D(
        n300), .Z(n190) );
  HS65_LS_AO22X9 U510 ( .A(dIn_h[8]), .B(n305), .C(\spm_out[MDATA][40] ), .D(
        n300), .Z(n191) );
  HS65_LS_AO22X9 U511 ( .A(dIn_h[9]), .B(n305), .C(\spm_out[MDATA][41] ), .D(
        n300), .Z(n192) );
  HS65_LS_AO22X9 U512 ( .A(dIn_h[10]), .B(n305), .C(\spm_out[MDATA][42] ), .D(
        n300), .Z(n193) );
  HS65_LS_AO22X9 U513 ( .A(dIn_h[11]), .B(n305), .C(\spm_out[MDATA][43] ), .D(
        n300), .Z(n194) );
  HS65_LS_AO22X9 U514 ( .A(dIn_h[12]), .B(n305), .C(\spm_out[MDATA][44] ), .D(
        n299), .Z(n195) );
  HS65_LS_AO22X9 U515 ( .A(dIn_h[13]), .B(n305), .C(\spm_out[MDATA][45] ), .D(
        n299), .Z(n196) );
  HS65_LS_AO22X9 U516 ( .A(dIn_h[14]), .B(n305), .C(\spm_out[MDATA][46] ), .D(
        n299), .Z(n197) );
  HS65_LS_AO22X9 U517 ( .A(dIn_h[15]), .B(n305), .C(\spm_out[MDATA][47] ), .D(
        n299), .Z(n198) );
  HS65_LS_AO22X9 U518 ( .A(dIn_h[16]), .B(n305), .C(\spm_out[MDATA][48] ), .D(
        n299), .Z(n199) );
  HS65_LS_AO22X9 U519 ( .A(dIn_h[17]), .B(n304), .C(\spm_out[MDATA][49] ), .D(
        n299), .Z(n200) );
  HS65_LS_AO22X9 U520 ( .A(dIn_h[18]), .B(n304), .C(\spm_out[MDATA][50] ), .D(
        n299), .Z(n201) );
  HS65_LS_AO22X9 U521 ( .A(dIn_h[19]), .B(n304), .C(\spm_out[MDATA][51] ), .D(
        n299), .Z(n202) );
  HS65_LS_AO22X9 U522 ( .A(dIn_h[20]), .B(n305), .C(\spm_out[MDATA][52] ), .D(
        n299), .Z(n203) );
  HS65_LS_AO22X9 U523 ( .A(dIn_h[21]), .B(n304), .C(\spm_out[MDATA][53] ), .D(
        n300), .Z(n204) );
  HS65_LS_AO22X9 U524 ( .A(dIn_h[22]), .B(n304), .C(\spm_out[MDATA][54] ), .D(
        n299), .Z(n205) );
  HS65_LS_AO22X9 U525 ( .A(dIn_h[23]), .B(n304), .C(\spm_out[MDATA][55] ), .D(
        n299), .Z(n206) );
  HS65_LS_AO22X9 U526 ( .A(dIn_h[24]), .B(n304), .C(\spm_out[MDATA][56] ), .D(
        n299), .Z(n207) );
  HS65_LS_AO22X9 U527 ( .A(dIn_h[25]), .B(n304), .C(\spm_out[MDATA][57] ), .D(
        n299), .Z(n208) );
  HS65_LS_AO22X9 U528 ( .A(dIn_h[26]), .B(n304), .C(\spm_out[MDATA][58] ), .D(
        n299), .Z(n209) );
  HS65_LS_AO22X9 U529 ( .A(dIn_h[27]), .B(n304), .C(\spm_out[MDATA][59] ), .D(
        n300), .Z(n210) );
  HS65_LS_AO22X9 U530 ( .A(dIn_h[28]), .B(n304), .C(\spm_out[MDATA][60] ), .D(
        n299), .Z(n211) );
  HS65_LS_AO22X9 U531 ( .A(dIn_h[29]), .B(n304), .C(\spm_out[MDATA][61] ), .D(
        n300), .Z(n212) );
  HS65_LS_AO22X9 U532 ( .A(dIn_h[30]), .B(n304), .C(\spm_out[MDATA][62] ), .D(
        n299), .Z(n213) );
  HS65_LS_AO22X9 U533 ( .A(dIn_h[31]), .B(n304), .C(\spm_out[MDATA][63] ), .D(
        n301), .Z(n214) );
  HS65_LS_AO22X9 U534 ( .A(phitIn[17]), .B(n297), .C(n295), .D(dIn_h[17]), .Z(
        n239) );
  HS65_LS_AO22X9 U535 ( .A(phitIn[18]), .B(n297), .C(n295), .D(dIn_h[18]), .Z(
        n241) );
  HS65_LS_AO22X9 U536 ( .A(phitIn[19]), .B(n297), .C(n295), .D(dIn_h[19]), .Z(
        n243) );
  HS65_LS_AO22X9 U537 ( .A(phitIn[20]), .B(n297), .C(n295), .D(dIn_h[20]), .Z(
        n245) );
  HS65_LS_AO22X9 U538 ( .A(phitIn[21]), .B(n298), .C(n295), .D(dIn_h[21]), .Z(
        n247) );
  HS65_LS_AO22X9 U539 ( .A(phitIn[22]), .B(n298), .C(n295), .D(dIn_h[22]), .Z(
        n249) );
  HS65_LS_AO22X9 U540 ( .A(phitIn[23]), .B(n298), .C(n295), .D(dIn_h[23]), .Z(
        n251) );
  HS65_LS_AO22X9 U541 ( .A(phitIn[0]), .B(n296), .C(n294), .D(dIn_h[0]), .Z(
        n222) );
  HS65_LS_AO22X9 U542 ( .A(phitIn[1]), .B(n297), .C(n294), .D(dIn_h[1]), .Z(
        n223) );
  HS65_LS_AO22X9 U543 ( .A(phitIn[2]), .B(n297), .C(n294), .D(dIn_h[2]), .Z(
        n224) );
  HS65_LS_AO22X9 U544 ( .A(phitIn[3]), .B(n297), .C(n294), .D(dIn_h[3]), .Z(
        n225) );
  HS65_LS_AO22X9 U545 ( .A(phitIn[4]), .B(n297), .C(n294), .D(dIn_h[4]), .Z(
        n226) );
  HS65_LS_AO22X9 U546 ( .A(phitIn[5]), .B(n297), .C(n294), .D(dIn_h[5]), .Z(
        n227) );
  HS65_LS_AO22X9 U547 ( .A(phitIn[6]), .B(n297), .C(n294), .D(dIn_h[6]), .Z(
        n228) );
  HS65_LS_AO22X9 U548 ( .A(phitIn[7]), .B(n297), .C(n294), .D(dIn_h[7]), .Z(
        n229) );
  HS65_LS_AO22X9 U549 ( .A(phitIn[8]), .B(n297), .C(n294), .D(dIn_h[8]), .Z(
        n230) );
  HS65_LS_AO22X9 U550 ( .A(phitIn[9]), .B(n297), .C(n294), .D(dIn_h[9]), .Z(
        n231) );
  HS65_LS_AO22X9 U551 ( .A(phitIn[10]), .B(n297), .C(n294), .D(dIn_h[10]), .Z(
        n232) );
  HS65_LS_AO22X9 U552 ( .A(phitIn[11]), .B(n297), .C(n294), .D(dIn_h[11]), .Z(
        n233) );
  HS65_LS_AO22X9 U553 ( .A(phitIn[12]), .B(n297), .C(n294), .D(dIn_h[12]), .Z(
        n234) );
  HS65_LS_AO22X9 U554 ( .A(phitIn[13]), .B(n297), .C(n295), .D(dIn_h[13]), .Z(
        n235) );
  HS65_LS_AO22X9 U555 ( .A(phitIn[14]), .B(n297), .C(n295), .D(dIn_h[14]), .Z(
        n236) );
  HS65_LS_AO22X9 U556 ( .A(phitIn[15]), .B(n297), .C(n295), .D(dIn_h[15]), .Z(
        n237) );
  HS65_LS_AO22X9 U557 ( .A(phitIn[16]), .B(n297), .C(n295), .D(dIn_h[16]), .Z(
        n238) );
  HS65_LS_AO22X9 U558 ( .A(phitIn[24]), .B(n298), .C(n295), .D(dIn_h[24]), .Z(
        n253) );
  HS65_LS_AO22X9 U559 ( .A(phitIn[25]), .B(n298), .C(n295), .D(dIn_h[25]), .Z(
        n254) );
  HS65_LS_AO22X9 U560 ( .A(phitIn[26]), .B(n298), .C(n294), .D(dIn_h[26]), .Z(
        n255) );
  HS65_LS_AO22X9 U561 ( .A(phitIn[27]), .B(n298), .C(n295), .D(dIn_h[27]), .Z(
        n256) );
  HS65_LS_AO22X9 U562 ( .A(phitIn[28]), .B(n298), .C(n294), .D(dIn_h[28]), .Z(
        n257) );
  HS65_LS_AO22X9 U563 ( .A(phitIn[29]), .B(n298), .C(n295), .D(dIn_h[29]), .Z(
        n258) );
  HS65_LS_AO22X9 U564 ( .A(phitIn[30]), .B(n298), .C(n294), .D(dIn_h[30]), .Z(
        n259) );
  HS65_LS_AO22X9 U565 ( .A(phitIn[31]), .B(n298), .C(n295), .D(dIn_h[31]), .Z(
        n260) );
  HS65_LS_AO22X9 U566 ( .A(n304), .B(address[0]), .C(n300), .D(flit_buf[64]), 
        .Z(n215) );
  HS65_LS_AO22X9 U567 ( .A(n304), .B(address[1]), .C(n299), .D(flit_buf[65]), 
        .Z(n216) );
  HS65_LS_AO22X9 U568 ( .A(n304), .B(address[2]), .C(n300), .D(flit_buf[66]), 
        .Z(n217) );
  HS65_LS_AO22X9 U569 ( .A(n304), .B(address[3]), .C(n299), .D(flit_buf[67]), 
        .Z(n218) );
  HS65_LS_AO22X9 U570 ( .A(n303), .B(address[4]), .C(n300), .D(flit_buf[68]), 
        .Z(n219) );
  HS65_LS_AO22X9 U571 ( .A(n302), .B(address[5]), .C(n299), .D(flit_buf[69]), 
        .Z(n220) );
  HS65_LS_AO22X9 U572 ( .A(n304), .B(address[6]), .C(n300), .D(flit_buf[70]), 
        .Z(n221) );
  HS65_LS_OR2X9 U573 ( .A(vld_pkt), .B(n646), .Z(n318) );
  HS65_LS_NAND2X7 U574 ( .A(\proc_in[MADDR][0] ), .B(n146), .Z(n71) );
  HS65_LS_NOR4ABX2 U575 ( .A(n653), .B(n150), .C(\proc_in[MADDR][26] ), .D(
        \proc_in[MADDR][24] ), .Z(n76) );
  HS65_LS_IVX9 U576 ( .A(\proc_in[MADDR][25] ), .Z(n653) );
  HS65_LS_NOR3X4 U577 ( .A(\proc_in[MADDR][27] ), .B(\proc_in[MADDR][31] ), 
        .C(\proc_in[MADDR][30] ), .Z(n150) );
  HS65_LS_NAND4ABX3 U578 ( .A(\proc_in[MADDR][29] ), .B(\proc_in[MADDR][26] ), 
        .C(n147), .D(n148), .Z(n82) );
  HS65_LS_NOR2X6 U579 ( .A(\proc_in[MADDR][31] ), .B(\proc_in[MADDR][30] ), 
        .Z(n147) );
  HS65_LS_NOR4ABX2 U580 ( .A(\proc_in[MADDR][28] ), .B(\proc_in[MADDR][27] ), 
        .C(\proc_in[MADDR][25] ), .D(\proc_in[MADDR][24] ), .Z(n148) );
  HS65_LS_NOR3AX2 U581 ( .A(n76), .B(n652), .C(\proc_in[MADDR][29] ), .Z(n322)
         );
  HS65_LS_NAND4ABX3 U582 ( .A(config_reg[3]), .B(n33), .C(config_reg[4]), .D(
        n590), .Z(n16) );
  HS65_LS_OA32X4 U583 ( .A(config_reg[0]), .B(config_reg[1]), .C(n647), .D(n36), .E(config_reg[2]), .Z(n33) );
  HS65_LS_IVX9 U584 ( .A(config_reg[2]), .Z(n647) );
  HS65_LSS_XNOR2X6 U585 ( .A(config_reg[1]), .B(config_reg[0]), .Z(n36) );
  HS65_LS_BFX9 U586 ( .A(na_reset), .Z(n335) );
  HS65_LS_BFX9 U587 ( .A(na_reset), .Z(n334) );
  HS65_LS_NAND2X7 U588 ( .A(n322), .B(\proc_in[MCMD][0] ), .Z(n38) );
  HS65_LS_IVX9 U589 ( .A(\proc_in[MDATA][15] ), .Z(n657) );
  HS65_LS_IVX9 U590 ( .A(\proc_in[MDATA][6] ), .Z(n666) );
  HS65_LS_IVX9 U591 ( .A(\proc_in[MDATA][7] ), .Z(n665) );
  HS65_LS_IVX9 U592 ( .A(\proc_in[MDATA][8] ), .Z(n664) );
  HS65_LS_IVX9 U593 ( .A(\proc_in[MDATA][9] ), .Z(n663) );
  HS65_LS_IVX9 U594 ( .A(\proc_in[MADDR][28] ), .Z(n652) );
  HS65_LS_AND3X9 U595 ( .A(n76), .B(n652), .C(\proc_in[MADDR][29] ), .Z(n146)
         );
  HS65_LS_IVX9 U596 ( .A(\proc_in[MDATA][14] ), .Z(n658) );
  HS65_LS_IVX9 U597 ( .A(\proc_in[MDATA][0] ), .Z(n672) );
  HS65_LS_IVX9 U598 ( .A(\proc_in[MDATA][1] ), .Z(n671) );
  HS65_LS_IVX9 U599 ( .A(\proc_in[MDATA][2] ), .Z(n670) );
  HS65_LS_IVX9 U600 ( .A(\proc_in[MDATA][3] ), .Z(n669) );
  HS65_LS_IVX9 U601 ( .A(\proc_in[MDATA][4] ), .Z(n668) );
  HS65_LS_IVX9 U602 ( .A(\proc_in[MDATA][5] ), .Z(n667) );
  HS65_LS_IVX9 U603 ( .A(\proc_in[MDATA][10] ), .Z(n662) );
  HS65_LS_IVX9 U604 ( .A(\proc_in[MDATA][11] ), .Z(n661) );
  HS65_LS_IVX9 U605 ( .A(\proc_in[MDATA][12] ), .Z(n660) );
  HS65_LS_IVX9 U606 ( .A(\proc_in[MDATA][13] ), .Z(n659) );
  HS65_LS_IVX9 U607 ( .A(\proc_in[MADDR][0] ), .Z(n656) );
  HS65_LS_IVX9 U608 ( .A(\proc_in[MADDR][1] ), .Z(n655) );
  HS65_LH_NAND2X2 U609 ( .A(n26), .B(n447), .Z(n360) );
  HS65_LH_AND2X4 U610 ( .A(n26), .B(n410), .Z(phit_togo[32]) );
  HS65_LS_AND2X18 U611 ( .A(n443), .B(n447), .Z(n118) );
  HS65_LS_IVX7 U612 ( .A(n456), .Z(n457) );
  HS65_LH_BFX2 U613 ( .A(n2), .Z(n132) );
  HS65_LS_BFX9 U614 ( .A(n132), .Z(n134) );
  HS65_LS_BFX9 U615 ( .A(n132), .Z(n133) );
  HS65_LS_BFX9 U616 ( .A(n132), .Z(n136) );
  HS65_LH_NAND2X2 U617 ( .A(n443), .B(n447), .Z(n444) );
  HS65_LH_CBI4I1X5 U618 ( .A(n444), .B(n359), .C(n301), .D(n358), .Z(n317) );
  HS65_LS_IVX18 U619 ( .A(\phase_prev[0] ), .Z(n448) );
  HS65_LS_NAND2X7 U620 ( .A(dma_rdata[39]), .B(n139), .Z(n588) );
  HS65_LS_IVX9 U621 ( .A(n588), .Z(n617) );
  HS65_LS_NAND2X7 U622 ( .A(dma_rdata[38]), .B(n138), .Z(n586) );
  HS65_LS_IVX9 U623 ( .A(n586), .Z(n616) );
  HS65_LS_NAND2X7 U624 ( .A(dma_rdata[37]), .B(n138), .Z(n584) );
  HS65_LS_IVX9 U625 ( .A(n584), .Z(n615) );
  HS65_LS_NAND2X7 U626 ( .A(dma_rdata[36]), .B(n138), .Z(n582) );
  HS65_LS_IVX9 U627 ( .A(n582), .Z(n614) );
  HS65_LS_NAND2X7 U628 ( .A(dma_rdata[35]), .B(n618), .Z(n580) );
  HS65_LS_IVX9 U629 ( .A(n580), .Z(n613) );
  HS65_LS_NAND2X7 U630 ( .A(dma_rdata[34]), .B(n618), .Z(n578) );
  HS65_LS_IVX9 U631 ( .A(n578), .Z(n612) );
  HS65_LS_NAND2X7 U632 ( .A(dma_rdata[33]), .B(n618), .Z(n576) );
  HS65_LS_IVX9 U633 ( .A(n576), .Z(n611) );
  HS65_LS_NAND2X7 U634 ( .A(dma_rdata[31]), .B(n139), .Z(n408) );
  HS65_LS_IVX9 U635 ( .A(n408), .Z(n610) );
  HS65_LS_NAND2X7 U636 ( .A(dma_rdata[30]), .B(n138), .Z(n406) );
  HS65_LS_IVX9 U637 ( .A(n406), .Z(n609) );
  HS65_LS_NAND2X7 U638 ( .A(dma_rdata[29]), .B(n139), .Z(n404) );
  HS65_LS_IVX9 U639 ( .A(n404), .Z(n608) );
  HS65_LS_NAND2X7 U640 ( .A(dma_rdata[28]), .B(n139), .Z(n402) );
  HS65_LS_IVX9 U641 ( .A(n402), .Z(n607) );
  HS65_LS_NAND2X7 U642 ( .A(dma_rdata[27]), .B(n138), .Z(n400) );
  HS65_LS_IVX9 U643 ( .A(n400), .Z(n606) );
  HS65_LS_NAND2X7 U644 ( .A(dma_rdata[26]), .B(n139), .Z(n398) );
  HS65_LS_IVX9 U645 ( .A(n398), .Z(n605) );
  HS65_LS_NAND2X7 U646 ( .A(dma_rdata[25]), .B(n138), .Z(n396) );
  HS65_LS_IVX9 U647 ( .A(n396), .Z(n604) );
  HS65_LS_NAND2X7 U648 ( .A(dma_rdata[24]), .B(n138), .Z(n394) );
  HS65_LS_IVX9 U649 ( .A(n394), .Z(n603) );
  HS65_LS_NAND2X7 U650 ( .A(dma_rdata[23]), .B(n139), .Z(n392) );
  HS65_LS_IVX9 U651 ( .A(n392), .Z(n602) );
  HS65_LS_NAND2X7 U652 ( .A(dma_rdata[22]), .B(n139), .Z(n390) );
  HS65_LS_IVX9 U653 ( .A(n390), .Z(n601) );
  HS65_LS_NAND2X7 U654 ( .A(dma_rdata[21]), .B(n138), .Z(n388) );
  HS65_LS_IVX9 U655 ( .A(n388), .Z(n600) );
  HS65_LS_NAND2X7 U656 ( .A(dma_rdata[20]), .B(n139), .Z(n386) );
  HS65_LS_IVX9 U657 ( .A(n386), .Z(n599) );
  HS65_LS_NAND2X7 U658 ( .A(dma_rdata[19]), .B(n618), .Z(n384) );
  HS65_LS_IVX9 U659 ( .A(n384), .Z(n598) );
  HS65_LS_NAND2X7 U660 ( .A(dma_rdata[18]), .B(n618), .Z(n382) );
  HS65_LS_IVX9 U661 ( .A(n382), .Z(n597) );
  HS65_LS_NAND2X7 U662 ( .A(dma_rdata[17]), .B(n618), .Z(n380) );
  HS65_LS_IVX9 U663 ( .A(n380), .Z(n596) );
  HS65_LS_IVX9 U664 ( .A(\proc_in[MCMD][0] ), .Z(n355) );
  HS65_LS_IVX9 U665 ( .A(n357), .Z(n356) );
  HS65_LS_NAND2X7 U666 ( .A(n141), .B(n4), .Z(n83) );
  HS65_LS_OAI22X6 U667 ( .A(n643), .B(n360), .C(n143), .D(n357), .Z(
        dma_raddr[1]) );
  HS65_LS_OAI22X6 U668 ( .A(n644), .B(n360), .C(n145), .D(n357), .Z(
        dma_raddr[0]) );
  HS65_LS_NAND2X7 U669 ( .A(dma_rdata[16]), .B(n139), .Z(n378) );
  HS65_LS_IVX9 U670 ( .A(n378), .Z(n593) );
  HS65_LS_IVX9 U671 ( .A(n307), .Z(n449) );
  HS65_LS_IVX9 U672 ( .A(vld_pkt), .Z(n359) );
  HS65_LS_IVX9 U673 ( .A(n309), .Z(n574) );
  HS65_LS_IVX9 U674 ( .A(n360), .Z(n595) );
  HS65_LS_IVX9 U675 ( .A(n308), .Z(n410) );
  HS65_LS_NAND2X7 U676 ( .A(n595), .B(n410), .Z(n409) );
  HS65_LS_IVX9 U677 ( .A(dOut_l[0]), .Z(n411) );
  HS65_LS_NAND2X7 U678 ( .A(\spm_in[SDATA][32] ), .B(n122), .Z(n361) );
  HS65_LS_OAI212X5 U679 ( .A(n128), .B(n411), .C(n324), .D(n640), .E(n361), 
        .Z(mux_out[0]) );
  HS65_LS_IVX9 U680 ( .A(dOut_l[1]), .Z(n412) );
  HS65_LS_NAND2X7 U681 ( .A(\spm_in[SDATA][33] ), .B(n122), .Z(n362) );
  HS65_LS_OAI212X5 U682 ( .A(n128), .B(n412), .C(n324), .D(n639), .E(n362), 
        .Z(mux_out[1]) );
  HS65_LS_IVX9 U683 ( .A(dOut_l[2]), .Z(n413) );
  HS65_LS_NAND2X7 U684 ( .A(\spm_in[SDATA][34] ), .B(n122), .Z(n363) );
  HS65_LS_OAI212X5 U685 ( .A(n128), .B(n413), .C(n324), .D(n638), .E(n363), 
        .Z(mux_out[2]) );
  HS65_LS_IVX9 U686 ( .A(dOut_l[3]), .Z(n414) );
  HS65_LS_NAND2X7 U687 ( .A(\spm_in[SDATA][35] ), .B(n122), .Z(n364) );
  HS65_LS_OAI212X5 U688 ( .A(n128), .B(n414), .C(n324), .D(n637), .E(n364), 
        .Z(mux_out[3]) );
  HS65_LS_IVX9 U689 ( .A(dOut_l[4]), .Z(n415) );
  HS65_LS_NAND2X7 U690 ( .A(\spm_in[SDATA][36] ), .B(n122), .Z(n365) );
  HS65_LS_OAI212X5 U691 ( .A(n128), .B(n415), .C(n324), .D(n636), .E(n365), 
        .Z(mux_out[4]) );
  HS65_LS_IVX9 U692 ( .A(dOut_l[5]), .Z(n416) );
  HS65_LS_NAND2X7 U693 ( .A(\spm_in[SDATA][37] ), .B(n122), .Z(n366) );
  HS65_LS_OAI212X5 U694 ( .A(n128), .B(n416), .C(n324), .D(n635), .E(n366), 
        .Z(mux_out[5]) );
  HS65_LS_IVX9 U695 ( .A(dOut_l[6]), .Z(n417) );
  HS65_LS_NAND2X7 U696 ( .A(\spm_in[SDATA][38] ), .B(n122), .Z(n367) );
  HS65_LS_OAI212X5 U697 ( .A(n128), .B(n417), .C(n324), .D(n634), .E(n367), 
        .Z(mux_out[6]) );
  HS65_LS_IVX9 U698 ( .A(dOut_l[7]), .Z(n418) );
  HS65_LS_NAND2X7 U699 ( .A(\spm_in[SDATA][39] ), .B(n122), .Z(n368) );
  HS65_LS_OAI212X5 U700 ( .A(n128), .B(n418), .C(n324), .D(n633), .E(n368), 
        .Z(mux_out[7]) );
  HS65_LS_IVX9 U701 ( .A(dOut_l[8]), .Z(n419) );
  HS65_LS_NAND2X7 U702 ( .A(\spm_in[SDATA][40] ), .B(n122), .Z(n369) );
  HS65_LS_OAI212X5 U703 ( .A(n128), .B(n419), .C(n324), .D(n632), .E(n369), 
        .Z(mux_out[8]) );
  HS65_LS_IVX9 U704 ( .A(dOut_l[9]), .Z(n420) );
  HS65_LS_NAND2X7 U705 ( .A(\spm_in[SDATA][41] ), .B(n122), .Z(n370) );
  HS65_LS_OAI212X5 U706 ( .A(n128), .B(n420), .C(n323), .D(n631), .E(n370), 
        .Z(mux_out[9]) );
  HS65_LS_IVX9 U707 ( .A(dOut_l[10]), .Z(n421) );
  HS65_LS_NAND2X7 U708 ( .A(\spm_in[SDATA][42] ), .B(n122), .Z(n371) );
  HS65_LS_OAI212X5 U709 ( .A(n128), .B(n421), .C(n323), .D(n630), .E(n371), 
        .Z(mux_out[10]) );
  HS65_LS_IVX9 U710 ( .A(dOut_l[11]), .Z(n422) );
  HS65_LS_NAND2X7 U711 ( .A(\spm_in[SDATA][43] ), .B(n122), .Z(n372) );
  HS65_LS_OAI212X5 U712 ( .A(n128), .B(n422), .C(n323), .D(n629), .E(n372), 
        .Z(mux_out[11]) );
  HS65_LS_IVX9 U713 ( .A(dOut_l[12]), .Z(n423) );
  HS65_LS_NAND2X7 U714 ( .A(\spm_in[SDATA][44] ), .B(n124), .Z(n373) );
  HS65_LS_OAI212X5 U715 ( .A(n129), .B(n423), .C(n323), .D(n628), .E(n373), 
        .Z(mux_out[12]) );
  HS65_LS_IVX9 U716 ( .A(dOut_l[13]), .Z(n424) );
  HS65_LS_NAND2X7 U717 ( .A(\spm_in[SDATA][45] ), .B(n124), .Z(n374) );
  HS65_LS_OAI212X5 U718 ( .A(n129), .B(n424), .C(n323), .D(n627), .E(n374), 
        .Z(mux_out[13]) );
  HS65_LS_IVX9 U719 ( .A(dOut_l[14]), .Z(n425) );
  HS65_LS_NAND2X7 U720 ( .A(\spm_in[SDATA][46] ), .B(n124), .Z(n375) );
  HS65_LS_OAI212X5 U721 ( .A(n129), .B(n425), .C(n323), .D(n626), .E(n375), 
        .Z(mux_out[14]) );
  HS65_LS_IVX9 U722 ( .A(dOut_l[15]), .Z(n426) );
  HS65_LS_NAND2X7 U723 ( .A(\spm_in[SDATA][47] ), .B(n124), .Z(n376) );
  HS65_LS_OAI212X5 U724 ( .A(n129), .B(n426), .C(n323), .D(n625), .E(n376), 
        .Z(mux_out[15]) );
  HS65_LS_IVX9 U725 ( .A(dOut_l[16]), .Z(n427) );
  HS65_LS_NAND2X7 U726 ( .A(\spm_in[SDATA][48] ), .B(n124), .Z(n377) );
  HS65_LS_OAI212X5 U727 ( .A(n129), .B(n427), .C(n323), .D(n378), .E(n377), 
        .Z(mux_out[16]) );
  HS65_LS_IVX9 U728 ( .A(dOut_l[17]), .Z(n428) );
  HS65_LS_NAND2X7 U729 ( .A(\spm_in[SDATA][49] ), .B(n124), .Z(n379) );
  HS65_LS_IVX9 U730 ( .A(dOut_l[18]), .Z(n429) );
  HS65_LS_NAND2X7 U731 ( .A(\spm_in[SDATA][50] ), .B(n124), .Z(n381) );
  HS65_LS_IVX9 U732 ( .A(dOut_l[19]), .Z(n430) );
  HS65_LS_NAND2X7 U733 ( .A(\spm_in[SDATA][51] ), .B(n124), .Z(n383) );
  HS65_LS_OAI212X5 U734 ( .A(n129), .B(n430), .C(n323), .D(n384), .E(n383), 
        .Z(mux_out[19]) );
  HS65_LS_IVX9 U735 ( .A(dOut_l[20]), .Z(n431) );
  HS65_LS_NAND2X7 U736 ( .A(\spm_in[SDATA][52] ), .B(n124), .Z(n385) );
  HS65_LS_OAI212X5 U737 ( .A(n129), .B(n431), .C(n323), .D(n386), .E(n385), 
        .Z(mux_out[20]) );
  HS65_LS_IVX9 U738 ( .A(dOut_l[21]), .Z(n432) );
  HS65_LS_NAND2X7 U739 ( .A(\spm_in[SDATA][53] ), .B(n124), .Z(n387) );
  HS65_LS_OAI212X5 U740 ( .A(n129), .B(n432), .C(n323), .D(n388), .E(n387), 
        .Z(mux_out[21]) );
  HS65_LS_IVX9 U741 ( .A(dOut_l[22]), .Z(n433) );
  HS65_LS_NAND2X7 U742 ( .A(\spm_in[SDATA][54] ), .B(n124), .Z(n389) );
  HS65_LS_OAI212X5 U743 ( .A(n129), .B(n433), .C(n323), .D(n390), .E(n389), 
        .Z(mux_out[22]) );
  HS65_LS_IVX9 U744 ( .A(dOut_l[23]), .Z(n434) );
  HS65_LS_NAND2X7 U745 ( .A(\spm_in[SDATA][55] ), .B(n124), .Z(n391) );
  HS65_LS_OAI212X5 U746 ( .A(n129), .B(n434), .C(n323), .D(n392), .E(n391), 
        .Z(mux_out[23]) );
  HS65_LS_IVX9 U747 ( .A(dOut_l[24]), .Z(n435) );
  HS65_LS_NAND2X7 U748 ( .A(\spm_in[SDATA][56] ), .B(n125), .Z(n393) );
  HS65_LS_OAI212X5 U749 ( .A(n130), .B(n435), .C(n323), .D(n394), .E(n393), 
        .Z(mux_out[24]) );
  HS65_LS_IVX9 U750 ( .A(dOut_l[25]), .Z(n436) );
  HS65_LS_NAND2X7 U751 ( .A(\spm_in[SDATA][57] ), .B(n125), .Z(n395) );
  HS65_LS_OAI212X5 U752 ( .A(n130), .B(n436), .C(n323), .D(n396), .E(n395), 
        .Z(mux_out[25]) );
  HS65_LS_IVX9 U753 ( .A(dOut_l[26]), .Z(n437) );
  HS65_LS_NAND2X7 U754 ( .A(\spm_in[SDATA][58] ), .B(n125), .Z(n397) );
  HS65_LS_OAI212X5 U755 ( .A(n130), .B(n437), .C(n323), .D(n398), .E(n397), 
        .Z(mux_out[26]) );
  HS65_LS_IVX9 U756 ( .A(dOut_l[27]), .Z(n438) );
  HS65_LS_NAND2X7 U757 ( .A(\spm_in[SDATA][59] ), .B(n125), .Z(n399) );
  HS65_LS_OAI212X5 U758 ( .A(n130), .B(n438), .C(n314), .D(n400), .E(n399), 
        .Z(mux_out[27]) );
  HS65_LS_IVX9 U759 ( .A(dOut_l[28]), .Z(n439) );
  HS65_LS_NAND2X7 U760 ( .A(\spm_in[SDATA][60] ), .B(n125), .Z(n401) );
  HS65_LS_OAI212X5 U761 ( .A(n130), .B(n439), .C(n323), .D(n402), .E(n401), 
        .Z(mux_out[28]) );
  HS65_LS_IVX9 U762 ( .A(dOut_l[29]), .Z(n440) );
  HS65_LS_NAND2X7 U763 ( .A(\spm_in[SDATA][61] ), .B(n125), .Z(n403) );
  HS65_LS_OAI212X5 U764 ( .A(n130), .B(n440), .C(n314), .D(n404), .E(n403), 
        .Z(mux_out[29]) );
  HS65_LS_IVX9 U765 ( .A(dOut_l[30]), .Z(n441) );
  HS65_LS_NAND2X7 U766 ( .A(\spm_in[SDATA][62] ), .B(n125), .Z(n405) );
  HS65_LS_OAI212X5 U767 ( .A(n130), .B(n441), .C(n323), .D(n406), .E(n405), 
        .Z(mux_out[30]) );
  HS65_LS_IVX9 U768 ( .A(dOut_l[31]), .Z(n442) );
  HS65_LS_NAND2X7 U769 ( .A(\spm_in[SDATA][63] ), .B(n125), .Z(n407) );
  HS65_LS_OAI212X5 U770 ( .A(n130), .B(n442), .C(n314), .D(n408), .E(n407), 
        .Z(mux_out[31]) );
  HS65_LS_MUX21I1X6 U771 ( .D0(n411), .D1(\spm_in[SDATA][0] ), .S0(n134), .Z(
        n261) );
  HS65_LS_MUX21I1X6 U772 ( .D0(n412), .D1(\spm_in[SDATA][1] ), .S0(n134), .Z(
        n262) );
  HS65_LS_MUX21I1X6 U773 ( .D0(n413), .D1(\spm_in[SDATA][2] ), .S0(n133), .Z(
        n263) );
  HS65_LS_MUX21I1X6 U774 ( .D0(n414), .D1(\spm_in[SDATA][3] ), .S0(n136), .Z(
        n264) );
  HS65_LS_MUX21I1X6 U775 ( .D0(n415), .D1(\spm_in[SDATA][4] ), .S0(n133), .Z(
        n265) );
  HS65_LS_MUX21I1X6 U776 ( .D0(n416), .D1(\spm_in[SDATA][5] ), .S0(n136), .Z(
        n266) );
  HS65_LS_MUX21I1X6 U777 ( .D0(n417), .D1(\spm_in[SDATA][6] ), .S0(n134), .Z(
        n267) );
  HS65_LS_MUX21I1X6 U778 ( .D0(n418), .D1(\spm_in[SDATA][7] ), .S0(n133), .Z(
        n268) );
  HS65_LS_MUX21I1X6 U779 ( .D0(n419), .D1(\spm_in[SDATA][8] ), .S0(n136), .Z(
        n269) );
  HS65_LS_MUX21I1X6 U780 ( .D0(n420), .D1(\spm_in[SDATA][9] ), .S0(n134), .Z(
        n270) );
  HS65_LS_MUX21I1X6 U781 ( .D0(n421), .D1(\spm_in[SDATA][10] ), .S0(n133), .Z(
        n271) );
  HS65_LS_MUX21I1X6 U782 ( .D0(n422), .D1(\spm_in[SDATA][11] ), .S0(n136), .Z(
        n272) );
  HS65_LS_MUX21I1X6 U783 ( .D0(n423), .D1(\spm_in[SDATA][12] ), .S0(n134), .Z(
        n273) );
  HS65_LS_MUX21I1X6 U784 ( .D0(n424), .D1(\spm_in[SDATA][13] ), .S0(n133), .Z(
        n274) );
  HS65_LS_MUX21I1X6 U785 ( .D0(n425), .D1(\spm_in[SDATA][14] ), .S0(n136), .Z(
        n275) );
  HS65_LS_MUX21I1X6 U786 ( .D0(n426), .D1(\spm_in[SDATA][15] ), .S0(n133), .Z(
        n276) );
  HS65_LS_MUX21I1X6 U787 ( .D0(n427), .D1(\spm_in[SDATA][16] ), .S0(n136), .Z(
        n277) );
  HS65_LS_MUX21I1X6 U788 ( .D0(n428), .D1(\spm_in[SDATA][17] ), .S0(n134), .Z(
        n278) );
  HS65_LS_MUX21I1X6 U789 ( .D0(n429), .D1(\spm_in[SDATA][18] ), .S0(n133), .Z(
        n279) );
  HS65_LS_MUX21I1X6 U790 ( .D0(n430), .D1(\spm_in[SDATA][19] ), .S0(n136), .Z(
        n280) );
  HS65_LS_MUX21I1X6 U791 ( .D0(n431), .D1(\spm_in[SDATA][20] ), .S0(n134), .Z(
        n281) );
  HS65_LS_MUX21I1X6 U792 ( .D0(n432), .D1(\spm_in[SDATA][21] ), .S0(n133), .Z(
        n282) );
  HS65_LS_MUX21I1X6 U793 ( .D0(n433), .D1(\spm_in[SDATA][22] ), .S0(n136), .Z(
        n283) );
  HS65_LS_MUX21I1X6 U794 ( .D0(n434), .D1(\spm_in[SDATA][23] ), .S0(n134), .Z(
        n284) );
  HS65_LS_MUX21I1X6 U795 ( .D0(n435), .D1(\spm_in[SDATA][24] ), .S0(n133), .Z(
        n285) );
  HS65_LS_MUX21I1X6 U796 ( .D0(n436), .D1(\spm_in[SDATA][25] ), .S0(n136), .Z(
        n286) );
  HS65_LS_MUX21I1X6 U797 ( .D0(n437), .D1(\spm_in[SDATA][26] ), .S0(n134), .Z(
        n287) );
  HS65_LS_MUX21I1X6 U798 ( .D0(n438), .D1(\spm_in[SDATA][27] ), .S0(n134), .Z(
        n288) );
  HS65_LS_MUX21I1X6 U799 ( .D0(n439), .D1(\spm_in[SDATA][28] ), .S0(n133), .Z(
        n289) );
  HS65_LS_MUX21I1X6 U800 ( .D0(n440), .D1(\spm_in[SDATA][29] ), .S0(n136), .Z(
        n290) );
  HS65_LS_MUX21I1X6 U801 ( .D0(n441), .D1(\spm_in[SDATA][30] ), .S0(n134), .Z(
        n291) );
  HS65_LS_MUX21I1X6 U802 ( .D0(n442), .D1(\spm_in[SDATA][31] ), .S0(n133), .Z(
        n292) );
  HS65_LS_IVX9 U803 ( .A(\phase_next[1] ), .Z(n452) );
  HS65_LS_IVX9 U804 ( .A(phitOut1[0]), .Z(n467) );
  HS65_LS_IVX9 U805 ( .A(phitOut0[0]), .Z(n466) );
  HS65_LS_IVX9 U806 ( .A(phitOut1[1]), .Z(n470) );
  HS65_LS_IVX9 U807 ( .A(phitOut0[1]), .Z(n469) );
  HS65_LS_IVX9 U808 ( .A(phitOut1[2]), .Z(n474) );
  HS65_LS_IVX9 U809 ( .A(phitOut0[2]), .Z(n473) );
  HS65_LS_IVX9 U810 ( .A(phitOut1[3]), .Z(n478) );
  HS65_LS_IVX9 U811 ( .A(phitOut0[3]), .Z(n477) );
  HS65_LS_IVX9 U812 ( .A(phitOut1[4]), .Z(n481) );
  HS65_LS_IVX9 U813 ( .A(phitOut0[4]), .Z(n480) );
  HS65_LS_OAI212X5 U814 ( .A(n481), .B(n114), .C(n27), .D(n480), .E(n479), .Z(
        pkt_out[4]) );
  HS65_LS_IVX9 U815 ( .A(phitOut1[5]), .Z(n484) );
  HS65_LS_IVX9 U816 ( .A(phitOut0[5]), .Z(n483) );
  HS65_LS_OAI212X5 U817 ( .A(n116), .B(n484), .C(n27), .D(n483), .E(n482), .Z(
        pkt_out[5]) );
  HS65_LS_IVX9 U818 ( .A(phitOut1[6]), .Z(n487) );
  HS65_LS_IVX9 U819 ( .A(phitOut0[6]), .Z(n486) );
  HS65_LS_OAI212X5 U820 ( .A(n113), .B(n487), .C(n27), .D(n486), .E(n485), .Z(
        pkt_out[6]) );
  HS65_LS_IVX9 U821 ( .A(phitOut1[7]), .Z(n490) );
  HS65_LS_IVX9 U822 ( .A(phitOut0[7]), .Z(n489) );
  HS65_LS_IVX9 U823 ( .A(phitOut1[8]), .Z(n493) );
  HS65_LS_IVX9 U824 ( .A(phitOut0[8]), .Z(n492) );
  HS65_LS_OAI212X5 U825 ( .A(n113), .B(n493), .C(n27), .D(n492), .E(n491), .Z(
        pkt_out[8]) );
  HS65_LS_IVX9 U826 ( .A(phitOut1[9]), .Z(n496) );
  HS65_LS_IVX9 U827 ( .A(phitOut0[9]), .Z(n495) );
  HS65_LS_OAI212X5 U828 ( .A(n496), .B(n113), .C(n27), .D(n495), .E(n494), .Z(
        pkt_out[9]) );
  HS65_LS_IVX9 U829 ( .A(phitOut1[10]), .Z(n499) );
  HS65_LS_IVX9 U830 ( .A(phitOut0[10]), .Z(n498) );
  HS65_LS_IVX9 U831 ( .A(phitOut1[11]), .Z(n502) );
  HS65_LS_IVX9 U832 ( .A(phitOut0[11]), .Z(n501) );
  HS65_LS_IVX9 U833 ( .A(phitOut1[12]), .Z(n505) );
  HS65_LS_IVX9 U834 ( .A(phitOut0[12]), .Z(n504) );
  HS65_LS_NAND2X7 U835 ( .A(phitOut2[12]), .B(n471), .Z(n503) );
  HS65_LS_OAI212X5 U836 ( .A(n113), .B(n505), .C(n27), .D(n504), .E(n503), .Z(
        pkt_out[12]) );
  HS65_LS_IVX9 U837 ( .A(phitOut1[13]), .Z(n508) );
  HS65_LS_IVX9 U838 ( .A(phitOut0[13]), .Z(n507) );
  HS65_LS_IVX9 U839 ( .A(phitOut1[14]), .Z(n511) );
  HS65_LS_IVX9 U840 ( .A(phitOut0[14]), .Z(n510) );
  HS65_LS_NAND2X7 U841 ( .A(phitOut2[14]), .B(n471), .Z(n509) );
  HS65_LS_OAI212X5 U842 ( .A(n511), .B(n117), .C(n27), .D(n510), .E(n509), .Z(
        pkt_out[14]) );
  HS65_LS_IVX9 U843 ( .A(phitOut1[15]), .Z(n514) );
  HS65_LS_IVX9 U844 ( .A(phitOut0[15]), .Z(n513) );
  HS65_LS_OAI212X5 U845 ( .A(n514), .B(n114), .C(n27), .D(n513), .E(n512), .Z(
        pkt_out[15]) );
  HS65_LS_IVX9 U846 ( .A(phitOut1[16]), .Z(n517) );
  HS65_LS_IVX9 U847 ( .A(phitOut0[16]), .Z(n516) );
  HS65_LS_OAI212X5 U848 ( .A(n116), .B(n517), .C(n27), .D(n516), .E(n515), .Z(
        pkt_out[16]) );
  HS65_LS_IVX9 U849 ( .A(phitOut1[17]), .Z(n520) );
  HS65_LS_IVX9 U850 ( .A(phitOut0[17]), .Z(n519) );
  HS65_LS_NAND2X7 U851 ( .A(phitOut2[17]), .B(n471), .Z(n518) );
  HS65_LS_OAI212X5 U852 ( .A(n113), .B(n520), .C(n27), .D(n519), .E(n518), .Z(
        pkt_out[17]) );
  HS65_LS_IVX9 U853 ( .A(phitOut1[18]), .Z(n523) );
  HS65_LS_IVX9 U854 ( .A(phitOut0[18]), .Z(n522) );
  HS65_LS_IVX9 U855 ( .A(phitOut1[19]), .Z(n527) );
  HS65_LS_IVX9 U856 ( .A(phitOut0[19]), .Z(n525) );
  HS65_LS_IVX9 U857 ( .A(phitOut1[20]), .Z(n530) );
  HS65_LS_IVX9 U858 ( .A(phitOut0[20]), .Z(n529) );
  HS65_LS_OAI212X5 U859 ( .A(n530), .B(n114), .C(n18), .D(n529), .E(n528), .Z(
        pkt_out[20]) );
  HS65_LS_IVX9 U860 ( .A(phitOut1[21]), .Z(n533) );
  HS65_LS_IVX9 U861 ( .A(phitOut0[21]), .Z(n532) );
  HS65_LS_NAND2X7 U862 ( .A(phitOut2[21]), .B(n471), .Z(n531) );
  HS65_LS_OAI212X5 U863 ( .A(n113), .B(n533), .C(n3), .D(n532), .E(n531), .Z(
        pkt_out[21]) );
  HS65_LS_IVX9 U864 ( .A(phitOut1[22]), .Z(n536) );
  HS65_LS_IVX9 U865 ( .A(phitOut0[22]), .Z(n535) );
  HS65_LS_NAND2X7 U866 ( .A(phitOut2[22]), .B(n471), .Z(n534) );
  HS65_LS_OAI212X5 U867 ( .A(n113), .B(n536), .C(n18), .D(n535), .E(n534), .Z(
        pkt_out[22]) );
  HS65_LS_IVX9 U868 ( .A(phitOut1[23]), .Z(n539) );
  HS65_LS_IVX9 U869 ( .A(phitOut0[23]), .Z(n538) );
  HS65_LS_NAND2X7 U870 ( .A(phitOut2[23]), .B(n471), .Z(n537) );
  HS65_LS_IVX9 U871 ( .A(phitOut1[24]), .Z(n542) );
  HS65_LS_IVX9 U872 ( .A(phitOut0[24]), .Z(n541) );
  HS65_LS_NAND2X7 U873 ( .A(phitOut2[24]), .B(n471), .Z(n540) );
  HS65_LS_IVX9 U874 ( .A(phitOut1[25]), .Z(n545) );
  HS65_LS_IVX9 U875 ( .A(phitOut0[25]), .Z(n544) );
  HS65_LS_IVX9 U876 ( .A(phitOut1[26]), .Z(n548) );
  HS65_LS_IVX9 U877 ( .A(phitOut0[26]), .Z(n547) );
  HS65_LS_NAND2X7 U878 ( .A(phitOut2[26]), .B(n471), .Z(n546) );
  HS65_LS_OAI212X5 U879 ( .A(n113), .B(n548), .C(n3), .D(n547), .E(n546), .Z(
        pkt_out[26]) );
  HS65_LS_IVX9 U880 ( .A(phitOut1[27]), .Z(n551) );
  HS65_LS_IVX9 U881 ( .A(phitOut0[27]), .Z(n550) );
  HS65_LS_IVX9 U882 ( .A(phitOut1[28]), .Z(n554) );
  HS65_LS_IVX9 U883 ( .A(phitOut0[28]), .Z(n553) );
  HS65_LS_OAI212X5 U884 ( .A(n116), .B(n554), .C(n18), .D(n553), .E(n552), .Z(
        pkt_out[28]) );
  HS65_LS_IVX9 U885 ( .A(phitOut1[29]), .Z(n557) );
  HS65_LS_IVX9 U886 ( .A(phitOut0[29]), .Z(n556) );
  HS65_LS_OAI212X5 U887 ( .A(n116), .B(n557), .C(n3), .D(n556), .E(n555), .Z(
        pkt_out[29]) );
  HS65_LS_IVX9 U888 ( .A(phitOut1[30]), .Z(n560) );
  HS65_LS_IVX9 U889 ( .A(phitOut0[30]), .Z(n559) );
  HS65_LS_OAI212X5 U890 ( .A(n113), .B(n560), .C(n559), .D(n18), .E(n558), .Z(
        pkt_out[30]) );
  HS65_LS_IVX9 U891 ( .A(phitOut1[31]), .Z(n563) );
  HS65_LS_IVX9 U892 ( .A(phitOut0[31]), .Z(n562) );
  HS65_LS_NAND2X7 U893 ( .A(phitOut2[31]), .B(n471), .Z(n561) );
  HS65_LS_OAI212X5 U894 ( .A(n113), .B(n563), .C(n3), .D(n562), .E(n561), .Z(
        pkt_out[31]) );
  HS65_LS_IVX9 U895 ( .A(phitOut1[32]), .Z(n566) );
  HS65_LS_IVX9 U896 ( .A(phitOut0[32]), .Z(n565) );
  HS65_LS_OAI212X5 U897 ( .A(n113), .B(n566), .C(n565), .D(n18), .E(n564), .Z(
        pkt_out[32]) );
  HS65_LS_IVX9 U898 ( .A(phitOut1[33]), .Z(n569) );
  HS65_LS_IVX9 U899 ( .A(phitOut0[33]), .Z(n568) );
  HS65_LS_OAI212X5 U900 ( .A(n116), .B(n569), .C(n3), .D(n568), .E(n567), .Z(
        pkt_out[33]) );
  HS65_LS_IVX9 U901 ( .A(phitOut1[34]), .Z(n572) );
  HS65_LS_IVX9 U902 ( .A(flit_buf[64]), .Z(n575) );
  HS65_LS_OAI22X6 U903 ( .A(n354), .B(n576), .C(n589), .D(n575), .Z(
        \spm_out[MADDR][0] ) );
  HS65_LS_IVX9 U904 ( .A(flit_buf[65]), .Z(n577) );
  HS65_LS_OAI22X6 U905 ( .A(n354), .B(n578), .C(n589), .D(n577), .Z(
        \spm_out[MADDR][1] ) );
  HS65_LS_IVX9 U906 ( .A(flit_buf[66]), .Z(n579) );
  HS65_LS_OAI22X6 U907 ( .A(n354), .B(n580), .C(n589), .D(n579), .Z(
        \spm_out[MADDR][2] ) );
  HS65_LS_IVX9 U908 ( .A(flit_buf[67]), .Z(n581) );
  HS65_LS_OAI22X6 U909 ( .A(n354), .B(n582), .C(n589), .D(n581), .Z(
        \spm_out[MADDR][3] ) );
  HS65_LS_IVX9 U910 ( .A(flit_buf[68]), .Z(n583) );
  HS65_LS_OAI22X6 U911 ( .A(n354), .B(n584), .C(n589), .D(n583), .Z(
        \spm_out[MADDR][4] ) );
  HS65_LS_IVX9 U912 ( .A(flit_buf[69]), .Z(n585) );
  HS65_LS_OAI22X6 U913 ( .A(n354), .B(n586), .C(n589), .D(n585), .Z(
        \spm_out[MADDR][5] ) );
  HS65_LS_IVX9 U914 ( .A(flit_buf[70]), .Z(n587) );
  HS65_LS_OAI22X6 U915 ( .A(n588), .B(n354), .C(n589), .D(n587), .Z(
        \spm_out[MADDR][6] ) );
  HS65_LS_IVX9 U916 ( .A(n589), .Z(\spm_out[MCMD][0] ) );
  HS65_LS_IVX9 U917 ( .A(n590), .Z(n592) );
  HS65_LS_OAI112X5 U918 ( .A(n38), .B(n592), .C(n40), .D(n591), .Z(
        \proc_out[SCMDACCEPT] ) );
endmodule


module latch_controller_1_0 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_0 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n1, n2, n3, n4;
  assign N0 = preset;

  latch_controller_1_0 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n4), .RN(n3), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n3), .Z(n2) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n1) );
  HS65_LS_OR2X9 U8 ( .A(n1), .B(n2), .Z(N5) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_IVX9 U3 ( .A(lt_enable), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(N0), .Z(n3) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n4), .Z(lt_gated) );
endmodule


module latch_controller_1_39 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_39 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n3, n4, n5, n6;
  assign N0 = preset;

  latch_controller_1_39 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n4), .RN(n3), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n3), .Z(n5) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n6), .B(n5), .Z(N5) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_IVX9 U3 ( .A(lt_enable), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(N0), .Z(n3) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n4), .Z(lt_gated) );
endmodule


module latch_controller_1_38 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_38 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n3, n4, n5, n6;
  assign N0 = preset;

  latch_controller_1_38 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n4), .RN(n3), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n3), .Z(n5) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n6), .B(n5), .Z(N5) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_IVX9 U3 ( .A(lt_enable), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(N0), .Z(n3) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n4), .Z(lt_gated) );
endmodule


module latch_controller_1_37 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_37 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n3, n4, n5, n6;
  assign N0 = preset;

  latch_controller_1_37 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n4), .RN(n3), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n3), .Z(n5) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n6), .B(n5), .Z(N5) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_IVX9 U3 ( .A(lt_enable), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(N0), .Z(n3) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n4), .Z(lt_gated) );
endmodule


module latch_controller_1_36 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_NOR2AX3 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_36 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n3, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_36 controller ( .preset(n3), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLRQX18 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(n3), .Z(n7) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_LDHQX18 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX18 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX18 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX18 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX18 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX18 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX18 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX18 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX18 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX18 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX18 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX18 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX18 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX18 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX18 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX18 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX18 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX18 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX18 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX4 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX18 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX18 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX18 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX4 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX4 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX18 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX18 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX18 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX18 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX18 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX18 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX18 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX18 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX18 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_IVX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_IVX9 U5 ( .A(N0), .Z(n4) );
  HS65_LS_NAND2X7 U9 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_comb_0_0_0 ( data_valid, data_in, preset, data_out, sel );
  input [34:0] data_in;
  output [34:0] data_out;
  output [4:0] sel;
  input data_valid, preset;
  wire   data_in_34, data_in_33, data_in_32, \data_in[31] , \data_in[30] ,
         \data_in[29] , \data_in[28] , \data_in[27] , \data_in[26] ,
         \data_in[25] , \data_in[24] , \data_in[23] , \data_in[22] ,
         \data_in[21] , \data_in[20] , \data_in[19] , \data_in[18] ,
         \data_in[17] , \data_in[16] , N23, N25, N26, N27, N28, n19, n20, n21,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;
  assign data_out[34] = data_in_34;
  assign data_in_34 = data_in[34];
  assign data_out[33] = data_in_33;
  assign data_in_33 = data_in[33];
  assign data_out[32] = data_in_32;
  assign data_in_32 = data_in[32];
  assign data_out[31] = \data_in[31] ;
  assign \data_in[31]  = data_in[31];
  assign data_out[30] = \data_in[30] ;
  assign \data_in[30]  = data_in[30];
  assign data_out[29] = \data_in[29] ;
  assign \data_in[29]  = data_in[29];
  assign data_out[28] = \data_in[28] ;
  assign \data_in[28]  = data_in[28];
  assign data_out[27] = \data_in[27] ;
  assign \data_in[27]  = data_in[27];
  assign data_out[26] = \data_in[26] ;
  assign \data_in[26]  = data_in[26];
  assign data_out[25] = \data_in[25] ;
  assign \data_in[25]  = data_in[25];
  assign data_out[24] = \data_in[24] ;
  assign \data_in[24]  = data_in[24];
  assign data_out[23] = \data_in[23] ;
  assign \data_in[23]  = data_in[23];
  assign data_out[22] = \data_in[22] ;
  assign \data_in[22]  = data_in[22];
  assign data_out[21] = \data_in[21] ;
  assign \data_in[21]  = data_in[21];
  assign data_out[20] = \data_in[20] ;
  assign \data_in[20]  = data_in[20];
  assign data_out[19] = \data_in[19] ;
  assign \data_in[19]  = data_in[19];
  assign data_out[18] = \data_in[18] ;
  assign \data_in[18]  = data_in[18];
  assign data_out[17] = \data_in[17] ;
  assign \data_in[17]  = data_in[17];
  assign data_out[16] = \data_in[16] ;
  assign \data_in[16]  = data_in[16];
  assign sel[0] = 1'b0;

  HS65_LS_LDHQX9 \sel_reg[4]  ( .G(N23), .D(N28), .Q(sel[4]) );
  HS65_LS_LDHQX9 \sel_reg[3]  ( .G(N23), .D(N27), .Q(sel[3]) );
  HS65_LS_LDHQX9 \sel_reg[2]  ( .G(N23), .D(N26), .Q(sel[2]) );
  HS65_LS_LDHQX9 \sel_reg[1]  ( .G(N23), .D(N25), .Q(sel[1]) );
  HS65_LS_NAND3AX6 U4 ( .A(preset), .B(n20), .C(n2), .Z(n21) );
  HS65_LS_OAI22X6 U5 ( .A(n9), .B(n19), .C(n2), .D(n11), .Z(data_out[7]) );
  HS65_LS_OAI22X6 U6 ( .A(n19), .B(n16), .C(n2), .D(n18), .Z(data_out[0]) );
  HS65_LS_OAI22X6 U7 ( .A(n19), .B(n15), .C(n2), .D(n17), .Z(data_out[1]) );
  HS65_LS_OAI22X6 U8 ( .A(n19), .B(n14), .C(n2), .D(n16), .Z(data_out[2]) );
  HS65_LS_OAI22X6 U9 ( .A(n19), .B(n13), .C(n2), .D(n15), .Z(data_out[3]) );
  HS65_LS_OAI22X6 U10 ( .A(n19), .B(n12), .C(n2), .D(n14), .Z(data_out[4]) );
  HS65_LS_OAI22X6 U11 ( .A(n19), .B(n11), .C(n2), .D(n13), .Z(data_out[5]) );
  HS65_LS_OAI22X6 U12 ( .A(n19), .B(n10), .C(n2), .D(n12), .Z(data_out[6]) );
  HS65_LS_OAI22X6 U13 ( .A(n19), .B(n8), .C(n2), .D(n10), .Z(data_out[8]) );
  HS65_LS_OAI22X6 U14 ( .A(n19), .B(n7), .C(n2), .D(n9), .Z(data_out[9]) );
  HS65_LS_OAI22X6 U15 ( .A(n19), .B(n6), .C(n2), .D(n8), .Z(data_out[10]) );
  HS65_LS_OAI22X6 U16 ( .A(n19), .B(n5), .C(n2), .D(n7), .Z(data_out[11]) );
  HS65_LS_OAI22X6 U17 ( .A(n19), .B(n4), .C(n2), .D(n6), .Z(data_out[12]) );
  HS65_LS_OAI22X6 U18 ( .A(n19), .B(n3), .C(n2), .D(n5), .Z(data_out[13]) );
  HS65_LS_IVX9 U19 ( .A(n19), .Z(n2) );
  HS65_LS_NOR3X4 U20 ( .A(n20), .B(preset), .C(n19), .Z(N28) );
  HS65_LS_NOR3X4 U21 ( .A(n21), .B(n17), .C(n18), .Z(N27) );
  HS65_LS_NAND2X7 U22 ( .A(n17), .B(n18), .Z(n20) );
  HS65_LS_NOR2X6 U23 ( .A(n2), .B(n4), .Z(data_out[14]) );
  HS65_LS_NOR2X6 U24 ( .A(n2), .B(n3), .Z(data_out[15]) );
  HS65_LS_NAND2X14 U25 ( .A(data_in_34), .B(data_in_33), .Z(n19) );
  HS65_LS_IVX9 U26 ( .A(data_in[1]), .Z(n17) );
  HS65_LS_IVX9 U27 ( .A(data_in[0]), .Z(n18) );
  HS65_LS_NOR2X6 U28 ( .A(data_in[1]), .B(n21), .Z(N25) );
  HS65_LS_NOR2X6 U29 ( .A(data_in[0]), .B(n21), .Z(N26) );
  HS65_LS_IVX9 U30 ( .A(data_in[9]), .Z(n9) );
  HS65_LS_IVX9 U31 ( .A(data_in[2]), .Z(n16) );
  HS65_LS_IVX9 U32 ( .A(data_in[3]), .Z(n15) );
  HS65_LS_IVX9 U33 ( .A(data_in[4]), .Z(n14) );
  HS65_LS_IVX9 U34 ( .A(data_in[5]), .Z(n13) );
  HS65_LS_IVX9 U35 ( .A(data_in[6]), .Z(n12) );
  HS65_LS_IVX9 U36 ( .A(data_in[7]), .Z(n11) );
  HS65_LS_IVX9 U37 ( .A(data_in[8]), .Z(n10) );
  HS65_LS_IVX9 U38 ( .A(data_in[10]), .Z(n8) );
  HS65_LS_IVX9 U39 ( .A(data_in[11]), .Z(n7) );
  HS65_LS_IVX9 U40 ( .A(data_in[12]), .Z(n6) );
  HS65_LS_IVX9 U41 ( .A(data_in[13]), .Z(n5) );
  HS65_LS_IVX9 U42 ( .A(data_in[14]), .Z(n4) );
  HS65_LS_IVX9 U43 ( .A(data_in[15]), .Z(n3) );
  HS65_LS_CB4I6X9 U44 ( .A(n2), .B(n1), .C(data_valid), .D(preset), .Z(N23) );
  HS65_LS_IVX9 U45 ( .A(data_in_34), .Z(n1) );
endmodule


module latch_controller_1_20 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_20 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_20 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n7) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_IVX9 U3 ( .A(N0), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_0_0_0 ( preset, .chan_in_f({\chan_in_f[REQ] , \chan_in_f[DATA][34] , 
        \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , 
        \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , 
        \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , 
        \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , 
        \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , 
        \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , 
        \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , 
        \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , 
        \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , 
        \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , 
        \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , 
        \chan_in_f[DATA][0] }), .chan_in_b(\chan_in_b[ACK] ), .chan_out_f({
        \chan_out_f[REQ] , \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , 
        \chan_out_f[DATA][32] , \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , 
        \chan_out_f[DATA][29] , \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , 
        \chan_out_f[DATA][26] , \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , 
        \chan_out_f[DATA][23] , \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , 
        \chan_out_f[DATA][20] , \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , 
        \chan_out_f[DATA][17] , \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , 
        \chan_out_f[DATA][14] , \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , 
        \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , 
        \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , 
        \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , 
        \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), 
    .chan_out_b(\chan_out_b[ACK] ), sel );
  output [4:0] sel;
  input preset, \chan_in_f[REQ] , \chan_in_f[DATA][34] , \chan_in_f[DATA][33] ,
         \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , \chan_in_f[DATA][30] ,
         \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , \chan_in_f[DATA][27] ,
         \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , \chan_in_f[DATA][24] ,
         \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , \chan_in_f[DATA][21] ,
         \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , \chan_in_f[DATA][18] ,
         \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , \chan_in_f[DATA][15] ,
         \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , \chan_in_f[DATA][12] ,
         \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , \chan_in_f[DATA][9] ,
         \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , \chan_in_f[DATA][6] ,
         \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , \chan_in_f[DATA][3] ,
         \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , \chan_in_f[DATA][0] ,
         \chan_out_b[ACK] ;
  output \chan_in_b[ACK] , \chan_out_f[REQ] , \chan_out_f[DATA][34] ,
         \chan_out_f[DATA][33] , \chan_out_f[DATA][32] ,
         \chan_out_f[DATA][31] , \chan_out_f[DATA][30] ,
         \chan_out_f[DATA][29] , \chan_out_f[DATA][28] ,
         \chan_out_f[DATA][27] , \chan_out_f[DATA][26] ,
         \chan_out_f[DATA][25] , \chan_out_f[DATA][24] ,
         \chan_out_f[DATA][23] , \chan_out_f[DATA][22] ,
         \chan_out_f[DATA][21] , \chan_out_f[DATA][20] ,
         \chan_out_f[DATA][19] , \chan_out_f[DATA][18] ,
         \chan_out_f[DATA][17] , \chan_out_f[DATA][16] ,
         \chan_out_f[DATA][15] , \chan_out_f[DATA][14] ,
         \chan_out_f[DATA][13] , \chan_out_f[DATA][12] ,
         \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] ,
         \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] ,
         \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] ,
         \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] ;
  wire   \chan_internal_f[REQ] , \chan_internal_f[DATA][34] ,
         \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] ,
         \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] ,
         \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] ,
         \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] ,
         \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] ,
         \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] ,
         \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] ,
         \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] ,
         \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] ,
         \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] ,
         \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] ,
         \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] ,
         \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] ,
         \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] ,
         \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] ,
         \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] ,
         \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] , req_n, lt_en,
         n1, n2, n3, n4, n5, n6, n7;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign sel[0] = 1'b0;

  hpu_comb_0_0_0 hpu_combinatorial ( .data_valid(lt_en), .data_in({
        \chan_in_f[DATA][34] , \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , 
        \chan_in_f[DATA][31] , \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , 
        \chan_in_f[DATA][28] , \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , 
        \chan_in_f[DATA][25] , \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , 
        \chan_in_f[DATA][22] , \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , 
        \chan_in_f[DATA][19] , \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , 
        \chan_in_f[DATA][16] , \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , 
        \chan_in_f[DATA][13] , \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , 
        \chan_in_f[DATA][10] , \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , 
        \chan_in_f[DATA][7] , \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , 
        \chan_in_f[DATA][4] , \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , 
        \chan_in_f[DATA][1] , \chan_in_f[DATA][0] }), .preset(n7), .data_out({
        \chan_internal_f[DATA][34] , \chan_internal_f[DATA][33] , 
        \chan_internal_f[DATA][32] , \chan_internal_f[DATA][31] , 
        \chan_internal_f[DATA][30] , \chan_internal_f[DATA][29] , 
        \chan_internal_f[DATA][28] , \chan_internal_f[DATA][27] , 
        \chan_internal_f[DATA][26] , \chan_internal_f[DATA][25] , 
        \chan_internal_f[DATA][24] , \chan_internal_f[DATA][23] , 
        \chan_internal_f[DATA][22] , \chan_internal_f[DATA][21] , 
        \chan_internal_f[DATA][20] , \chan_internal_f[DATA][19] , 
        \chan_internal_f[DATA][18] , \chan_internal_f[DATA][17] , 
        \chan_internal_f[DATA][16] , \chan_internal_f[DATA][15] , 
        \chan_internal_f[DATA][14] , \chan_internal_f[DATA][13] , 
        \chan_internal_f[DATA][12] , \chan_internal_f[DATA][11] , 
        \chan_internal_f[DATA][10] , \chan_internal_f[DATA][9] , 
        \chan_internal_f[DATA][8] , \chan_internal_f[DATA][7] , 
        \chan_internal_f[DATA][6] , \chan_internal_f[DATA][5] , 
        \chan_internal_f[DATA][4] , \chan_internal_f[DATA][3] , 
        \chan_internal_f[DATA][2] , \chan_internal_f[DATA][1] , 
        \chan_internal_f[DATA][0] }), .sel({sel[4:1], SYNOPSYS_UNCONNECTED__0}) );
  channel_latch_1_xxxxxxxxx_20 token_latch ( .preset(n7), .left_in({
        \chan_internal_f[REQ] , \chan_internal_f[DATA][34] , 
        \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] , 
        \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] , 
        \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] , 
        \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] , 
        \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] , 
        \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] , 
        \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] , 
        \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] , 
        \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] , 
        \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] , 
        \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] , 
        \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] , 
        \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] , 
        \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] , 
        \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] , 
        \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] , 
        \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] }), .left_out(
        \chan_in_b[ACK] ), .right_out({\chan_out_f[REQ] , 
        \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , \chan_out_f[DATA][32] , 
        \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , \chan_out_f[DATA][29] , 
        \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , \chan_out_f[DATA][26] , 
        \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , \chan_out_f[DATA][23] , 
        \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , \chan_out_f[DATA][20] , 
        \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , \chan_out_f[DATA][17] , 
        \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , \chan_out_f[DATA][14] , 
        \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , \chan_out_f[DATA][11] , 
        \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , \chan_out_f[DATA][8] , 
        \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , \chan_out_f[DATA][5] , 
        \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , \chan_out_f[DATA][2] , 
        \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), .right_in(
        \chan_out_b[ACK] ), .lt_enable(lt_en) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chan_internal_f[REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(\chan_in_f[REQ] ), .Z(req_n) );
  HS65_LS_BFX9 U1 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U2 ( .A(n3), .Z(n2) );
  HS65_LS_BFX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_BFX9 U4 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U6 ( .A(req_n), .Z(n6) );
  HS65_LS_BFX9 U7 ( .A(preset), .Z(n7) );
endmodule


module hpu_comb_0_2_0 ( data_valid, data_in, preset, data_out, sel );
  input [34:0] data_in;
  output [34:0] data_out;
  output [4:0] sel;
  input data_valid, preset;
  wire   data_in_34, data_in_33, data_in_32, \data_in[31] , \data_in[30] ,
         \data_in[29] , \data_in[28] , \data_in[27] , \data_in[26] ,
         \data_in[25] , \data_in[24] , \data_in[23] , \data_in[22] ,
         \data_in[21] , \data_in[20] , \data_in[19] , \data_in[18] ,
         \data_in[17] , \data_in[16] , N26, N27, N28, N30, N31, n11, n12, n13,
         n14, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  assign data_out[34] = data_in_34;
  assign data_in_34 = data_in[34];
  assign data_out[33] = data_in_33;
  assign data_in_33 = data_in[33];
  assign data_out[32] = data_in_32;
  assign data_in_32 = data_in[32];
  assign data_out[31] = \data_in[31] ;
  assign \data_in[31]  = data_in[31];
  assign data_out[30] = \data_in[30] ;
  assign \data_in[30]  = data_in[30];
  assign data_out[29] = \data_in[29] ;
  assign \data_in[29]  = data_in[29];
  assign data_out[28] = \data_in[28] ;
  assign \data_in[28]  = data_in[28];
  assign data_out[27] = \data_in[27] ;
  assign \data_in[27]  = data_in[27];
  assign data_out[26] = \data_in[26] ;
  assign \data_in[26]  = data_in[26];
  assign data_out[25] = \data_in[25] ;
  assign \data_in[25]  = data_in[25];
  assign data_out[24] = \data_in[24] ;
  assign \data_in[24]  = data_in[24];
  assign data_out[23] = \data_in[23] ;
  assign \data_in[23]  = data_in[23];
  assign data_out[22] = \data_in[22] ;
  assign \data_in[22]  = data_in[22];
  assign data_out[21] = \data_in[21] ;
  assign \data_in[21]  = data_in[21];
  assign data_out[20] = \data_in[20] ;
  assign \data_in[20]  = data_in[20];
  assign data_out[19] = \data_in[19] ;
  assign \data_in[19]  = data_in[19];
  assign data_out[18] = \data_in[18] ;
  assign \data_in[18]  = data_in[18];
  assign data_out[17] = \data_in[17] ;
  assign \data_in[17]  = data_in[17];
  assign data_out[16] = \data_in[16] ;
  assign \data_in[16]  = data_in[16];
  assign sel[2] = 1'b0;

  HS65_LS_LDHQX9 \sel_reg[4]  ( .G(N26), .D(N31), .Q(sel[4]) );
  HS65_LS_LDHQX9 \sel_reg[3]  ( .G(N26), .D(N30), .Q(sel[3]) );
  HS65_LS_LDHQX9 \sel_reg[1]  ( .G(N26), .D(N28), .Q(sel[1]) );
  HS65_LS_LDHQX9 \sel_reg[0]  ( .G(N26), .D(N27), .Q(sel[0]) );
  HS65_LS_OAI22X6 U4 ( .A(n11), .B(n9), .C(n2), .D(n10), .Z(data_out[0]) );
  HS65_LS_OAI22X6 U5 ( .A(n11), .B(n8), .C(n2), .D(n9), .Z(data_out[2]) );
  HS65_LS_OAI22X6 U6 ( .A(n11), .B(n7), .C(n2), .D(n8), .Z(data_out[4]) );
  HS65_LS_OAI22X6 U7 ( .A(n11), .B(n6), .C(n2), .D(n7), .Z(data_out[6]) );
  HS65_LS_OAI22X6 U8 ( .A(n11), .B(n5), .C(n2), .D(n6), .Z(data_out[8]) );
  HS65_LS_OAI22X6 U9 ( .A(n11), .B(n4), .C(n2), .D(n5), .Z(data_out[10]) );
  HS65_LS_OAI22X6 U10 ( .A(n11), .B(n3), .C(n2), .D(n4), .Z(data_out[12]) );
  HS65_LS_NAND3AX6 U11 ( .A(preset), .B(n12), .C(n2), .Z(n13) );
  HS65_LS_NOR3X4 U12 ( .A(n12), .B(preset), .C(n11), .Z(N31) );
  HS65_LS_IVX9 U13 ( .A(n11), .Z(n2) );
  HS65_LS_NOR3X4 U14 ( .A(n13), .B(n10), .C(n14), .Z(N30) );
  HS65_LS_NOR2AX3 U15 ( .A(n14), .B(n13), .Z(N28) );
  HS65_LS_NOR2X6 U16 ( .A(n2), .B(n3), .Z(data_out[14]) );
  HS65_LS_NAND2X14 U17 ( .A(data_in_34), .B(data_in_33), .Z(n11) );
  HS65_LS_IVX9 U18 ( .A(data_in[0]), .Z(n10) );
  HS65_LS_NAND2X7 U19 ( .A(data_in[1]), .B(n10), .Z(n12) );
  HS65_LS_NOR2X6 U20 ( .A(n10), .B(data_in[1]), .Z(n14) );
  HS65_LS_NOR2X6 U21 ( .A(data_in[0]), .B(n13), .Z(N27) );
  HS65_LS_IVX9 U22 ( .A(data_in[2]), .Z(n9) );
  HS65_LS_IVX9 U23 ( .A(data_in[4]), .Z(n8) );
  HS65_LS_IVX9 U24 ( .A(data_in[6]), .Z(n7) );
  HS65_LS_IVX9 U25 ( .A(data_in[8]), .Z(n6) );
  HS65_LS_IVX9 U26 ( .A(data_in[10]), .Z(n5) );
  HS65_LS_IVX9 U27 ( .A(data_in[12]), .Z(n4) );
  HS65_LS_IVX9 U28 ( .A(data_in[14]), .Z(n3) );
  HS65_LS_AO22X9 U29 ( .A(n2), .B(data_in[3]), .C(n11), .D(data_in[1]), .Z(
        data_out[1]) );
  HS65_LS_AO22X9 U30 ( .A(n2), .B(data_in[5]), .C(n11), .D(data_in[3]), .Z(
        data_out[3]) );
  HS65_LS_AO22X9 U31 ( .A(n2), .B(data_in[7]), .C(n11), .D(data_in[5]), .Z(
        data_out[5]) );
  HS65_LS_AO22X9 U32 ( .A(data_in[9]), .B(n2), .C(n11), .D(data_in[7]), .Z(
        data_out[7]) );
  HS65_LS_AO22X9 U33 ( .A(n2), .B(data_in[11]), .C(n11), .D(data_in[9]), .Z(
        data_out[9]) );
  HS65_LS_AO22X9 U34 ( .A(n2), .B(data_in[13]), .C(n11), .D(data_in[11]), .Z(
        data_out[11]) );
  HS65_LS_AO22X9 U35 ( .A(n2), .B(data_in[15]), .C(n11), .D(data_in[13]), .Z(
        data_out[13]) );
  HS65_LS_AND2X4 U36 ( .A(data_in[15]), .B(n11), .Z(data_out[15]) );
  HS65_LS_CB4I6X9 U37 ( .A(n2), .B(n1), .C(data_valid), .D(preset), .Z(N26) );
  HS65_LS_IVX9 U38 ( .A(data_in_34), .Z(n1) );
endmodule


module latch_controller_1_19 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_19 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_19 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n7) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_IVX9 U3 ( .A(N0), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_0_2_0 ( preset, .chan_in_f({\chan_in_f[REQ] , \chan_in_f[DATA][34] , 
        \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , 
        \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , 
        \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , 
        \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , 
        \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , 
        \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , 
        \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , 
        \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , 
        \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , 
        \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , 
        \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , 
        \chan_in_f[DATA][0] }), .chan_in_b(\chan_in_b[ACK] ), .chan_out_f({
        \chan_out_f[REQ] , \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , 
        \chan_out_f[DATA][32] , \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , 
        \chan_out_f[DATA][29] , \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , 
        \chan_out_f[DATA][26] , \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , 
        \chan_out_f[DATA][23] , \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , 
        \chan_out_f[DATA][20] , \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , 
        \chan_out_f[DATA][17] , \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , 
        \chan_out_f[DATA][14] , \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , 
        \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , 
        \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , 
        \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , 
        \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), 
    .chan_out_b(\chan_out_b[ACK] ), sel );
  output [4:0] sel;
  input preset, \chan_in_f[REQ] , \chan_in_f[DATA][34] , \chan_in_f[DATA][33] ,
         \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , \chan_in_f[DATA][30] ,
         \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , \chan_in_f[DATA][27] ,
         \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , \chan_in_f[DATA][24] ,
         \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , \chan_in_f[DATA][21] ,
         \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , \chan_in_f[DATA][18] ,
         \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , \chan_in_f[DATA][15] ,
         \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , \chan_in_f[DATA][12] ,
         \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , \chan_in_f[DATA][9] ,
         \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , \chan_in_f[DATA][6] ,
         \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , \chan_in_f[DATA][3] ,
         \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , \chan_in_f[DATA][0] ,
         \chan_out_b[ACK] ;
  output \chan_in_b[ACK] , \chan_out_f[REQ] , \chan_out_f[DATA][34] ,
         \chan_out_f[DATA][33] , \chan_out_f[DATA][32] ,
         \chan_out_f[DATA][31] , \chan_out_f[DATA][30] ,
         \chan_out_f[DATA][29] , \chan_out_f[DATA][28] ,
         \chan_out_f[DATA][27] , \chan_out_f[DATA][26] ,
         \chan_out_f[DATA][25] , \chan_out_f[DATA][24] ,
         \chan_out_f[DATA][23] , \chan_out_f[DATA][22] ,
         \chan_out_f[DATA][21] , \chan_out_f[DATA][20] ,
         \chan_out_f[DATA][19] , \chan_out_f[DATA][18] ,
         \chan_out_f[DATA][17] , \chan_out_f[DATA][16] ,
         \chan_out_f[DATA][15] , \chan_out_f[DATA][14] ,
         \chan_out_f[DATA][13] , \chan_out_f[DATA][12] ,
         \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] ,
         \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] ,
         \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] ,
         \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] ;
  wire   \chan_internal_f[REQ] , \chan_internal_f[DATA][34] ,
         \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] ,
         \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] ,
         \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] ,
         \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] ,
         \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] ,
         \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] ,
         \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] ,
         \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] ,
         \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] ,
         \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] ,
         \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] ,
         \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] ,
         \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] ,
         \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] ,
         \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] ,
         \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] ,
         \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] , req_n, lt_en,
         n1, n2, n3, n4, n5, n6, n7;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign sel[2] = 1'b0;

  hpu_comb_0_2_0 hpu_combinatorial ( .data_valid(lt_en), .data_in({
        \chan_in_f[DATA][34] , \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , 
        \chan_in_f[DATA][31] , \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , 
        \chan_in_f[DATA][28] , \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , 
        \chan_in_f[DATA][25] , \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , 
        \chan_in_f[DATA][22] , \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , 
        \chan_in_f[DATA][19] , \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , 
        \chan_in_f[DATA][16] , \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , 
        \chan_in_f[DATA][13] , \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , 
        \chan_in_f[DATA][10] , \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , 
        \chan_in_f[DATA][7] , \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , 
        \chan_in_f[DATA][4] , \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , 
        \chan_in_f[DATA][1] , \chan_in_f[DATA][0] }), .preset(n7), .data_out({
        \chan_internal_f[DATA][34] , \chan_internal_f[DATA][33] , 
        \chan_internal_f[DATA][32] , \chan_internal_f[DATA][31] , 
        \chan_internal_f[DATA][30] , \chan_internal_f[DATA][29] , 
        \chan_internal_f[DATA][28] , \chan_internal_f[DATA][27] , 
        \chan_internal_f[DATA][26] , \chan_internal_f[DATA][25] , 
        \chan_internal_f[DATA][24] , \chan_internal_f[DATA][23] , 
        \chan_internal_f[DATA][22] , \chan_internal_f[DATA][21] , 
        \chan_internal_f[DATA][20] , \chan_internal_f[DATA][19] , 
        \chan_internal_f[DATA][18] , \chan_internal_f[DATA][17] , 
        \chan_internal_f[DATA][16] , \chan_internal_f[DATA][15] , 
        \chan_internal_f[DATA][14] , \chan_internal_f[DATA][13] , 
        \chan_internal_f[DATA][12] , \chan_internal_f[DATA][11] , 
        \chan_internal_f[DATA][10] , \chan_internal_f[DATA][9] , 
        \chan_internal_f[DATA][8] , \chan_internal_f[DATA][7] , 
        \chan_internal_f[DATA][6] , \chan_internal_f[DATA][5] , 
        \chan_internal_f[DATA][4] , \chan_internal_f[DATA][3] , 
        \chan_internal_f[DATA][2] , \chan_internal_f[DATA][1] , 
        \chan_internal_f[DATA][0] }), .sel({sel[4:3], SYNOPSYS_UNCONNECTED__0, 
        sel[1:0]}) );
  channel_latch_1_xxxxxxxxx_19 token_latch ( .preset(n7), .left_in({
        \chan_internal_f[REQ] , \chan_internal_f[DATA][34] , 
        \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] , 
        \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] , 
        \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] , 
        \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] , 
        \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] , 
        \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] , 
        \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] , 
        \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] , 
        \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] , 
        \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] , 
        \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] , 
        \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] , 
        \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] , 
        \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] , 
        \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] , 
        \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] , 
        \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] }), .left_out(
        \chan_in_b[ACK] ), .right_out({\chan_out_f[REQ] , 
        \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , \chan_out_f[DATA][32] , 
        \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , \chan_out_f[DATA][29] , 
        \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , \chan_out_f[DATA][26] , 
        \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , \chan_out_f[DATA][23] , 
        \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , \chan_out_f[DATA][20] , 
        \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , \chan_out_f[DATA][17] , 
        \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , \chan_out_f[DATA][14] , 
        \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , \chan_out_f[DATA][11] , 
        \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , \chan_out_f[DATA][8] , 
        \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , \chan_out_f[DATA][5] , 
        \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , \chan_out_f[DATA][2] , 
        \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), .right_in(
        \chan_out_b[ACK] ), .lt_enable(lt_en) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chan_internal_f[REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(\chan_in_f[REQ] ), .Z(req_n) );
  HS65_LS_BFX9 U1 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U2 ( .A(n3), .Z(n2) );
  HS65_LS_BFX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_BFX9 U4 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U6 ( .A(req_n), .Z(n6) );
  HS65_LS_BFX9 U7 ( .A(preset), .Z(n7) );
endmodule


module hpu_comb_0_1_0 ( data_valid, data_in, preset, data_out, sel );
  input [34:0] data_in;
  output [34:0] data_out;
  output [4:0] sel;
  input data_valid, preset;
  wire   data_in_34, data_in_33, data_in_32, \data_in[31] , \data_in[30] ,
         \data_in[29] , \data_in[28] , \data_in[27] , \data_in[26] ,
         \data_in[25] , \data_in[24] , \data_in[23] , \data_in[22] ,
         \data_in[21] , \data_in[20] , \data_in[19] , \data_in[18] ,
         \data_in[17] , \data_in[16] , N23, N24, N26, N27, N28, n11, n12, n13,
         n14, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  assign data_out[34] = data_in_34;
  assign data_in_34 = data_in[34];
  assign data_out[33] = data_in_33;
  assign data_in_33 = data_in[33];
  assign data_out[32] = data_in_32;
  assign data_in_32 = data_in[32];
  assign data_out[31] = \data_in[31] ;
  assign \data_in[31]  = data_in[31];
  assign data_out[30] = \data_in[30] ;
  assign \data_in[30]  = data_in[30];
  assign data_out[29] = \data_in[29] ;
  assign \data_in[29]  = data_in[29];
  assign data_out[28] = \data_in[28] ;
  assign \data_in[28]  = data_in[28];
  assign data_out[27] = \data_in[27] ;
  assign \data_in[27]  = data_in[27];
  assign data_out[26] = \data_in[26] ;
  assign \data_in[26]  = data_in[26];
  assign data_out[25] = \data_in[25] ;
  assign \data_in[25]  = data_in[25];
  assign data_out[24] = \data_in[24] ;
  assign \data_in[24]  = data_in[24];
  assign data_out[23] = \data_in[23] ;
  assign \data_in[23]  = data_in[23];
  assign data_out[22] = \data_in[22] ;
  assign \data_in[22]  = data_in[22];
  assign data_out[21] = \data_in[21] ;
  assign \data_in[21]  = data_in[21];
  assign data_out[20] = \data_in[20] ;
  assign \data_in[20]  = data_in[20];
  assign data_out[19] = \data_in[19] ;
  assign \data_in[19]  = data_in[19];
  assign data_out[18] = \data_in[18] ;
  assign \data_in[18]  = data_in[18];
  assign data_out[17] = \data_in[17] ;
  assign \data_in[17]  = data_in[17];
  assign data_out[16] = \data_in[16] ;
  assign \data_in[16]  = data_in[16];
  assign sel[1] = 1'b0;

  HS65_LS_LDHQX9 \sel_reg[4]  ( .G(N23), .D(N28), .Q(sel[4]) );
  HS65_LS_LDHQX9 \sel_reg[3]  ( .G(N23), .D(N27), .Q(sel[3]) );
  HS65_LS_LDHQX9 \sel_reg[2]  ( .G(N23), .D(N26), .Q(sel[2]) );
  HS65_LS_LDHQX9 \sel_reg[0]  ( .G(N23), .D(N24), .Q(sel[0]) );
  HS65_LS_OAI22X6 U4 ( .A(n6), .B(n11), .C(n2), .D(n7), .Z(data_out[7]) );
  HS65_LS_OAI22X6 U5 ( .A(n11), .B(n9), .C(n2), .D(n10), .Z(data_out[1]) );
  HS65_LS_OAI22X6 U6 ( .A(n11), .B(n8), .C(n2), .D(n9), .Z(data_out[3]) );
  HS65_LS_OAI22X6 U7 ( .A(n11), .B(n7), .C(n2), .D(n8), .Z(data_out[5]) );
  HS65_LS_OAI22X6 U8 ( .A(n11), .B(n5), .C(n2), .D(n6), .Z(data_out[9]) );
  HS65_LS_OAI22X6 U9 ( .A(n11), .B(n4), .C(n2), .D(n5), .Z(data_out[11]) );
  HS65_LS_OAI22X6 U10 ( .A(n11), .B(n3), .C(n2), .D(n4), .Z(data_out[13]) );
  HS65_LS_NAND3AX6 U11 ( .A(preset), .B(n12), .C(n2), .Z(n13) );
  HS65_LS_NOR3X4 U12 ( .A(n12), .B(preset), .C(n11), .Z(N28) );
  HS65_LS_IVX9 U13 ( .A(n11), .Z(n2) );
  HS65_LS_NOR3X4 U14 ( .A(n13), .B(n10), .C(n14), .Z(N27) );
  HS65_LS_NOR2AX3 U15 ( .A(n14), .B(n13), .Z(N26) );
  HS65_LS_NOR2X6 U16 ( .A(n2), .B(n3), .Z(data_out[15]) );
  HS65_LS_NAND2X14 U17 ( .A(data_in_34), .B(data_in_33), .Z(n11) );
  HS65_LS_IVX9 U18 ( .A(data_in[1]), .Z(n10) );
  HS65_LS_NAND2X7 U19 ( .A(data_in[0]), .B(n10), .Z(n12) );
  HS65_LS_NOR2X6 U20 ( .A(n10), .B(data_in[0]), .Z(n14) );
  HS65_LS_NOR2X6 U21 ( .A(data_in[1]), .B(n13), .Z(N24) );
  HS65_LS_IVX9 U22 ( .A(data_in[9]), .Z(n6) );
  HS65_LS_IVX9 U23 ( .A(data_in[3]), .Z(n9) );
  HS65_LS_IVX9 U24 ( .A(data_in[5]), .Z(n8) );
  HS65_LS_IVX9 U25 ( .A(data_in[7]), .Z(n7) );
  HS65_LS_IVX9 U26 ( .A(data_in[11]), .Z(n5) );
  HS65_LS_IVX9 U27 ( .A(data_in[13]), .Z(n4) );
  HS65_LS_IVX9 U28 ( .A(data_in[15]), .Z(n3) );
  HS65_LS_AO22X9 U29 ( .A(n2), .B(data_in[2]), .C(n11), .D(data_in[0]), .Z(
        data_out[0]) );
  HS65_LS_AO22X9 U30 ( .A(n2), .B(data_in[4]), .C(n11), .D(data_in[2]), .Z(
        data_out[2]) );
  HS65_LS_AO22X9 U31 ( .A(n2), .B(data_in[6]), .C(n11), .D(data_in[4]), .Z(
        data_out[4]) );
  HS65_LS_AO22X9 U32 ( .A(n2), .B(data_in[8]), .C(n11), .D(data_in[6]), .Z(
        data_out[6]) );
  HS65_LS_AO22X9 U33 ( .A(n2), .B(data_in[10]), .C(n11), .D(data_in[8]), .Z(
        data_out[8]) );
  HS65_LS_AO22X9 U34 ( .A(n2), .B(data_in[12]), .C(n11), .D(data_in[10]), .Z(
        data_out[10]) );
  HS65_LS_AO22X9 U35 ( .A(n2), .B(data_in[14]), .C(n11), .D(data_in[12]), .Z(
        data_out[12]) );
  HS65_LS_AND2X4 U36 ( .A(data_in[14]), .B(n11), .Z(data_out[14]) );
  HS65_LS_CB4I6X9 U37 ( .A(n2), .B(n1), .C(data_valid), .D(preset), .Z(N23) );
  HS65_LS_IVX9 U38 ( .A(data_in_34), .Z(n1) );
endmodule


module latch_controller_1_18 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_18 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_18 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n7) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_IVX9 U3 ( .A(N0), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_0_1_0 ( preset, .chan_in_f({\chan_in_f[REQ] , \chan_in_f[DATA][34] , 
        \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , 
        \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , 
        \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , 
        \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , 
        \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , 
        \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , 
        \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , 
        \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , 
        \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , 
        \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , 
        \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , 
        \chan_in_f[DATA][0] }), .chan_in_b(\chan_in_b[ACK] ), .chan_out_f({
        \chan_out_f[REQ] , \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , 
        \chan_out_f[DATA][32] , \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , 
        \chan_out_f[DATA][29] , \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , 
        \chan_out_f[DATA][26] , \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , 
        \chan_out_f[DATA][23] , \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , 
        \chan_out_f[DATA][20] , \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , 
        \chan_out_f[DATA][17] , \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , 
        \chan_out_f[DATA][14] , \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , 
        \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , 
        \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , 
        \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , 
        \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), 
    .chan_out_b(\chan_out_b[ACK] ), sel );
  output [4:0] sel;
  input preset, \chan_in_f[REQ] , \chan_in_f[DATA][34] , \chan_in_f[DATA][33] ,
         \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , \chan_in_f[DATA][30] ,
         \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , \chan_in_f[DATA][27] ,
         \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , \chan_in_f[DATA][24] ,
         \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , \chan_in_f[DATA][21] ,
         \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , \chan_in_f[DATA][18] ,
         \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , \chan_in_f[DATA][15] ,
         \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , \chan_in_f[DATA][12] ,
         \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , \chan_in_f[DATA][9] ,
         \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , \chan_in_f[DATA][6] ,
         \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , \chan_in_f[DATA][3] ,
         \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , \chan_in_f[DATA][0] ,
         \chan_out_b[ACK] ;
  output \chan_in_b[ACK] , \chan_out_f[REQ] , \chan_out_f[DATA][34] ,
         \chan_out_f[DATA][33] , \chan_out_f[DATA][32] ,
         \chan_out_f[DATA][31] , \chan_out_f[DATA][30] ,
         \chan_out_f[DATA][29] , \chan_out_f[DATA][28] ,
         \chan_out_f[DATA][27] , \chan_out_f[DATA][26] ,
         \chan_out_f[DATA][25] , \chan_out_f[DATA][24] ,
         \chan_out_f[DATA][23] , \chan_out_f[DATA][22] ,
         \chan_out_f[DATA][21] , \chan_out_f[DATA][20] ,
         \chan_out_f[DATA][19] , \chan_out_f[DATA][18] ,
         \chan_out_f[DATA][17] , \chan_out_f[DATA][16] ,
         \chan_out_f[DATA][15] , \chan_out_f[DATA][14] ,
         \chan_out_f[DATA][13] , \chan_out_f[DATA][12] ,
         \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] ,
         \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] ,
         \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] ,
         \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] ;
  wire   \chan_internal_f[REQ] , \chan_internal_f[DATA][34] ,
         \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] ,
         \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] ,
         \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] ,
         \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] ,
         \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] ,
         \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] ,
         \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] ,
         \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] ,
         \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] ,
         \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] ,
         \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] ,
         \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] ,
         \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] ,
         \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] ,
         \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] ,
         \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] ,
         \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] , req_n, lt_en,
         n1, n2, n3, n4, n5, n6, n7;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign sel[1] = 1'b0;

  hpu_comb_0_1_0 hpu_combinatorial ( .data_valid(lt_en), .data_in({
        \chan_in_f[DATA][34] , \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , 
        \chan_in_f[DATA][31] , \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , 
        \chan_in_f[DATA][28] , \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , 
        \chan_in_f[DATA][25] , \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , 
        \chan_in_f[DATA][22] , \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , 
        \chan_in_f[DATA][19] , \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , 
        \chan_in_f[DATA][16] , \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , 
        \chan_in_f[DATA][13] , \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , 
        \chan_in_f[DATA][10] , \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , 
        \chan_in_f[DATA][7] , \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , 
        \chan_in_f[DATA][4] , \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , 
        \chan_in_f[DATA][1] , \chan_in_f[DATA][0] }), .preset(n7), .data_out({
        \chan_internal_f[DATA][34] , \chan_internal_f[DATA][33] , 
        \chan_internal_f[DATA][32] , \chan_internal_f[DATA][31] , 
        \chan_internal_f[DATA][30] , \chan_internal_f[DATA][29] , 
        \chan_internal_f[DATA][28] , \chan_internal_f[DATA][27] , 
        \chan_internal_f[DATA][26] , \chan_internal_f[DATA][25] , 
        \chan_internal_f[DATA][24] , \chan_internal_f[DATA][23] , 
        \chan_internal_f[DATA][22] , \chan_internal_f[DATA][21] , 
        \chan_internal_f[DATA][20] , \chan_internal_f[DATA][19] , 
        \chan_internal_f[DATA][18] , \chan_internal_f[DATA][17] , 
        \chan_internal_f[DATA][16] , \chan_internal_f[DATA][15] , 
        \chan_internal_f[DATA][14] , \chan_internal_f[DATA][13] , 
        \chan_internal_f[DATA][12] , \chan_internal_f[DATA][11] , 
        \chan_internal_f[DATA][10] , \chan_internal_f[DATA][9] , 
        \chan_internal_f[DATA][8] , \chan_internal_f[DATA][7] , 
        \chan_internal_f[DATA][6] , \chan_internal_f[DATA][5] , 
        \chan_internal_f[DATA][4] , \chan_internal_f[DATA][3] , 
        \chan_internal_f[DATA][2] , \chan_internal_f[DATA][1] , 
        \chan_internal_f[DATA][0] }), .sel({sel[4:2], SYNOPSYS_UNCONNECTED__0, 
        sel[0]}) );
  channel_latch_1_xxxxxxxxx_18 token_latch ( .preset(n7), .left_in({
        \chan_internal_f[REQ] , \chan_internal_f[DATA][34] , 
        \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] , 
        \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] , 
        \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] , 
        \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] , 
        \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] , 
        \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] , 
        \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] , 
        \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] , 
        \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] , 
        \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] , 
        \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] , 
        \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] , 
        \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] , 
        \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] , 
        \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] , 
        \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] , 
        \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] }), .left_out(
        \chan_in_b[ACK] ), .right_out({\chan_out_f[REQ] , 
        \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , \chan_out_f[DATA][32] , 
        \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , \chan_out_f[DATA][29] , 
        \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , \chan_out_f[DATA][26] , 
        \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , \chan_out_f[DATA][23] , 
        \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , \chan_out_f[DATA][20] , 
        \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , \chan_out_f[DATA][17] , 
        \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , \chan_out_f[DATA][14] , 
        \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , \chan_out_f[DATA][11] , 
        \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , \chan_out_f[DATA][8] , 
        \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , \chan_out_f[DATA][5] , 
        \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , \chan_out_f[DATA][2] , 
        \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), .right_in(
        \chan_out_b[ACK] ), .lt_enable(lt_en) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chan_internal_f[REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(\chan_in_f[REQ] ), .Z(req_n) );
  HS65_LS_BFX9 U1 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U2 ( .A(n3), .Z(n2) );
  HS65_LS_BFX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_BFX9 U4 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U6 ( .A(req_n), .Z(n6) );
  HS65_LS_BFX9 U7 ( .A(preset), .Z(n7) );
endmodule


module hpu_comb_0_3_0 ( data_valid, data_in, preset, data_out, sel );
  input [34:0] data_in;
  output [34:0] data_out;
  output [4:0] sel;
  input data_valid, preset;
  wire   data_in_34, data_in_33, data_in_32, \data_in[31] , \data_in[30] ,
         \data_in[29] , \data_in[28] , \data_in[27] , \data_in[26] ,
         \data_in[25] , \data_in[24] , \data_in[23] , \data_in[22] ,
         \data_in[21] , \data_in[20] , \data_in[19] , \data_in[18] ,
         \data_in[17] , \data_in[16] , N25, N26, N27, N28, N30, n11, n12, n13,
         n14, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  assign data_out[34] = data_in_34;
  assign data_in_34 = data_in[34];
  assign data_out[33] = data_in_33;
  assign data_in_33 = data_in[33];
  assign data_out[32] = data_in_32;
  assign data_in_32 = data_in[32];
  assign data_out[31] = \data_in[31] ;
  assign \data_in[31]  = data_in[31];
  assign data_out[30] = \data_in[30] ;
  assign \data_in[30]  = data_in[30];
  assign data_out[29] = \data_in[29] ;
  assign \data_in[29]  = data_in[29];
  assign data_out[28] = \data_in[28] ;
  assign \data_in[28]  = data_in[28];
  assign data_out[27] = \data_in[27] ;
  assign \data_in[27]  = data_in[27];
  assign data_out[26] = \data_in[26] ;
  assign \data_in[26]  = data_in[26];
  assign data_out[25] = \data_in[25] ;
  assign \data_in[25]  = data_in[25];
  assign data_out[24] = \data_in[24] ;
  assign \data_in[24]  = data_in[24];
  assign data_out[23] = \data_in[23] ;
  assign \data_in[23]  = data_in[23];
  assign data_out[22] = \data_in[22] ;
  assign \data_in[22]  = data_in[22];
  assign data_out[21] = \data_in[21] ;
  assign \data_in[21]  = data_in[21];
  assign data_out[20] = \data_in[20] ;
  assign \data_in[20]  = data_in[20];
  assign data_out[19] = \data_in[19] ;
  assign \data_in[19]  = data_in[19];
  assign data_out[18] = \data_in[18] ;
  assign \data_in[18]  = data_in[18];
  assign data_out[17] = \data_in[17] ;
  assign \data_in[17]  = data_in[17];
  assign data_out[16] = \data_in[16] ;
  assign \data_in[16]  = data_in[16];
  assign sel[3] = 1'b0;

  HS65_LS_LDHQX9 \sel_reg[4]  ( .G(N25), .D(N30), .Q(sel[4]) );
  HS65_LS_LDHQX9 \sel_reg[2]  ( .G(N25), .D(N28), .Q(sel[2]) );
  HS65_LS_LDHQX9 \sel_reg[1]  ( .G(N25), .D(N27), .Q(sel[1]) );
  HS65_LS_LDHQX9 \sel_reg[0]  ( .G(N25), .D(N26), .Q(sel[0]) );
  HS65_LS_OAI22X6 U4 ( .A(n11), .B(n9), .C(n2), .D(n10), .Z(data_out[0]) );
  HS65_LS_OAI22X6 U5 ( .A(n11), .B(n8), .C(n2), .D(n9), .Z(data_out[2]) );
  HS65_LS_OAI22X6 U6 ( .A(n11), .B(n7), .C(n2), .D(n8), .Z(data_out[4]) );
  HS65_LS_OAI22X6 U7 ( .A(n11), .B(n6), .C(n2), .D(n7), .Z(data_out[6]) );
  HS65_LS_OAI22X6 U8 ( .A(n11), .B(n5), .C(n2), .D(n6), .Z(data_out[8]) );
  HS65_LS_OAI22X6 U9 ( .A(n11), .B(n4), .C(n2), .D(n5), .Z(data_out[10]) );
  HS65_LS_OAI22X6 U10 ( .A(n11), .B(n3), .C(n2), .D(n4), .Z(data_out[12]) );
  HS65_LS_NAND3AX6 U11 ( .A(preset), .B(n12), .C(n2), .Z(n13) );
  HS65_LS_NOR3X4 U12 ( .A(n12), .B(preset), .C(n11), .Z(N30) );
  HS65_LS_IVX9 U13 ( .A(n11), .Z(n2) );
  HS65_LS_NOR2X6 U14 ( .A(n10), .B(n13), .Z(N27) );
  HS65_LS_NOR2AX3 U15 ( .A(n14), .B(n13), .Z(N26) );
  HS65_LS_NOR2X6 U16 ( .A(n2), .B(n3), .Z(data_out[14]) );
  HS65_LS_NAND2X14 U17 ( .A(data_in_34), .B(data_in_33), .Z(n11) );
  HS65_LS_NOR3X4 U18 ( .A(n13), .B(data_in[0]), .C(n14), .Z(N28) );
  HS65_LS_NAND2X7 U19 ( .A(data_in[0]), .B(data_in[1]), .Z(n12) );
  HS65_LS_NOR2X6 U20 ( .A(data_in[1]), .B(data_in[0]), .Z(n14) );
  HS65_LS_IVX9 U21 ( .A(data_in[0]), .Z(n10) );
  HS65_LS_IVX9 U22 ( .A(data_in[2]), .Z(n9) );
  HS65_LS_IVX9 U23 ( .A(data_in[4]), .Z(n8) );
  HS65_LS_IVX9 U24 ( .A(data_in[6]), .Z(n7) );
  HS65_LS_IVX9 U25 ( .A(data_in[8]), .Z(n6) );
  HS65_LS_IVX9 U26 ( .A(data_in[10]), .Z(n5) );
  HS65_LS_IVX9 U27 ( .A(data_in[12]), .Z(n4) );
  HS65_LS_IVX9 U28 ( .A(data_in[14]), .Z(n3) );
  HS65_LS_AO22X9 U29 ( .A(n2), .B(data_in[3]), .C(n11), .D(data_in[1]), .Z(
        data_out[1]) );
  HS65_LS_AO22X9 U30 ( .A(n2), .B(data_in[5]), .C(n11), .D(data_in[3]), .Z(
        data_out[3]) );
  HS65_LS_AO22X9 U31 ( .A(n2), .B(data_in[7]), .C(n11), .D(data_in[5]), .Z(
        data_out[5]) );
  HS65_LS_AO22X9 U32 ( .A(data_in[9]), .B(n2), .C(n11), .D(data_in[7]), .Z(
        data_out[7]) );
  HS65_LS_AO22X9 U33 ( .A(n2), .B(data_in[11]), .C(n11), .D(data_in[9]), .Z(
        data_out[9]) );
  HS65_LS_AO22X9 U34 ( .A(n2), .B(data_in[13]), .C(n11), .D(data_in[11]), .Z(
        data_out[11]) );
  HS65_LS_AO22X9 U35 ( .A(n2), .B(data_in[15]), .C(n11), .D(data_in[13]), .Z(
        data_out[13]) );
  HS65_LS_AND2X4 U36 ( .A(data_in[15]), .B(n11), .Z(data_out[15]) );
  HS65_LS_CB4I6X9 U37 ( .A(n2), .B(n1), .C(data_valid), .D(preset), .Z(N25) );
  HS65_LS_IVX9 U38 ( .A(data_in_34), .Z(n1) );
endmodule


module latch_controller_1_17 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_17 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_17 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n7) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_IVX9 U3 ( .A(N0), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_0_3_0 ( preset, .chan_in_f({\chan_in_f[REQ] , \chan_in_f[DATA][34] , 
        \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , 
        \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , 
        \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , 
        \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , 
        \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , 
        \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , 
        \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , 
        \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , 
        \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , 
        \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , 
        \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , 
        \chan_in_f[DATA][0] }), .chan_in_b(\chan_in_b[ACK] ), .chan_out_f({
        \chan_out_f[REQ] , \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , 
        \chan_out_f[DATA][32] , \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , 
        \chan_out_f[DATA][29] , \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , 
        \chan_out_f[DATA][26] , \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , 
        \chan_out_f[DATA][23] , \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , 
        \chan_out_f[DATA][20] , \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , 
        \chan_out_f[DATA][17] , \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , 
        \chan_out_f[DATA][14] , \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , 
        \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , 
        \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , 
        \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , 
        \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), 
    .chan_out_b(\chan_out_b[ACK] ), sel );
  output [4:0] sel;
  input preset, \chan_in_f[REQ] , \chan_in_f[DATA][34] , \chan_in_f[DATA][33] ,
         \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , \chan_in_f[DATA][30] ,
         \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , \chan_in_f[DATA][27] ,
         \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , \chan_in_f[DATA][24] ,
         \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , \chan_in_f[DATA][21] ,
         \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , \chan_in_f[DATA][18] ,
         \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , \chan_in_f[DATA][15] ,
         \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , \chan_in_f[DATA][12] ,
         \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , \chan_in_f[DATA][9] ,
         \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , \chan_in_f[DATA][6] ,
         \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , \chan_in_f[DATA][3] ,
         \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , \chan_in_f[DATA][0] ,
         \chan_out_b[ACK] ;
  output \chan_in_b[ACK] , \chan_out_f[REQ] , \chan_out_f[DATA][34] ,
         \chan_out_f[DATA][33] , \chan_out_f[DATA][32] ,
         \chan_out_f[DATA][31] , \chan_out_f[DATA][30] ,
         \chan_out_f[DATA][29] , \chan_out_f[DATA][28] ,
         \chan_out_f[DATA][27] , \chan_out_f[DATA][26] ,
         \chan_out_f[DATA][25] , \chan_out_f[DATA][24] ,
         \chan_out_f[DATA][23] , \chan_out_f[DATA][22] ,
         \chan_out_f[DATA][21] , \chan_out_f[DATA][20] ,
         \chan_out_f[DATA][19] , \chan_out_f[DATA][18] ,
         \chan_out_f[DATA][17] , \chan_out_f[DATA][16] ,
         \chan_out_f[DATA][15] , \chan_out_f[DATA][14] ,
         \chan_out_f[DATA][13] , \chan_out_f[DATA][12] ,
         \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] ,
         \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] ,
         \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] ,
         \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] ;
  wire   \chan_internal_f[REQ] , \chan_internal_f[DATA][34] ,
         \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] ,
         \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] ,
         \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] ,
         \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] ,
         \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] ,
         \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] ,
         \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] ,
         \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] ,
         \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] ,
         \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] ,
         \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] ,
         \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] ,
         \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] ,
         \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] ,
         \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] ,
         \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] ,
         \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] , req_n, lt_en,
         n1, n2, n3, n4, n5, n6, n7;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign sel[3] = 1'b0;

  hpu_comb_0_3_0 hpu_combinatorial ( .data_valid(lt_en), .data_in({
        \chan_in_f[DATA][34] , \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , 
        \chan_in_f[DATA][31] , \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , 
        \chan_in_f[DATA][28] , \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , 
        \chan_in_f[DATA][25] , \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , 
        \chan_in_f[DATA][22] , \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , 
        \chan_in_f[DATA][19] , \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , 
        \chan_in_f[DATA][16] , \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , 
        \chan_in_f[DATA][13] , \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , 
        \chan_in_f[DATA][10] , \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , 
        \chan_in_f[DATA][7] , \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , 
        \chan_in_f[DATA][4] , \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , 
        \chan_in_f[DATA][1] , \chan_in_f[DATA][0] }), .preset(n7), .data_out({
        \chan_internal_f[DATA][34] , \chan_internal_f[DATA][33] , 
        \chan_internal_f[DATA][32] , \chan_internal_f[DATA][31] , 
        \chan_internal_f[DATA][30] , \chan_internal_f[DATA][29] , 
        \chan_internal_f[DATA][28] , \chan_internal_f[DATA][27] , 
        \chan_internal_f[DATA][26] , \chan_internal_f[DATA][25] , 
        \chan_internal_f[DATA][24] , \chan_internal_f[DATA][23] , 
        \chan_internal_f[DATA][22] , \chan_internal_f[DATA][21] , 
        \chan_internal_f[DATA][20] , \chan_internal_f[DATA][19] , 
        \chan_internal_f[DATA][18] , \chan_internal_f[DATA][17] , 
        \chan_internal_f[DATA][16] , \chan_internal_f[DATA][15] , 
        \chan_internal_f[DATA][14] , \chan_internal_f[DATA][13] , 
        \chan_internal_f[DATA][12] , \chan_internal_f[DATA][11] , 
        \chan_internal_f[DATA][10] , \chan_internal_f[DATA][9] , 
        \chan_internal_f[DATA][8] , \chan_internal_f[DATA][7] , 
        \chan_internal_f[DATA][6] , \chan_internal_f[DATA][5] , 
        \chan_internal_f[DATA][4] , \chan_internal_f[DATA][3] , 
        \chan_internal_f[DATA][2] , \chan_internal_f[DATA][1] , 
        \chan_internal_f[DATA][0] }), .sel({sel[4], SYNOPSYS_UNCONNECTED__0, 
        sel[2:0]}) );
  channel_latch_1_xxxxxxxxx_17 token_latch ( .preset(n7), .left_in({
        \chan_internal_f[REQ] , \chan_internal_f[DATA][34] , 
        \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] , 
        \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] , 
        \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] , 
        \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] , 
        \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] , 
        \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] , 
        \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] , 
        \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] , 
        \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] , 
        \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] , 
        \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] , 
        \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] , 
        \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] , 
        \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] , 
        \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] , 
        \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] , 
        \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] }), .left_out(
        \chan_in_b[ACK] ), .right_out({\chan_out_f[REQ] , 
        \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , \chan_out_f[DATA][32] , 
        \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , \chan_out_f[DATA][29] , 
        \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , \chan_out_f[DATA][26] , 
        \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , \chan_out_f[DATA][23] , 
        \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , \chan_out_f[DATA][20] , 
        \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , \chan_out_f[DATA][17] , 
        \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , \chan_out_f[DATA][14] , 
        \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , \chan_out_f[DATA][11] , 
        \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , \chan_out_f[DATA][8] , 
        \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , \chan_out_f[DATA][5] , 
        \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , \chan_out_f[DATA][2] , 
        \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), .right_in(
        \chan_out_b[ACK] ), .lt_enable(lt_en) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chan_internal_f[REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(\chan_in_f[REQ] ), .Z(req_n) );
  HS65_LS_BFX9 U1 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U2 ( .A(n3), .Z(n2) );
  HS65_LS_BFX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_BFX9 U4 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U6 ( .A(req_n), .Z(n6) );
  HS65_LS_BFX9 U7 ( .A(preset), .Z(n7) );
endmodule


module hpu_comb_1_x_0 ( data_valid, data_in, preset, data_out, sel );
  input [34:0] data_in;
  output [34:0] data_out;
  output [4:0] sel;
  input data_valid, preset;
  wire   data_in_34, data_in_33, data_in_32, \data_in[31] , \data_in[30] ,
         \data_in[29] , \data_in[28] , \data_in[27] , \data_in[26] ,
         \data_in[25] , \data_in[24] , \data_in[23] , \data_in[22] ,
         \data_in[21] , \data_in[20] , \data_in[19] , \data_in[18] ,
         \data_in[17] , \data_in[16] , N19, N20, N21, N22, N23, n19, n20, n21,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;
  assign data_out[34] = data_in_34;
  assign data_in_34 = data_in[34];
  assign data_out[33] = data_in_33;
  assign data_in_33 = data_in[33];
  assign data_out[32] = data_in_32;
  assign data_in_32 = data_in[32];
  assign data_out[31] = \data_in[31] ;
  assign \data_in[31]  = data_in[31];
  assign data_out[30] = \data_in[30] ;
  assign \data_in[30]  = data_in[30];
  assign data_out[29] = \data_in[29] ;
  assign \data_in[29]  = data_in[29];
  assign data_out[28] = \data_in[28] ;
  assign \data_in[28]  = data_in[28];
  assign data_out[27] = \data_in[27] ;
  assign \data_in[27]  = data_in[27];
  assign data_out[26] = \data_in[26] ;
  assign \data_in[26]  = data_in[26];
  assign data_out[25] = \data_in[25] ;
  assign \data_in[25]  = data_in[25];
  assign data_out[24] = \data_in[24] ;
  assign \data_in[24]  = data_in[24];
  assign data_out[23] = \data_in[23] ;
  assign \data_in[23]  = data_in[23];
  assign data_out[22] = \data_in[22] ;
  assign \data_in[22]  = data_in[22];
  assign data_out[21] = \data_in[21] ;
  assign \data_in[21]  = data_in[21];
  assign data_out[20] = \data_in[20] ;
  assign \data_in[20]  = data_in[20];
  assign data_out[19] = \data_in[19] ;
  assign \data_in[19]  = data_in[19];
  assign data_out[18] = \data_in[18] ;
  assign \data_in[18]  = data_in[18];
  assign data_out[17] = \data_in[17] ;
  assign \data_in[17]  = data_in[17];
  assign data_out[16] = \data_in[16] ;
  assign \data_in[16]  = data_in[16];
  assign sel[4] = 1'b0;

  HS65_LS_LDHQX9 \sel_reg[3]  ( .G(N19), .D(N23), .Q(sel[3]) );
  HS65_LS_LDHQX9 \sel_reg[2]  ( .G(N19), .D(N22), .Q(sel[2]) );
  HS65_LS_LDHQX9 \sel_reg[1]  ( .G(N19), .D(N21), .Q(sel[1]) );
  HS65_LS_LDHQX9 \sel_reg[0]  ( .G(N19), .D(N20), .Q(sel[0]) );
  HS65_LS_NAND2X21 U4 ( .A(data_in_34), .B(data_in_33), .Z(n19) );
  HS65_LS_NAND3AX6 U5 ( .A(preset), .B(n21), .C(n2), .Z(n20) );
  HS65_LS_OAI22X6 U6 ( .A(n9), .B(n19), .C(n2), .D(n11), .Z(data_out[7]) );
  HS65_LS_OAI22X6 U7 ( .A(n19), .B(n16), .C(n2), .D(n18), .Z(data_out[0]) );
  HS65_LS_OAI22X6 U8 ( .A(n19), .B(n15), .C(n2), .D(n17), .Z(data_out[1]) );
  HS65_LS_OAI22X6 U9 ( .A(n19), .B(n14), .C(n2), .D(n16), .Z(data_out[2]) );
  HS65_LS_OAI22X6 U10 ( .A(n19), .B(n13), .C(n2), .D(n15), .Z(data_out[3]) );
  HS65_LS_OAI22X6 U11 ( .A(n19), .B(n12), .C(n2), .D(n14), .Z(data_out[4]) );
  HS65_LS_OAI22X6 U12 ( .A(n19), .B(n11), .C(n2), .D(n13), .Z(data_out[5]) );
  HS65_LS_OAI22X6 U13 ( .A(n19), .B(n10), .C(n2), .D(n12), .Z(data_out[6]) );
  HS65_LS_OAI22X6 U14 ( .A(n19), .B(n8), .C(n2), .D(n10), .Z(data_out[8]) );
  HS65_LS_OAI22X6 U15 ( .A(n19), .B(n7), .C(n2), .D(n9), .Z(data_out[9]) );
  HS65_LS_OAI22X6 U16 ( .A(n19), .B(n6), .C(n2), .D(n8), .Z(data_out[10]) );
  HS65_LS_OAI22X6 U17 ( .A(n19), .B(n5), .C(n2), .D(n7), .Z(data_out[11]) );
  HS65_LS_OAI22X6 U18 ( .A(n19), .B(n4), .C(n2), .D(n6), .Z(data_out[12]) );
  HS65_LS_OAI22X6 U19 ( .A(n19), .B(n3), .C(n2), .D(n5), .Z(data_out[13]) );
  HS65_LS_IVX9 U20 ( .A(n19), .Z(n2) );
  HS65_LS_NOR3X4 U21 ( .A(n21), .B(preset), .C(n19), .Z(N20) );
  HS65_LS_NOR3X4 U22 ( .A(n20), .B(n17), .C(n18), .Z(N23) );
  HS65_LS_NAND2X7 U23 ( .A(n17), .B(n18), .Z(n21) );
  HS65_LS_NOR2X6 U24 ( .A(n2), .B(n4), .Z(data_out[14]) );
  HS65_LS_NOR2X6 U25 ( .A(n2), .B(n3), .Z(data_out[15]) );
  HS65_LS_IVX9 U26 ( .A(data_in[1]), .Z(n17) );
  HS65_LS_IVX9 U27 ( .A(data_in[0]), .Z(n18) );
  HS65_LS_NOR2X6 U28 ( .A(data_in[1]), .B(n20), .Z(N21) );
  HS65_LS_NOR2X6 U29 ( .A(data_in[0]), .B(n20), .Z(N22) );
  HS65_LS_IVX9 U30 ( .A(data_in[9]), .Z(n9) );
  HS65_LS_IVX9 U31 ( .A(data_in[2]), .Z(n16) );
  HS65_LS_IVX9 U32 ( .A(data_in[3]), .Z(n15) );
  HS65_LS_IVX9 U33 ( .A(data_in[4]), .Z(n14) );
  HS65_LS_IVX9 U34 ( .A(data_in[5]), .Z(n13) );
  HS65_LS_IVX9 U35 ( .A(data_in[7]), .Z(n11) );
  HS65_LS_IVX9 U36 ( .A(data_in[10]), .Z(n8) );
  HS65_LS_IVX9 U37 ( .A(data_in[12]), .Z(n6) );
  HS65_LS_IVX9 U38 ( .A(data_in[13]), .Z(n5) );
  HS65_LS_IVX9 U39 ( .A(data_in[14]), .Z(n4) );
  HS65_LS_IVX9 U40 ( .A(data_in[15]), .Z(n3) );
  HS65_LS_IVX9 U41 ( .A(data_in[6]), .Z(n12) );
  HS65_LS_IVX9 U42 ( .A(data_in[8]), .Z(n10) );
  HS65_LS_IVX9 U43 ( .A(data_in[11]), .Z(n7) );
  HS65_LS_CB4I6X9 U44 ( .A(n2), .B(n1), .C(data_valid), .D(preset), .Z(N19) );
  HS65_LS_IVX9 U45 ( .A(data_in_34), .Z(n1) );
endmodule


module latch_controller_1_16 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_16 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_16 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n7) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_IVX9 U3 ( .A(N0), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_1_x_0 ( preset, .chan_in_f({\chan_in_f[REQ] , \chan_in_f[DATA][34] , 
        \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , 
        \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , 
        \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , 
        \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , 
        \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , 
        \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , 
        \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , 
        \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , 
        \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , 
        \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , 
        \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , 
        \chan_in_f[DATA][0] }), .chan_in_b(\chan_in_b[ACK] ), .chan_out_f({
        \chan_out_f[REQ] , \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , 
        \chan_out_f[DATA][32] , \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , 
        \chan_out_f[DATA][29] , \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , 
        \chan_out_f[DATA][26] , \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , 
        \chan_out_f[DATA][23] , \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , 
        \chan_out_f[DATA][20] , \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , 
        \chan_out_f[DATA][17] , \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , 
        \chan_out_f[DATA][14] , \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , 
        \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , 
        \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , 
        \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , 
        \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), 
    .chan_out_b(\chan_out_b[ACK] ), sel );
  output [4:0] sel;
  input preset, \chan_in_f[REQ] , \chan_in_f[DATA][34] , \chan_in_f[DATA][33] ,
         \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , \chan_in_f[DATA][30] ,
         \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , \chan_in_f[DATA][27] ,
         \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , \chan_in_f[DATA][24] ,
         \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , \chan_in_f[DATA][21] ,
         \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , \chan_in_f[DATA][18] ,
         \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , \chan_in_f[DATA][15] ,
         \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , \chan_in_f[DATA][12] ,
         \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , \chan_in_f[DATA][9] ,
         \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , \chan_in_f[DATA][6] ,
         \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , \chan_in_f[DATA][3] ,
         \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , \chan_in_f[DATA][0] ,
         \chan_out_b[ACK] ;
  output \chan_in_b[ACK] , \chan_out_f[REQ] , \chan_out_f[DATA][34] ,
         \chan_out_f[DATA][33] , \chan_out_f[DATA][32] ,
         \chan_out_f[DATA][31] , \chan_out_f[DATA][30] ,
         \chan_out_f[DATA][29] , \chan_out_f[DATA][28] ,
         \chan_out_f[DATA][27] , \chan_out_f[DATA][26] ,
         \chan_out_f[DATA][25] , \chan_out_f[DATA][24] ,
         \chan_out_f[DATA][23] , \chan_out_f[DATA][22] ,
         \chan_out_f[DATA][21] , \chan_out_f[DATA][20] ,
         \chan_out_f[DATA][19] , \chan_out_f[DATA][18] ,
         \chan_out_f[DATA][17] , \chan_out_f[DATA][16] ,
         \chan_out_f[DATA][15] , \chan_out_f[DATA][14] ,
         \chan_out_f[DATA][13] , \chan_out_f[DATA][12] ,
         \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] ,
         \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] ,
         \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] ,
         \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] ;
  wire   \chan_internal_f[REQ] , \chan_internal_f[DATA][34] ,
         \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] ,
         \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] ,
         \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] ,
         \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] ,
         \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] ,
         \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] ,
         \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] ,
         \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] ,
         \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] ,
         \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] ,
         \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] ,
         \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] ,
         \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] ,
         \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] ,
         \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] ,
         \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] ,
         \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] , req_n, lt_en,
         n1, n2, n3, n4, n5, n6, n7;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign sel[4] = 1'b0;

  hpu_comb_1_x_0 hpu_combinatorial ( .data_valid(lt_en), .data_in({
        \chan_in_f[DATA][34] , \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , 
        \chan_in_f[DATA][31] , \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , 
        \chan_in_f[DATA][28] , \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , 
        \chan_in_f[DATA][25] , \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , 
        \chan_in_f[DATA][22] , \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , 
        \chan_in_f[DATA][19] , \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , 
        \chan_in_f[DATA][16] , \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , 
        \chan_in_f[DATA][13] , \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , 
        \chan_in_f[DATA][10] , \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , 
        \chan_in_f[DATA][7] , \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , 
        \chan_in_f[DATA][4] , \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , 
        \chan_in_f[DATA][1] , \chan_in_f[DATA][0] }), .preset(n7), .data_out({
        \chan_internal_f[DATA][34] , \chan_internal_f[DATA][33] , 
        \chan_internal_f[DATA][32] , \chan_internal_f[DATA][31] , 
        \chan_internal_f[DATA][30] , \chan_internal_f[DATA][29] , 
        \chan_internal_f[DATA][28] , \chan_internal_f[DATA][27] , 
        \chan_internal_f[DATA][26] , \chan_internal_f[DATA][25] , 
        \chan_internal_f[DATA][24] , \chan_internal_f[DATA][23] , 
        \chan_internal_f[DATA][22] , \chan_internal_f[DATA][21] , 
        \chan_internal_f[DATA][20] , \chan_internal_f[DATA][19] , 
        \chan_internal_f[DATA][18] , \chan_internal_f[DATA][17] , 
        \chan_internal_f[DATA][16] , \chan_internal_f[DATA][15] , 
        \chan_internal_f[DATA][14] , \chan_internal_f[DATA][13] , 
        \chan_internal_f[DATA][12] , \chan_internal_f[DATA][11] , 
        \chan_internal_f[DATA][10] , \chan_internal_f[DATA][9] , 
        \chan_internal_f[DATA][8] , \chan_internal_f[DATA][7] , 
        \chan_internal_f[DATA][6] , \chan_internal_f[DATA][5] , 
        \chan_internal_f[DATA][4] , \chan_internal_f[DATA][3] , 
        \chan_internal_f[DATA][2] , \chan_internal_f[DATA][1] , 
        \chan_internal_f[DATA][0] }), .sel({SYNOPSYS_UNCONNECTED__0, sel[3:0]}) );
  channel_latch_1_xxxxxxxxx_16 token_latch ( .preset(n7), .left_in({
        \chan_internal_f[REQ] , \chan_internal_f[DATA][34] , 
        \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] , 
        \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] , 
        \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] , 
        \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] , 
        \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] , 
        \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] , 
        \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] , 
        \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] , 
        \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] , 
        \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] , 
        \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] , 
        \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] , 
        \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] , 
        \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] , 
        \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] , 
        \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] , 
        \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] }), .left_out(
        \chan_in_b[ACK] ), .right_out({\chan_out_f[REQ] , 
        \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , \chan_out_f[DATA][32] , 
        \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , \chan_out_f[DATA][29] , 
        \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , \chan_out_f[DATA][26] , 
        \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , \chan_out_f[DATA][23] , 
        \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , \chan_out_f[DATA][20] , 
        \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , \chan_out_f[DATA][17] , 
        \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , \chan_out_f[DATA][14] , 
        \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , \chan_out_f[DATA][11] , 
        \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , \chan_out_f[DATA][8] , 
        \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , \chan_out_f[DATA][5] , 
        \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , \chan_out_f[DATA][2] , 
        \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), .right_in(
        \chan_out_b[ACK] ), .lt_enable(lt_en) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chan_internal_f[REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(\chan_in_f[REQ] ), .Z(req_n) );
  HS65_LS_BFX9 U1 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U2 ( .A(n3), .Z(n2) );
  HS65_LS_BFX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_BFX9 U4 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U6 ( .A(req_n), .Z(n6) );
  HS65_LS_BFX9 U7 ( .A(preset), .Z(n7) );
endmodule


module sr_latch_1_0 ( s, r, q, qn );
  input s, r;
  output q, qn;
  wire   N3, n1;

  HS65_LS_AND2X4 C9 ( .A(n1), .B(N3), .Z(qn) );
  HS65_LH_NOR2X3 U1 ( .A(r), .B(qn), .Z(q) );
  HS65_LS_IVX9 U2 ( .A(q), .Z(N3) );
  HS65_LS_IVX9 U3 ( .A(s), .Z(n1) );
endmodule


module c_gate_generic_1_5_0 ( preset, \input , \output  );
  input [4:0] \input ;
  input preset;
  output \output ;
  wire   set, reset, n2, n3, n1;

  sr_latch_1_0 latch ( .s(set), .r(reset), .q(\output ) );
  HS65_LS_NOR3X4 U3 ( .A(\input [3]), .B(preset), .C(\input [4]), .Z(n3) );
  HS65_LS_NOR4ABX2 U4 ( .A(n1), .B(n3), .C(\input [2]), .D(\input [1]), .Z(
        reset) );
  HS65_LS_AO31X9 U5 ( .A(n2), .B(\input [3]), .C(\input [4]), .D(preset), .Z(
        set) );
  HS65_LS_IVX9 U6 ( .A(\input [0]), .Z(n1) );
  HS65_LS_AND3X9 U7 ( .A(\input [1]), .B(\input [0]), .C(\input [2]), .Z(n2)
         );
endmodule


module sr_latch_1_7 ( s, r, q, qn );
  input s, r;
  output q, qn;
  wire   N3, n1;

  HS65_LS_AND2X4 C9 ( .A(n1), .B(N3), .Z(qn) );
  HS65_LS_IVX9 U1 ( .A(q), .Z(N3) );
  HS65_LS_IVX9 U2 ( .A(s), .Z(n1) );
  HS65_LS_NOR2X6 U3 ( .A(r), .B(qn), .Z(q) );
endmodule


module c_gate_generic_1_5_7 ( preset, \input , \output  );
  input [4:0] \input ;
  input preset;
  output \output ;
  wire   set, reset, n1, n4, n5;

  sr_latch_1_7 latch ( .s(set), .r(reset), .q(\output ) );
  HS65_LS_NOR3X4 U3 ( .A(\input [3]), .B(preset), .C(\input [4]), .Z(n4) );
  HS65_LS_NOR4ABX2 U4 ( .A(n1), .B(n4), .C(\input [2]), .D(\input [1]), .Z(
        reset) );
  HS65_LS_AO31X9 U5 ( .A(n5), .B(\input [3]), .C(\input [4]), .D(preset), .Z(
        set) );
  HS65_LS_IVX9 U6 ( .A(\input [0]), .Z(n1) );
  HS65_LS_AND3X9 U7 ( .A(\input [1]), .B(\input [0]), .C(\input [2]), .Z(n5)
         );
endmodule


module crossbar_0 ( preset, .switch_sel({\switch_sel[4][4] , 
        \switch_sel[4][3] , \switch_sel[4][2] , \switch_sel[4][1] , 
        \switch_sel[4][0] , \switch_sel[3][4] , \switch_sel[3][3] , 
        \switch_sel[3][2] , \switch_sel[3][1] , \switch_sel[3][0] , 
        \switch_sel[2][4] , \switch_sel[2][3] , \switch_sel[2][2] , 
        \switch_sel[2][1] , \switch_sel[2][0] , \switch_sel[1][4] , 
        \switch_sel[1][3] , \switch_sel[1][2] , \switch_sel[1][1] , 
        \switch_sel[1][0] , \switch_sel[0][4] , \switch_sel[0][3] , 
        \switch_sel[0][2] , \switch_sel[0][1] , \switch_sel[0][0] }), 
    .chs_in_f({\chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] , 
        \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] , 
        \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] , 
        \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] , 
        \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] , 
        \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] , 
        \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] , 
        \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] , 
        \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] , 
        \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] , 
        \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] , 
        \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] , 
        \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] , 
        \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] , \chs_in_f[4][DATA][7] , 
        \chs_in_f[4][DATA][6] , \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] , 
        \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] , \chs_in_f[4][DATA][1] , 
        \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] , \chs_in_f[3][DATA][34] , 
        \chs_in_f[3][DATA][33] , \chs_in_f[3][DATA][32] , 
        \chs_in_f[3][DATA][31] , \chs_in_f[3][DATA][30] , 
        \chs_in_f[3][DATA][29] , \chs_in_f[3][DATA][28] , 
        \chs_in_f[3][DATA][27] , \chs_in_f[3][DATA][26] , 
        \chs_in_f[3][DATA][25] , \chs_in_f[3][DATA][24] , 
        \chs_in_f[3][DATA][23] , \chs_in_f[3][DATA][22] , 
        \chs_in_f[3][DATA][21] , \chs_in_f[3][DATA][20] , 
        \chs_in_f[3][DATA][19] , \chs_in_f[3][DATA][18] , 
        \chs_in_f[3][DATA][17] , \chs_in_f[3][DATA][16] , 
        \chs_in_f[3][DATA][15] , \chs_in_f[3][DATA][14] , 
        \chs_in_f[3][DATA][13] , \chs_in_f[3][DATA][12] , 
        \chs_in_f[3][DATA][11] , \chs_in_f[3][DATA][10] , 
        \chs_in_f[3][DATA][9] , \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] , 
        \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] , \chs_in_f[3][DATA][4] , 
        \chs_in_f[3][DATA][3] , \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] , 
        \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] , 
        \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] , 
        \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] , 
        \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] , 
        \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] , 
        \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] , 
        \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] , 
        \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] , 
        \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] , 
        \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] , 
        \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] , 
        \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] , 
        \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] , 
        \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] , \chs_in_f[2][DATA][7] , 
        \chs_in_f[2][DATA][6] , \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] , 
        \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] , \chs_in_f[2][DATA][1] , 
        \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] , \chs_in_f[1][DATA][34] , 
        \chs_in_f[1][DATA][33] , \chs_in_f[1][DATA][32] , 
        \chs_in_f[1][DATA][31] , \chs_in_f[1][DATA][30] , 
        \chs_in_f[1][DATA][29] , \chs_in_f[1][DATA][28] , 
        \chs_in_f[1][DATA][27] , \chs_in_f[1][DATA][26] , 
        \chs_in_f[1][DATA][25] , \chs_in_f[1][DATA][24] , 
        \chs_in_f[1][DATA][23] , \chs_in_f[1][DATA][22] , 
        \chs_in_f[1][DATA][21] , \chs_in_f[1][DATA][20] , 
        \chs_in_f[1][DATA][19] , \chs_in_f[1][DATA][18] , 
        \chs_in_f[1][DATA][17] , \chs_in_f[1][DATA][16] , 
        \chs_in_f[1][DATA][15] , \chs_in_f[1][DATA][14] , 
        \chs_in_f[1][DATA][13] , \chs_in_f[1][DATA][12] , 
        \chs_in_f[1][DATA][11] , \chs_in_f[1][DATA][10] , 
        \chs_in_f[1][DATA][9] , \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] , 
        \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] , \chs_in_f[1][DATA][4] , 
        \chs_in_f[1][DATA][3] , \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] , 
        \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] , 
        \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] , 
        \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] , 
        \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] , 
        \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] , 
        \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] , 
        \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] , 
        \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] , 
        \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] , 
        \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] , 
        \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] , 
        \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] , 
        \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] , 
        \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] , \chs_in_f[0][DATA][7] , 
        \chs_in_f[0][DATA][6] , \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] , 
        \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] , \chs_in_f[0][DATA][1] , 
        \chs_in_f[0][DATA][0] }), .chs_in_b({\chs_in_b[4][ACK] , 
        \chs_in_b[3][ACK] , \chs_in_b[2][ACK] , \chs_in_b[1][ACK] , 
        \chs_in_b[0][ACK] }), .chs_out_f({\chs_out_f[4][REQ] , 
        \chs_out_f[4][DATA][34] , \chs_out_f[4][DATA][33] , 
        \chs_out_f[4][DATA][32] , \chs_out_f[4][DATA][31] , 
        \chs_out_f[4][DATA][30] , \chs_out_f[4][DATA][29] , 
        \chs_out_f[4][DATA][28] , \chs_out_f[4][DATA][27] , 
        \chs_out_f[4][DATA][26] , \chs_out_f[4][DATA][25] , 
        \chs_out_f[4][DATA][24] , \chs_out_f[4][DATA][23] , 
        \chs_out_f[4][DATA][22] , \chs_out_f[4][DATA][21] , 
        \chs_out_f[4][DATA][20] , \chs_out_f[4][DATA][19] , 
        \chs_out_f[4][DATA][18] , \chs_out_f[4][DATA][17] , 
        \chs_out_f[4][DATA][16] , \chs_out_f[4][DATA][15] , 
        \chs_out_f[4][DATA][14] , \chs_out_f[4][DATA][13] , 
        \chs_out_f[4][DATA][12] , \chs_out_f[4][DATA][11] , 
        \chs_out_f[4][DATA][10] , \chs_out_f[4][DATA][9] , 
        \chs_out_f[4][DATA][8] , \chs_out_f[4][DATA][7] , 
        \chs_out_f[4][DATA][6] , \chs_out_f[4][DATA][5] , 
        \chs_out_f[4][DATA][4] , \chs_out_f[4][DATA][3] , 
        \chs_out_f[4][DATA][2] , \chs_out_f[4][DATA][1] , 
        \chs_out_f[4][DATA][0] , \chs_out_f[3][REQ] , \chs_out_f[3][DATA][34] , 
        \chs_out_f[3][DATA][33] , \chs_out_f[3][DATA][32] , 
        \chs_out_f[3][DATA][31] , \chs_out_f[3][DATA][30] , 
        \chs_out_f[3][DATA][29] , \chs_out_f[3][DATA][28] , 
        \chs_out_f[3][DATA][27] , \chs_out_f[3][DATA][26] , 
        \chs_out_f[3][DATA][25] , \chs_out_f[3][DATA][24] , 
        \chs_out_f[3][DATA][23] , \chs_out_f[3][DATA][22] , 
        \chs_out_f[3][DATA][21] , \chs_out_f[3][DATA][20] , 
        \chs_out_f[3][DATA][19] , \chs_out_f[3][DATA][18] , 
        \chs_out_f[3][DATA][17] , \chs_out_f[3][DATA][16] , 
        \chs_out_f[3][DATA][15] , \chs_out_f[3][DATA][14] , 
        \chs_out_f[3][DATA][13] , \chs_out_f[3][DATA][12] , 
        \chs_out_f[3][DATA][11] , \chs_out_f[3][DATA][10] , 
        \chs_out_f[3][DATA][9] , \chs_out_f[3][DATA][8] , 
        \chs_out_f[3][DATA][7] , \chs_out_f[3][DATA][6] , 
        \chs_out_f[3][DATA][5] , \chs_out_f[3][DATA][4] , 
        \chs_out_f[3][DATA][3] , \chs_out_f[3][DATA][2] , 
        \chs_out_f[3][DATA][1] , \chs_out_f[3][DATA][0] , \chs_out_f[2][REQ] , 
        \chs_out_f[2][DATA][34] , \chs_out_f[2][DATA][33] , 
        \chs_out_f[2][DATA][32] , \chs_out_f[2][DATA][31] , 
        \chs_out_f[2][DATA][30] , \chs_out_f[2][DATA][29] , 
        \chs_out_f[2][DATA][28] , \chs_out_f[2][DATA][27] , 
        \chs_out_f[2][DATA][26] , \chs_out_f[2][DATA][25] , 
        \chs_out_f[2][DATA][24] , \chs_out_f[2][DATA][23] , 
        \chs_out_f[2][DATA][22] , \chs_out_f[2][DATA][21] , 
        \chs_out_f[2][DATA][20] , \chs_out_f[2][DATA][19] , 
        \chs_out_f[2][DATA][18] , \chs_out_f[2][DATA][17] , 
        \chs_out_f[2][DATA][16] , \chs_out_f[2][DATA][15] , 
        \chs_out_f[2][DATA][14] , \chs_out_f[2][DATA][13] , 
        \chs_out_f[2][DATA][12] , \chs_out_f[2][DATA][11] , 
        \chs_out_f[2][DATA][10] , \chs_out_f[2][DATA][9] , 
        \chs_out_f[2][DATA][8] , \chs_out_f[2][DATA][7] , 
        \chs_out_f[2][DATA][6] , \chs_out_f[2][DATA][5] , 
        \chs_out_f[2][DATA][4] , \chs_out_f[2][DATA][3] , 
        \chs_out_f[2][DATA][2] , \chs_out_f[2][DATA][1] , 
        \chs_out_f[2][DATA][0] , \chs_out_f[1][REQ] , \chs_out_f[1][DATA][34] , 
        \chs_out_f[1][DATA][33] , \chs_out_f[1][DATA][32] , 
        \chs_out_f[1][DATA][31] , \chs_out_f[1][DATA][30] , 
        \chs_out_f[1][DATA][29] , \chs_out_f[1][DATA][28] , 
        \chs_out_f[1][DATA][27] , \chs_out_f[1][DATA][26] , 
        \chs_out_f[1][DATA][25] , \chs_out_f[1][DATA][24] , 
        \chs_out_f[1][DATA][23] , \chs_out_f[1][DATA][22] , 
        \chs_out_f[1][DATA][21] , \chs_out_f[1][DATA][20] , 
        \chs_out_f[1][DATA][19] , \chs_out_f[1][DATA][18] , 
        \chs_out_f[1][DATA][17] , \chs_out_f[1][DATA][16] , 
        \chs_out_f[1][DATA][15] , \chs_out_f[1][DATA][14] , 
        \chs_out_f[1][DATA][13] , \chs_out_f[1][DATA][12] , 
        \chs_out_f[1][DATA][11] , \chs_out_f[1][DATA][10] , 
        \chs_out_f[1][DATA][9] , \chs_out_f[1][DATA][8] , 
        \chs_out_f[1][DATA][7] , \chs_out_f[1][DATA][6] , 
        \chs_out_f[1][DATA][5] , \chs_out_f[1][DATA][4] , 
        \chs_out_f[1][DATA][3] , \chs_out_f[1][DATA][2] , 
        \chs_out_f[1][DATA][1] , \chs_out_f[1][DATA][0] , \chs_out_f[0][REQ] , 
        \chs_out_f[0][DATA][34] , \chs_out_f[0][DATA][33] , 
        \chs_out_f[0][DATA][32] , \chs_out_f[0][DATA][31] , 
        \chs_out_f[0][DATA][30] , \chs_out_f[0][DATA][29] , 
        \chs_out_f[0][DATA][28] , \chs_out_f[0][DATA][27] , 
        \chs_out_f[0][DATA][26] , \chs_out_f[0][DATA][25] , 
        \chs_out_f[0][DATA][24] , \chs_out_f[0][DATA][23] , 
        \chs_out_f[0][DATA][22] , \chs_out_f[0][DATA][21] , 
        \chs_out_f[0][DATA][20] , \chs_out_f[0][DATA][19] , 
        \chs_out_f[0][DATA][18] , \chs_out_f[0][DATA][17] , 
        \chs_out_f[0][DATA][16] , \chs_out_f[0][DATA][15] , 
        \chs_out_f[0][DATA][14] , \chs_out_f[0][DATA][13] , 
        \chs_out_f[0][DATA][12] , \chs_out_f[0][DATA][11] , 
        \chs_out_f[0][DATA][10] , \chs_out_f[0][DATA][9] , 
        \chs_out_f[0][DATA][8] , \chs_out_f[0][DATA][7] , 
        \chs_out_f[0][DATA][6] , \chs_out_f[0][DATA][5] , 
        \chs_out_f[0][DATA][4] , \chs_out_f[0][DATA][3] , 
        \chs_out_f[0][DATA][2] , \chs_out_f[0][DATA][1] , 
        \chs_out_f[0][DATA][0] }), .chs_out_b({\chs_out_b[4][ACK] , 
        \chs_out_b[3][ACK] , \chs_out_b[2][ACK] , \chs_out_b[1][ACK] , 
        \chs_out_b[0][ACK] }) );
  input preset, \switch_sel[4][4] , \switch_sel[4][3] , \switch_sel[4][2] ,
         \switch_sel[4][1] , \switch_sel[4][0] , \switch_sel[3][4] ,
         \switch_sel[3][3] , \switch_sel[3][2] , \switch_sel[3][1] ,
         \switch_sel[3][0] , \switch_sel[2][4] , \switch_sel[2][3] ,
         \switch_sel[2][2] , \switch_sel[2][1] , \switch_sel[2][0] ,
         \switch_sel[1][4] , \switch_sel[1][3] , \switch_sel[1][2] ,
         \switch_sel[1][1] , \switch_sel[1][0] , \switch_sel[0][4] ,
         \switch_sel[0][3] , \switch_sel[0][2] , \switch_sel[0][1] ,
         \switch_sel[0][0] , \chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] ,
         \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] ,
         \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] ,
         \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] ,
         \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] ,
         \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] ,
         \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] ,
         \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] ,
         \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] ,
         \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] ,
         \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] ,
         \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] ,
         \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] ,
         \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] ,
         \chs_in_f[4][DATA][7] , \chs_in_f[4][DATA][6] ,
         \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] ,
         \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] ,
         \chs_in_f[4][DATA][1] , \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] ,
         \chs_in_f[3][DATA][34] , \chs_in_f[3][DATA][33] ,
         \chs_in_f[3][DATA][32] , \chs_in_f[3][DATA][31] ,
         \chs_in_f[3][DATA][30] , \chs_in_f[3][DATA][29] ,
         \chs_in_f[3][DATA][28] , \chs_in_f[3][DATA][27] ,
         \chs_in_f[3][DATA][26] , \chs_in_f[3][DATA][25] ,
         \chs_in_f[3][DATA][24] , \chs_in_f[3][DATA][23] ,
         \chs_in_f[3][DATA][22] , \chs_in_f[3][DATA][21] ,
         \chs_in_f[3][DATA][20] , \chs_in_f[3][DATA][19] ,
         \chs_in_f[3][DATA][18] , \chs_in_f[3][DATA][17] ,
         \chs_in_f[3][DATA][16] , \chs_in_f[3][DATA][15] ,
         \chs_in_f[3][DATA][14] , \chs_in_f[3][DATA][13] ,
         \chs_in_f[3][DATA][12] , \chs_in_f[3][DATA][11] ,
         \chs_in_f[3][DATA][10] , \chs_in_f[3][DATA][9] ,
         \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] ,
         \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] ,
         \chs_in_f[3][DATA][4] , \chs_in_f[3][DATA][3] ,
         \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] ,
         \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] ,
         \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] ,
         \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] ,
         \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] ,
         \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] ,
         \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] ,
         \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] ,
         \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] ,
         \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] ,
         \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] ,
         \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] ,
         \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] ,
         \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] ,
         \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] ,
         \chs_in_f[2][DATA][7] , \chs_in_f[2][DATA][6] ,
         \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] ,
         \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] ,
         \chs_in_f[2][DATA][1] , \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] ,
         \chs_in_f[1][DATA][34] , \chs_in_f[1][DATA][33] ,
         \chs_in_f[1][DATA][32] , \chs_in_f[1][DATA][31] ,
         \chs_in_f[1][DATA][30] , \chs_in_f[1][DATA][29] ,
         \chs_in_f[1][DATA][28] , \chs_in_f[1][DATA][27] ,
         \chs_in_f[1][DATA][26] , \chs_in_f[1][DATA][25] ,
         \chs_in_f[1][DATA][24] , \chs_in_f[1][DATA][23] ,
         \chs_in_f[1][DATA][22] , \chs_in_f[1][DATA][21] ,
         \chs_in_f[1][DATA][20] , \chs_in_f[1][DATA][19] ,
         \chs_in_f[1][DATA][18] , \chs_in_f[1][DATA][17] ,
         \chs_in_f[1][DATA][16] , \chs_in_f[1][DATA][15] ,
         \chs_in_f[1][DATA][14] , \chs_in_f[1][DATA][13] ,
         \chs_in_f[1][DATA][12] , \chs_in_f[1][DATA][11] ,
         \chs_in_f[1][DATA][10] , \chs_in_f[1][DATA][9] ,
         \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] ,
         \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] ,
         \chs_in_f[1][DATA][4] , \chs_in_f[1][DATA][3] ,
         \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] ,
         \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] ,
         \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] ,
         \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] ,
         \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] ,
         \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] ,
         \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] ,
         \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] ,
         \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] ,
         \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] ,
         \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] ,
         \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] ,
         \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] ,
         \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] ,
         \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] ,
         \chs_in_f[0][DATA][7] , \chs_in_f[0][DATA][6] ,
         \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] ,
         \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] ,
         \chs_in_f[0][DATA][1] , \chs_in_f[0][DATA][0] , \chs_out_b[4][ACK] ,
         \chs_out_b[3][ACK] , \chs_out_b[2][ACK] , \chs_out_b[1][ACK] ,
         \chs_out_b[0][ACK] ;
  output \chs_in_b[4][ACK] , \chs_in_b[3][ACK] , \chs_in_b[2][ACK] ,
         \chs_in_b[1][ACK] , \chs_in_b[0][ACK] , \chs_out_f[4][REQ] ,
         \chs_out_f[4][DATA][34] , \chs_out_f[4][DATA][33] ,
         \chs_out_f[4][DATA][32] , \chs_out_f[4][DATA][31] ,
         \chs_out_f[4][DATA][30] , \chs_out_f[4][DATA][29] ,
         \chs_out_f[4][DATA][28] , \chs_out_f[4][DATA][27] ,
         \chs_out_f[4][DATA][26] , \chs_out_f[4][DATA][25] ,
         \chs_out_f[4][DATA][24] , \chs_out_f[4][DATA][23] ,
         \chs_out_f[4][DATA][22] , \chs_out_f[4][DATA][21] ,
         \chs_out_f[4][DATA][20] , \chs_out_f[4][DATA][19] ,
         \chs_out_f[4][DATA][18] , \chs_out_f[4][DATA][17] ,
         \chs_out_f[4][DATA][16] , \chs_out_f[4][DATA][15] ,
         \chs_out_f[4][DATA][14] , \chs_out_f[4][DATA][13] ,
         \chs_out_f[4][DATA][12] , \chs_out_f[4][DATA][11] ,
         \chs_out_f[4][DATA][10] , \chs_out_f[4][DATA][9] ,
         \chs_out_f[4][DATA][8] , \chs_out_f[4][DATA][7] ,
         \chs_out_f[4][DATA][6] , \chs_out_f[4][DATA][5] ,
         \chs_out_f[4][DATA][4] , \chs_out_f[4][DATA][3] ,
         \chs_out_f[4][DATA][2] , \chs_out_f[4][DATA][1] ,
         \chs_out_f[4][DATA][0] , \chs_out_f[3][REQ] ,
         \chs_out_f[3][DATA][34] , \chs_out_f[3][DATA][33] ,
         \chs_out_f[3][DATA][32] , \chs_out_f[3][DATA][31] ,
         \chs_out_f[3][DATA][30] , \chs_out_f[3][DATA][29] ,
         \chs_out_f[3][DATA][28] , \chs_out_f[3][DATA][27] ,
         \chs_out_f[3][DATA][26] , \chs_out_f[3][DATA][25] ,
         \chs_out_f[3][DATA][24] , \chs_out_f[3][DATA][23] ,
         \chs_out_f[3][DATA][22] , \chs_out_f[3][DATA][21] ,
         \chs_out_f[3][DATA][20] , \chs_out_f[3][DATA][19] ,
         \chs_out_f[3][DATA][18] , \chs_out_f[3][DATA][17] ,
         \chs_out_f[3][DATA][16] , \chs_out_f[3][DATA][15] ,
         \chs_out_f[3][DATA][14] , \chs_out_f[3][DATA][13] ,
         \chs_out_f[3][DATA][12] , \chs_out_f[3][DATA][11] ,
         \chs_out_f[3][DATA][10] , \chs_out_f[3][DATA][9] ,
         \chs_out_f[3][DATA][8] , \chs_out_f[3][DATA][7] ,
         \chs_out_f[3][DATA][6] , \chs_out_f[3][DATA][5] ,
         \chs_out_f[3][DATA][4] , \chs_out_f[3][DATA][3] ,
         \chs_out_f[3][DATA][2] , \chs_out_f[3][DATA][1] ,
         \chs_out_f[3][DATA][0] , \chs_out_f[2][REQ] ,
         \chs_out_f[2][DATA][34] , \chs_out_f[2][DATA][33] ,
         \chs_out_f[2][DATA][32] , \chs_out_f[2][DATA][31] ,
         \chs_out_f[2][DATA][30] , \chs_out_f[2][DATA][29] ,
         \chs_out_f[2][DATA][28] , \chs_out_f[2][DATA][27] ,
         \chs_out_f[2][DATA][26] , \chs_out_f[2][DATA][25] ,
         \chs_out_f[2][DATA][24] , \chs_out_f[2][DATA][23] ,
         \chs_out_f[2][DATA][22] , \chs_out_f[2][DATA][21] ,
         \chs_out_f[2][DATA][20] , \chs_out_f[2][DATA][19] ,
         \chs_out_f[2][DATA][18] , \chs_out_f[2][DATA][17] ,
         \chs_out_f[2][DATA][16] , \chs_out_f[2][DATA][15] ,
         \chs_out_f[2][DATA][14] , \chs_out_f[2][DATA][13] ,
         \chs_out_f[2][DATA][12] , \chs_out_f[2][DATA][11] ,
         \chs_out_f[2][DATA][10] , \chs_out_f[2][DATA][9] ,
         \chs_out_f[2][DATA][8] , \chs_out_f[2][DATA][7] ,
         \chs_out_f[2][DATA][6] , \chs_out_f[2][DATA][5] ,
         \chs_out_f[2][DATA][4] , \chs_out_f[2][DATA][3] ,
         \chs_out_f[2][DATA][2] , \chs_out_f[2][DATA][1] ,
         \chs_out_f[2][DATA][0] , \chs_out_f[1][REQ] ,
         \chs_out_f[1][DATA][34] , \chs_out_f[1][DATA][33] ,
         \chs_out_f[1][DATA][32] , \chs_out_f[1][DATA][31] ,
         \chs_out_f[1][DATA][30] , \chs_out_f[1][DATA][29] ,
         \chs_out_f[1][DATA][28] , \chs_out_f[1][DATA][27] ,
         \chs_out_f[1][DATA][26] , \chs_out_f[1][DATA][25] ,
         \chs_out_f[1][DATA][24] , \chs_out_f[1][DATA][23] ,
         \chs_out_f[1][DATA][22] , \chs_out_f[1][DATA][21] ,
         \chs_out_f[1][DATA][20] , \chs_out_f[1][DATA][19] ,
         \chs_out_f[1][DATA][18] , \chs_out_f[1][DATA][17] ,
         \chs_out_f[1][DATA][16] , \chs_out_f[1][DATA][15] ,
         \chs_out_f[1][DATA][14] , \chs_out_f[1][DATA][13] ,
         \chs_out_f[1][DATA][12] , \chs_out_f[1][DATA][11] ,
         \chs_out_f[1][DATA][10] , \chs_out_f[1][DATA][9] ,
         \chs_out_f[1][DATA][8] , \chs_out_f[1][DATA][7] ,
         \chs_out_f[1][DATA][6] , \chs_out_f[1][DATA][5] ,
         \chs_out_f[1][DATA][4] , \chs_out_f[1][DATA][3] ,
         \chs_out_f[1][DATA][2] , \chs_out_f[1][DATA][1] ,
         \chs_out_f[1][DATA][0] , \chs_out_f[0][REQ] ,
         \chs_out_f[0][DATA][34] , \chs_out_f[0][DATA][33] ,
         \chs_out_f[0][DATA][32] , \chs_out_f[0][DATA][31] ,
         \chs_out_f[0][DATA][30] , \chs_out_f[0][DATA][29] ,
         \chs_out_f[0][DATA][28] , \chs_out_f[0][DATA][27] ,
         \chs_out_f[0][DATA][26] , \chs_out_f[0][DATA][25] ,
         \chs_out_f[0][DATA][24] , \chs_out_f[0][DATA][23] ,
         \chs_out_f[0][DATA][22] , \chs_out_f[0][DATA][21] ,
         \chs_out_f[0][DATA][20] , \chs_out_f[0][DATA][19] ,
         \chs_out_f[0][DATA][18] , \chs_out_f[0][DATA][17] ,
         \chs_out_f[0][DATA][16] , \chs_out_f[0][DATA][15] ,
         \chs_out_f[0][DATA][14] , \chs_out_f[0][DATA][13] ,
         \chs_out_f[0][DATA][12] , \chs_out_f[0][DATA][11] ,
         \chs_out_f[0][DATA][10] , \chs_out_f[0][DATA][9] ,
         \chs_out_f[0][DATA][8] , \chs_out_f[0][DATA][7] ,
         \chs_out_f[0][DATA][6] , \chs_out_f[0][DATA][5] ,
         \chs_out_f[0][DATA][4] , \chs_out_f[0][DATA][3] ,
         \chs_out_f[0][DATA][2] , \chs_out_f[0][DATA][1] ,
         \chs_out_f[0][DATA][0] ;
  wire   \chs_in_b[4][ACK] , \chs_out_f[4][REQ] , synced_req, del, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335;
  assign \chs_in_b[0][ACK]  = \chs_in_b[4][ACK] ;
  assign \chs_in_b[1][ACK]  = \chs_in_b[4][ACK] ;
  assign \chs_in_b[2][ACK]  = \chs_in_b[4][ACK] ;
  assign \chs_in_b[3][ACK]  = \chs_in_b[4][ACK] ;
  assign \chs_out_f[0][REQ]  = \chs_out_f[4][REQ] ;
  assign \chs_out_f[1][REQ]  = \chs_out_f[4][REQ] ;
  assign \chs_out_f[2][REQ]  = \chs_out_f[4][REQ] ;
  assign \chs_out_f[3][REQ]  = \chs_out_f[4][REQ] ;

  c_gate_generic_1_5_0 c_sync_req ( .preset(preset), .\input ({
        \chs_in_f[4][REQ] , \chs_in_f[3][REQ] , \chs_in_f[2][REQ] , 
        \chs_in_f[1][REQ] , \chs_in_f[0][REQ] }), .\output (synced_req) );
  c_gate_generic_1_5_7 c_sync_ack ( .preset(preset), .\input ({
        \chs_out_b[4][ACK] , \chs_out_b[3][ACK] , \chs_out_b[2][ACK] , 
        \chs_out_b[1][ACK] , \chs_out_b[0][ACK] }), .\output (
        \chs_in_b[4][ACK] ) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chs_out_f[4][REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(synced_req), .Z(del) );
  HS65_LS_IVX9 U2 ( .A(\switch_sel[3][2] ), .Z(n332) );
  HS65_LS_IVX9 U3 ( .A(\switch_sel[3][1] ), .Z(n333) );
  HS65_LS_IVX9 U4 ( .A(\switch_sel[3][0] ), .Z(n334) );
  HS65_LS_IVX9 U5 ( .A(\switch_sel[3][4] ), .Z(n331) );
  HS65_LS_BFX9 U6 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U7 ( .A(del), .Z(n2) );
  HS65_LS_BFX7 U8 ( .A(n329), .Z(n12) );
  HS65_LS_BFX7 U9 ( .A(n329), .Z(n13) );
  HS65_LS_BFX9 U10 ( .A(\switch_sel[0][3] ), .Z(n41) );
  HS65_LS_BFX9 U11 ( .A(\switch_sel[1][3] ), .Z(n57) );
  HS65_LS_BFX9 U12 ( .A(\switch_sel[1][2] ), .Z(n53) );
  HS65_LS_BFX9 U13 ( .A(\switch_sel[0][1] ), .Z(n33) );
  HS65_LS_BFX9 U14 ( .A(\switch_sel[1][0] ), .Z(n49) );
  HS65_LS_BFX9 U15 ( .A(\switch_sel[0][4] ), .Z(n45) );
  HS65_LS_BFX9 U16 ( .A(\switch_sel[1][4] ), .Z(n61) );
  HS65_LS_BFX9 U17 ( .A(n331), .Z(n18) );
  HS65_LS_BFX9 U18 ( .A(n331), .Z(n19) );
  HS65_LS_BFX9 U19 ( .A(n61), .Z(n62) );
  HS65_LS_BFX9 U20 ( .A(n61), .Z(n63) );
  HS65_LS_BFX9 U21 ( .A(n77), .Z(n78) );
  HS65_LS_BFX9 U22 ( .A(n77), .Z(n79) );
  HS65_LS_BFX9 U23 ( .A(n45), .Z(n46) );
  HS65_LS_BFX9 U24 ( .A(n45), .Z(n47) );
  HS65_LS_BFX9 U25 ( .A(n332), .Z(n21) );
  HS65_LS_BFX9 U26 ( .A(n332), .Z(n22) );
  HS65_LS_BFX9 U27 ( .A(n333), .Z(n24) );
  HS65_LS_BFX9 U28 ( .A(n333), .Z(n25) );
  HS65_LS_BFX9 U29 ( .A(n334), .Z(n27) );
  HS65_LS_BFX9 U30 ( .A(n334), .Z(n28) );
  HS65_LS_BFX9 U31 ( .A(n57), .Z(n58) );
  HS65_LS_BFX9 U32 ( .A(n57), .Z(n59) );
  HS65_LS_BFX9 U33 ( .A(n53), .Z(n54) );
  HS65_LS_BFX9 U34 ( .A(n53), .Z(n55) );
  HS65_LS_BFX9 U35 ( .A(n49), .Z(n50) );
  HS65_LS_BFX9 U36 ( .A(n49), .Z(n51) );
  HS65_LS_BFX9 U37 ( .A(n73), .Z(n74) );
  HS65_LS_BFX9 U38 ( .A(n73), .Z(n75) );
  HS65_LS_BFX9 U39 ( .A(n69), .Z(n70) );
  HS65_LS_BFX9 U40 ( .A(n69), .Z(n71) );
  HS65_LS_BFX9 U41 ( .A(n65), .Z(n66) );
  HS65_LS_BFX9 U42 ( .A(n65), .Z(n67) );
  HS65_LS_BFX9 U43 ( .A(n331), .Z(n20) );
  HS65_LS_BFX9 U44 ( .A(n41), .Z(n42) );
  HS65_LS_BFX9 U45 ( .A(n41), .Z(n43) );
  HS65_LS_BFX9 U46 ( .A(n37), .Z(n38) );
  HS65_LS_BFX9 U47 ( .A(n37), .Z(n39) );
  HS65_LS_BFX9 U48 ( .A(n33), .Z(n34) );
  HS65_LS_BFX9 U49 ( .A(n33), .Z(n35) );
  HS65_LS_BFX9 U50 ( .A(n45), .Z(n48) );
  HS65_LS_BFX9 U51 ( .A(n326), .Z(n3) );
  HS65_LS_BFX9 U52 ( .A(n326), .Z(n4) );
  HS65_LS_BFX9 U53 ( .A(n327), .Z(n6) );
  HS65_LS_BFX9 U54 ( .A(n327), .Z(n7) );
  HS65_LS_BFX9 U55 ( .A(n328), .Z(n9) );
  HS65_LS_BFX9 U56 ( .A(n328), .Z(n10) );
  HS65_LS_BFX9 U57 ( .A(n57), .Z(n60) );
  HS65_LS_BFX9 U58 ( .A(n53), .Z(n56) );
  HS65_LS_BFX9 U59 ( .A(n49), .Z(n52) );
  HS65_LS_BFX9 U60 ( .A(n73), .Z(n76) );
  HS65_LS_BFX9 U61 ( .A(n69), .Z(n72) );
  HS65_LS_BFX9 U62 ( .A(n65), .Z(n68) );
  HS65_LS_BFX9 U63 ( .A(n41), .Z(n44) );
  HS65_LS_BFX9 U64 ( .A(n37), .Z(n40) );
  HS65_LS_BFX9 U65 ( .A(n33), .Z(n36) );
  HS65_LS_BFX9 U66 ( .A(n326), .Z(n5) );
  HS65_LS_BFX9 U67 ( .A(n327), .Z(n8) );
  HS65_LS_BFX9 U68 ( .A(n328), .Z(n11) );
  HS65_LS_BFX9 U69 ( .A(n329), .Z(n14) );
  HS65_LS_BFX9 U70 ( .A(n332), .Z(n23) );
  HS65_LS_BFX9 U71 ( .A(n333), .Z(n26) );
  HS65_LS_BFX9 U72 ( .A(n334), .Z(n29) );
  HS65_LS_BFX9 U73 ( .A(n61), .Z(n64) );
  HS65_LS_BFX9 U74 ( .A(n77), .Z(n80) );
  HS65_LS_BFX9 U75 ( .A(n330), .Z(n15) );
  HS65_LS_BFX9 U76 ( .A(n330), .Z(n16) );
  HS65_LS_BFX9 U77 ( .A(n335), .Z(n30) );
  HS65_LS_BFX9 U78 ( .A(n335), .Z(n31) );
  HS65_LS_BFX9 U79 ( .A(n330), .Z(n17) );
  HS65_LS_BFX9 U80 ( .A(n335), .Z(n32) );
  HS65_LS_IVX9 U81 ( .A(\switch_sel[4][3] ), .Z(n326) );
  HS65_LS_IVX9 U82 ( .A(\switch_sel[4][2] ), .Z(n327) );
  HS65_LS_IVX9 U83 ( .A(\switch_sel[4][1] ), .Z(n328) );
  HS65_LS_IVX9 U84 ( .A(\switch_sel[4][0] ), .Z(n329) );
  HS65_LS_AOI222X2 U85 ( .A(\chs_in_f[2][DATA][34] ), .B(n78), .C(
        \chs_in_f[0][DATA][34] ), .D(n48), .E(\chs_in_f[1][DATA][34] ), .F(n62), .Z(n88) );
  HS65_LS_OAI212X5 U86 ( .A(n281), .B(n20), .C(n316), .D(n17), .E(n81), .Z(
        \chs_out_f[4][DATA][9] ) );
  HS65_LS_AOI222X2 U87 ( .A(n78), .B(\chs_in_f[2][DATA][9] ), .C(n48), .D(
        \chs_in_f[0][DATA][9] ), .E(n62), .F(\chs_in_f[1][DATA][9] ), .Z(n81)
         );
  HS65_LS_AOI222X2 U88 ( .A(n76), .B(\chs_in_f[2][DATA][34] ), .C(n44), .D(
        \chs_in_f[0][DATA][34] ), .E(n60), .F(\chs_in_f[1][DATA][34] ), .Z(
        n123) );
  HS65_LS_AOI222X2 U89 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][34] ), 
        .C(n40), .D(\chs_in_f[0][DATA][34] ), .E(n56), .F(
        \chs_in_f[1][DATA][34] ), .Z(n158) );
  HS65_LS_AOI222X2 U90 ( .A(n72), .B(\chs_in_f[2][DATA][34] ), .C(n36), .D(
        \chs_in_f[0][DATA][34] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][34] ), .Z(n193) );
  HS65_LS_AOI222X2 U91 ( .A(n68), .B(\chs_in_f[2][DATA][34] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][34] ), .E(n52), .F(
        \chs_in_f[1][DATA][34] ), .Z(n228) );
  HS65_LS_IVX9 U92 ( .A(\chs_in_f[3][DATA][9] ), .Z(n281) );
  HS65_LS_IVX9 U93 ( .A(\chs_in_f[3][DATA][34] ), .Z(n256) );
  HS65_LS_IVX9 U94 ( .A(\chs_in_f[3][DATA][0] ), .Z(n290) );
  HS65_LS_IVX9 U95 ( .A(\chs_in_f[3][DATA][1] ), .Z(n289) );
  HS65_LS_IVX9 U96 ( .A(\chs_in_f[3][DATA][2] ), .Z(n288) );
  HS65_LS_IVX9 U97 ( .A(\chs_in_f[3][DATA][3] ), .Z(n287) );
  HS65_LS_IVX9 U98 ( .A(\chs_in_f[3][DATA][4] ), .Z(n286) );
  HS65_LS_IVX9 U99 ( .A(\chs_in_f[3][DATA][5] ), .Z(n285) );
  HS65_LS_IVX9 U100 ( .A(\chs_in_f[3][DATA][6] ), .Z(n284) );
  HS65_LS_IVX9 U101 ( .A(\chs_in_f[3][DATA][7] ), .Z(n283) );
  HS65_LS_IVX9 U102 ( .A(\chs_in_f[3][DATA][8] ), .Z(n282) );
  HS65_LS_IVX9 U103 ( .A(\chs_in_f[3][DATA][10] ), .Z(n280) );
  HS65_LS_IVX9 U104 ( .A(\chs_in_f[3][DATA][11] ), .Z(n279) );
  HS65_LS_IVX9 U105 ( .A(\chs_in_f[3][DATA][12] ), .Z(n278) );
  HS65_LS_IVX9 U106 ( .A(\chs_in_f[3][DATA][13] ), .Z(n277) );
  HS65_LS_IVX9 U107 ( .A(\chs_in_f[3][DATA][14] ), .Z(n276) );
  HS65_LS_IVX9 U108 ( .A(\chs_in_f[3][DATA][15] ), .Z(n275) );
  HS65_LS_IVX9 U109 ( .A(\chs_in_f[3][DATA][16] ), .Z(n274) );
  HS65_LS_IVX9 U110 ( .A(\chs_in_f[3][DATA][17] ), .Z(n273) );
  HS65_LS_IVX9 U111 ( .A(\chs_in_f[3][DATA][18] ), .Z(n272) );
  HS65_LS_IVX9 U112 ( .A(\chs_in_f[3][DATA][19] ), .Z(n271) );
  HS65_LS_IVX9 U113 ( .A(\chs_in_f[3][DATA][20] ), .Z(n270) );
  HS65_LS_IVX9 U114 ( .A(\chs_in_f[3][DATA][21] ), .Z(n269) );
  HS65_LS_IVX9 U115 ( .A(\chs_in_f[3][DATA][22] ), .Z(n268) );
  HS65_LS_IVX9 U116 ( .A(\chs_in_f[3][DATA][23] ), .Z(n267) );
  HS65_LS_IVX9 U117 ( .A(\chs_in_f[3][DATA][24] ), .Z(n266) );
  HS65_LS_IVX9 U118 ( .A(\chs_in_f[3][DATA][25] ), .Z(n265) );
  HS65_LS_IVX9 U119 ( .A(\chs_in_f[3][DATA][26] ), .Z(n264) );
  HS65_LS_IVX9 U120 ( .A(\chs_in_f[3][DATA][27] ), .Z(n263) );
  HS65_LS_IVX9 U121 ( .A(\chs_in_f[3][DATA][28] ), .Z(n262) );
  HS65_LS_IVX9 U122 ( .A(\chs_in_f[3][DATA][29] ), .Z(n261) );
  HS65_LS_IVX9 U123 ( .A(\chs_in_f[3][DATA][30] ), .Z(n260) );
  HS65_LS_IVX9 U124 ( .A(\chs_in_f[3][DATA][31] ), .Z(n259) );
  HS65_LS_IVX9 U125 ( .A(\chs_in_f[3][DATA][32] ), .Z(n258) );
  HS65_LS_IVX9 U126 ( .A(\chs_in_f[3][DATA][33] ), .Z(n257) );
  HS65_LS_IVX9 U127 ( .A(\chs_in_f[4][DATA][9] ), .Z(n316) );
  HS65_LS_IVX9 U128 ( .A(\chs_in_f[4][DATA][34] ), .Z(n291) );
  HS65_LS_IVX9 U129 ( .A(\chs_in_f[4][DATA][0] ), .Z(n325) );
  HS65_LS_IVX9 U130 ( .A(\chs_in_f[4][DATA][1] ), .Z(n324) );
  HS65_LS_IVX9 U131 ( .A(\chs_in_f[4][DATA][2] ), .Z(n323) );
  HS65_LS_IVX9 U132 ( .A(\chs_in_f[4][DATA][3] ), .Z(n322) );
  HS65_LS_IVX9 U133 ( .A(\chs_in_f[4][DATA][4] ), .Z(n321) );
  HS65_LS_IVX9 U134 ( .A(\chs_in_f[4][DATA][5] ), .Z(n320) );
  HS65_LS_IVX9 U135 ( .A(\chs_in_f[4][DATA][6] ), .Z(n319) );
  HS65_LS_IVX9 U136 ( .A(\chs_in_f[4][DATA][7] ), .Z(n318) );
  HS65_LS_IVX9 U137 ( .A(\chs_in_f[4][DATA][8] ), .Z(n317) );
  HS65_LS_IVX9 U138 ( .A(\chs_in_f[4][DATA][10] ), .Z(n315) );
  HS65_LS_IVX9 U139 ( .A(\chs_in_f[4][DATA][11] ), .Z(n314) );
  HS65_LS_IVX9 U140 ( .A(\chs_in_f[4][DATA][12] ), .Z(n313) );
  HS65_LS_IVX9 U141 ( .A(\chs_in_f[4][DATA][13] ), .Z(n312) );
  HS65_LS_IVX9 U142 ( .A(\chs_in_f[4][DATA][14] ), .Z(n311) );
  HS65_LS_IVX9 U143 ( .A(\chs_in_f[4][DATA][15] ), .Z(n310) );
  HS65_LS_IVX9 U144 ( .A(\chs_in_f[4][DATA][33] ), .Z(n292) );
  HS65_LS_IVX9 U145 ( .A(\chs_in_f[4][DATA][16] ), .Z(n309) );
  HS65_LS_IVX9 U146 ( .A(\chs_in_f[4][DATA][17] ), .Z(n308) );
  HS65_LS_IVX9 U147 ( .A(\chs_in_f[4][DATA][18] ), .Z(n307) );
  HS65_LS_IVX9 U148 ( .A(\chs_in_f[4][DATA][19] ), .Z(n306) );
  HS65_LS_IVX9 U149 ( .A(\chs_in_f[4][DATA][20] ), .Z(n305) );
  HS65_LS_IVX9 U150 ( .A(\chs_in_f[4][DATA][21] ), .Z(n304) );
  HS65_LS_IVX9 U151 ( .A(\chs_in_f[4][DATA][22] ), .Z(n303) );
  HS65_LS_IVX9 U152 ( .A(\chs_in_f[4][DATA][23] ), .Z(n302) );
  HS65_LS_IVX9 U153 ( .A(\chs_in_f[4][DATA][24] ), .Z(n301) );
  HS65_LS_IVX9 U154 ( .A(\chs_in_f[4][DATA][25] ), .Z(n300) );
  HS65_LS_IVX9 U155 ( .A(\chs_in_f[4][DATA][26] ), .Z(n299) );
  HS65_LS_IVX9 U156 ( .A(\chs_in_f[4][DATA][27] ), .Z(n298) );
  HS65_LS_IVX9 U157 ( .A(\chs_in_f[4][DATA][28] ), .Z(n297) );
  HS65_LS_IVX9 U158 ( .A(\chs_in_f[4][DATA][29] ), .Z(n296) );
  HS65_LS_IVX9 U159 ( .A(\chs_in_f[4][DATA][30] ), .Z(n295) );
  HS65_LS_IVX9 U160 ( .A(\chs_in_f[4][DATA][31] ), .Z(n294) );
  HS65_LS_IVX9 U161 ( .A(\chs_in_f[4][DATA][32] ), .Z(n293) );
  HS65_LS_BFX18 U162 ( .A(\switch_sel[2][3] ), .Z(n73) );
  HS65_LS_BFX18 U163 ( .A(\switch_sel[0][2] ), .Z(n37) );
  HS65_LS_BFX18 U164 ( .A(\switch_sel[2][1] ), .Z(n69) );
  HS65_LS_BFX18 U165 ( .A(\switch_sel[2][0] ), .Z(n65) );
  HS65_LS_BFX18 U166 ( .A(\switch_sel[2][4] ), .Z(n77) );
  HS65_LS_OAI212X5 U167 ( .A(n18), .B(n290), .C(n15), .D(n325), .E(n115), .Z(
        \chs_out_f[4][DATA][0] ) );
  HS65_LS_AOI222X2 U168 ( .A(\chs_in_f[2][DATA][0] ), .B(n80), .C(
        \chs_in_f[0][DATA][0] ), .D(n46), .E(\chs_in_f[1][DATA][0] ), .F(n64), 
        .Z(n115) );
  HS65_LS_OAI212X5 U169 ( .A(n18), .B(n289), .C(n15), .D(n324), .E(n104), .Z(
        \chs_out_f[4][DATA][1] ) );
  HS65_LS_AOI222X2 U170 ( .A(\chs_in_f[2][DATA][1] ), .B(n79), .C(
        \chs_in_f[0][DATA][1] ), .D(n46), .E(\chs_in_f[1][DATA][1] ), .F(n63), 
        .Z(n104) );
  HS65_LS_OAI212X5 U171 ( .A(n19), .B(n288), .C(n16), .D(n323), .E(n93), .Z(
        \chs_out_f[4][DATA][2] ) );
  HS65_LS_AOI222X2 U172 ( .A(\chs_in_f[2][DATA][2] ), .B(n78), .C(
        \chs_in_f[0][DATA][2] ), .D(n47), .E(\chs_in_f[1][DATA][2] ), .F(n62), 
        .Z(n93) );
  HS65_LS_OAI212X5 U173 ( .A(n20), .B(n287), .C(n17), .D(n322), .E(n87), .Z(
        \chs_out_f[4][DATA][3] ) );
  HS65_LS_AOI222X2 U174 ( .A(\chs_in_f[2][DATA][3] ), .B(n78), .C(
        \chs_in_f[0][DATA][3] ), .D(n48), .E(\chs_in_f[1][DATA][3] ), .F(n62), 
        .Z(n87) );
  HS65_LS_OAI212X5 U175 ( .A(n20), .B(n286), .C(n17), .D(n321), .E(n86), .Z(
        \chs_out_f[4][DATA][4] ) );
  HS65_LS_AOI222X2 U176 ( .A(\chs_in_f[2][DATA][4] ), .B(n78), .C(
        \chs_in_f[0][DATA][4] ), .D(n48), .E(\chs_in_f[1][DATA][4] ), .F(n62), 
        .Z(n86) );
  HS65_LS_OAI212X5 U177 ( .A(n20), .B(n285), .C(n17), .D(n320), .E(n85), .Z(
        \chs_out_f[4][DATA][5] ) );
  HS65_LS_AOI222X2 U178 ( .A(\chs_in_f[2][DATA][5] ), .B(n78), .C(
        \chs_in_f[0][DATA][5] ), .D(n48), .E(\chs_in_f[1][DATA][5] ), .F(n62), 
        .Z(n85) );
  HS65_LS_OAI212X5 U179 ( .A(n20), .B(n284), .C(n17), .D(n319), .E(n84), .Z(
        \chs_out_f[4][DATA][6] ) );
  HS65_LS_AOI222X2 U180 ( .A(\chs_in_f[2][DATA][6] ), .B(n78), .C(
        \chs_in_f[0][DATA][6] ), .D(n48), .E(\chs_in_f[1][DATA][6] ), .F(n62), 
        .Z(n84) );
  HS65_LS_OAI212X5 U181 ( .A(n20), .B(n283), .C(n17), .D(n318), .E(n83), .Z(
        \chs_out_f[4][DATA][7] ) );
  HS65_LS_AOI222X2 U182 ( .A(\chs_in_f[2][DATA][7] ), .B(n78), .C(
        \chs_in_f[0][DATA][7] ), .D(n48), .E(\chs_in_f[1][DATA][7] ), .F(n62), 
        .Z(n83) );
  HS65_LS_OAI212X5 U183 ( .A(n20), .B(n282), .C(n17), .D(n317), .E(n82), .Z(
        \chs_out_f[4][DATA][8] ) );
  HS65_LS_AOI222X2 U184 ( .A(\chs_in_f[2][DATA][8] ), .B(n78), .C(
        \chs_in_f[0][DATA][8] ), .D(n48), .E(\chs_in_f[1][DATA][8] ), .F(n62), 
        .Z(n82) );
  HS65_LS_OAI212X5 U185 ( .A(n18), .B(n280), .C(n15), .D(n315), .E(n114), .Z(
        \chs_out_f[4][DATA][10] ) );
  HS65_LS_AOI222X2 U186 ( .A(\chs_in_f[2][DATA][10] ), .B(n80), .C(
        \chs_in_f[0][DATA][10] ), .D(n46), .E(\chs_in_f[1][DATA][10] ), .F(n64), .Z(n114) );
  HS65_LS_OAI212X5 U187 ( .A(n18), .B(n279), .C(n15), .D(n314), .E(n113), .Z(
        \chs_out_f[4][DATA][11] ) );
  HS65_LS_AOI222X2 U188 ( .A(\chs_in_f[2][DATA][11] ), .B(n80), .C(
        \chs_in_f[0][DATA][11] ), .D(n46), .E(\chs_in_f[1][DATA][11] ), .F(n64), .Z(n113) );
  HS65_LS_OAI212X5 U189 ( .A(n18), .B(n278), .C(n15), .D(n313), .E(n112), .Z(
        \chs_out_f[4][DATA][12] ) );
  HS65_LS_AOI222X2 U190 ( .A(\chs_in_f[2][DATA][12] ), .B(n80), .C(
        \chs_in_f[0][DATA][12] ), .D(n46), .E(\chs_in_f[1][DATA][12] ), .F(n64), .Z(n112) );
  HS65_LS_OAI212X5 U191 ( .A(n18), .B(n277), .C(n15), .D(n312), .E(n111), .Z(
        \chs_out_f[4][DATA][13] ) );
  HS65_LS_AOI222X2 U192 ( .A(\chs_in_f[2][DATA][13] ), .B(n80), .C(
        \chs_in_f[0][DATA][13] ), .D(n46), .E(\chs_in_f[1][DATA][13] ), .F(n64), .Z(n111) );
  HS65_LS_OAI212X5 U193 ( .A(n18), .B(n276), .C(n15), .D(n311), .E(n110), .Z(
        \chs_out_f[4][DATA][14] ) );
  HS65_LS_AOI222X2 U194 ( .A(\chs_in_f[2][DATA][14] ), .B(n80), .C(
        \chs_in_f[0][DATA][14] ), .D(n46), .E(\chs_in_f[1][DATA][14] ), .F(n64), .Z(n110) );
  HS65_LS_OAI212X5 U195 ( .A(n18), .B(n275), .C(n15), .D(n310), .E(n109), .Z(
        \chs_out_f[4][DATA][15] ) );
  HS65_LS_AOI222X2 U196 ( .A(\chs_in_f[2][DATA][15] ), .B(n80), .C(
        \chs_in_f[0][DATA][15] ), .D(n46), .E(\chs_in_f[1][DATA][15] ), .F(n64), .Z(n109) );
  HS65_LS_OAI212X5 U197 ( .A(n18), .B(n274), .C(n15), .D(n309), .E(n108), .Z(
        \chs_out_f[4][DATA][16] ) );
  HS65_LS_AOI222X2 U198 ( .A(\chs_in_f[2][DATA][16] ), .B(n80), .C(
        \chs_in_f[0][DATA][16] ), .D(n46), .E(\chs_in_f[1][DATA][16] ), .F(n64), .Z(n108) );
  HS65_LS_OAI212X5 U199 ( .A(n18), .B(n273), .C(n15), .D(n308), .E(n107), .Z(
        \chs_out_f[4][DATA][17] ) );
  HS65_LS_AOI222X2 U200 ( .A(\chs_in_f[2][DATA][17] ), .B(n80), .C(
        \chs_in_f[0][DATA][17] ), .D(n46), .E(\chs_in_f[1][DATA][17] ), .F(n64), .Z(n107) );
  HS65_LS_OAI212X5 U201 ( .A(n18), .B(n272), .C(n15), .D(n307), .E(n106), .Z(
        \chs_out_f[4][DATA][18] ) );
  HS65_LS_AOI222X2 U202 ( .A(\chs_in_f[2][DATA][18] ), .B(n79), .C(
        \chs_in_f[0][DATA][18] ), .D(n46), .E(\chs_in_f[1][DATA][18] ), .F(n63), .Z(n106) );
  HS65_LS_OAI212X5 U203 ( .A(n18), .B(n271), .C(n15), .D(n306), .E(n105), .Z(
        \chs_out_f[4][DATA][19] ) );
  HS65_LS_AOI222X2 U204 ( .A(\chs_in_f[2][DATA][19] ), .B(n79), .C(
        \chs_in_f[0][DATA][19] ), .D(n46), .E(\chs_in_f[1][DATA][19] ), .F(n63), .Z(n105) );
  HS65_LS_OAI212X5 U205 ( .A(n19), .B(n270), .C(n15), .D(n305), .E(n103), .Z(
        \chs_out_f[4][DATA][20] ) );
  HS65_LS_AOI222X2 U206 ( .A(\chs_in_f[2][DATA][20] ), .B(n79), .C(
        \chs_in_f[0][DATA][20] ), .D(n47), .E(\chs_in_f[1][DATA][20] ), .F(n63), .Z(n103) );
  HS65_LS_OAI212X5 U207 ( .A(n19), .B(n269), .C(n16), .D(n304), .E(n102), .Z(
        \chs_out_f[4][DATA][21] ) );
  HS65_LS_AOI222X2 U208 ( .A(\chs_in_f[2][DATA][21] ), .B(n79), .C(
        \chs_in_f[0][DATA][21] ), .D(n47), .E(\chs_in_f[1][DATA][21] ), .F(n63), .Z(n102) );
  HS65_LS_OAI212X5 U209 ( .A(n19), .B(n268), .C(n16), .D(n303), .E(n101), .Z(
        \chs_out_f[4][DATA][22] ) );
  HS65_LS_AOI222X2 U210 ( .A(\chs_in_f[2][DATA][22] ), .B(n79), .C(
        \chs_in_f[0][DATA][22] ), .D(n47), .E(\chs_in_f[1][DATA][22] ), .F(n63), .Z(n101) );
  HS65_LS_OAI212X5 U211 ( .A(n19), .B(n267), .C(n16), .D(n302), .E(n100), .Z(
        \chs_out_f[4][DATA][23] ) );
  HS65_LS_AOI222X2 U212 ( .A(\chs_in_f[2][DATA][23] ), .B(n79), .C(
        \chs_in_f[0][DATA][23] ), .D(n47), .E(\chs_in_f[1][DATA][23] ), .F(n63), .Z(n100) );
  HS65_LS_OAI212X5 U213 ( .A(n19), .B(n266), .C(n16), .D(n301), .E(n99), .Z(
        \chs_out_f[4][DATA][24] ) );
  HS65_LS_AOI222X2 U214 ( .A(\chs_in_f[2][DATA][24] ), .B(n79), .C(
        \chs_in_f[0][DATA][24] ), .D(n47), .E(\chs_in_f[1][DATA][24] ), .F(n63), .Z(n99) );
  HS65_LS_OAI212X5 U215 ( .A(n19), .B(n265), .C(n16), .D(n300), .E(n98), .Z(
        \chs_out_f[4][DATA][25] ) );
  HS65_LS_AOI222X2 U216 ( .A(\chs_in_f[2][DATA][25] ), .B(n79), .C(
        \chs_in_f[0][DATA][25] ), .D(n47), .E(\chs_in_f[1][DATA][25] ), .F(n63), .Z(n98) );
  HS65_LS_OAI212X5 U217 ( .A(n19), .B(n264), .C(n16), .D(n299), .E(n97), .Z(
        \chs_out_f[4][DATA][26] ) );
  HS65_LS_AOI222X2 U218 ( .A(\chs_in_f[2][DATA][26] ), .B(n79), .C(
        \chs_in_f[0][DATA][26] ), .D(n47), .E(\chs_in_f[1][DATA][26] ), .F(n63), .Z(n97) );
  HS65_LS_OAI212X5 U219 ( .A(n19), .B(n263), .C(n16), .D(n298), .E(n96), .Z(
        \chs_out_f[4][DATA][27] ) );
  HS65_LS_AOI222X2 U220 ( .A(\chs_in_f[2][DATA][27] ), .B(n79), .C(
        \chs_in_f[0][DATA][27] ), .D(n47), .E(\chs_in_f[1][DATA][27] ), .F(n63), .Z(n96) );
  HS65_LS_OAI212X5 U221 ( .A(n19), .B(n262), .C(n16), .D(n297), .E(n95), .Z(
        \chs_out_f[4][DATA][28] ) );
  HS65_LS_AOI222X2 U222 ( .A(\chs_in_f[2][DATA][28] ), .B(n79), .C(
        \chs_in_f[0][DATA][28] ), .D(n47), .E(\chs_in_f[1][DATA][28] ), .F(n63), .Z(n95) );
  HS65_LS_OAI212X5 U223 ( .A(n19), .B(n261), .C(n16), .D(n296), .E(n94), .Z(
        \chs_out_f[4][DATA][29] ) );
  HS65_LS_AOI222X2 U224 ( .A(\chs_in_f[2][DATA][29] ), .B(n79), .C(
        \chs_in_f[0][DATA][29] ), .D(n47), .E(\chs_in_f[1][DATA][29] ), .F(n63), .Z(n94) );
  HS65_LS_OAI212X5 U225 ( .A(n19), .B(n260), .C(n16), .D(n295), .E(n92), .Z(
        \chs_out_f[4][DATA][30] ) );
  HS65_LS_AOI222X2 U226 ( .A(\chs_in_f[2][DATA][30] ), .B(n78), .C(
        \chs_in_f[0][DATA][30] ), .D(n47), .E(\chs_in_f[1][DATA][30] ), .F(n62), .Z(n92) );
  HS65_LS_OAI212X5 U227 ( .A(n20), .B(n259), .C(n16), .D(n294), .E(n91), .Z(
        \chs_out_f[4][DATA][31] ) );
  HS65_LS_AOI222X2 U228 ( .A(\chs_in_f[2][DATA][31] ), .B(n78), .C(
        \chs_in_f[0][DATA][31] ), .D(n48), .E(\chs_in_f[1][DATA][31] ), .F(n62), .Z(n91) );
  HS65_LS_OAI212X5 U229 ( .A(n20), .B(n258), .C(n16), .D(n293), .E(n90), .Z(
        \chs_out_f[4][DATA][32] ) );
  HS65_LS_AOI222X2 U230 ( .A(\chs_in_f[2][DATA][32] ), .B(n78), .C(
        \chs_in_f[0][DATA][32] ), .D(n48), .E(\chs_in_f[1][DATA][32] ), .F(n62), .Z(n90) );
  HS65_LS_OAI212X5 U231 ( .A(n20), .B(n257), .C(n17), .D(n292), .E(n89), .Z(
        \chs_out_f[4][DATA][33] ) );
  HS65_LS_AOI222X2 U232 ( .A(\chs_in_f[2][DATA][33] ), .B(n78), .C(
        \chs_in_f[0][DATA][33] ), .D(n48), .E(\chs_in_f[1][DATA][33] ), .F(n62), .Z(n89) );
  HS65_LS_OAI212X5 U233 ( .A(n281), .B(n23), .C(n316), .D(n8), .E(n151), .Z(
        \chs_out_f[2][DATA][9] ) );
  HS65_LS_AOI222X2 U234 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][9] ), 
        .C(n40), .D(\chs_in_f[0][DATA][9] ), .E(n56), .F(
        \chs_in_f[1][DATA][9] ), .Z(n151) );
  HS65_LS_OAI212X5 U235 ( .A(n281), .B(n26), .C(n316), .D(n11), .E(n186), .Z(
        \chs_out_f[1][DATA][9] ) );
  HS65_LS_AOI222X2 U236 ( .A(n72), .B(\chs_in_f[2][DATA][9] ), .C(n36), .D(
        \chs_in_f[0][DATA][9] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][9] ), .Z(n186) );
  HS65_LS_OAI212X5 U237 ( .A(n281), .B(n29), .C(n316), .D(n14), .E(n221), .Z(
        \chs_out_f[0][DATA][9] ) );
  HS65_LS_AOI222X2 U238 ( .A(n68), .B(\chs_in_f[2][DATA][9] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][9] ), .E(n52), .F(
        \chs_in_f[1][DATA][9] ), .Z(n221) );
  HS65_LS_OAI212X5 U239 ( .A(n290), .B(n21), .C(n325), .D(n6), .E(n185), .Z(
        \chs_out_f[2][DATA][0] ) );
  HS65_LS_AOI222X2 U240 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][0] ), 
        .C(n38), .D(\chs_in_f[0][DATA][0] ), .E(n54), .F(
        \chs_in_f[1][DATA][0] ), .Z(n185) );
  HS65_LS_OAI212X5 U241 ( .A(n289), .B(n21), .C(n324), .D(n6), .E(n174), .Z(
        \chs_out_f[2][DATA][1] ) );
  HS65_LS_AOI222X2 U242 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][1] ), 
        .C(n38), .D(\chs_in_f[0][DATA][1] ), .E(n54), .F(
        \chs_in_f[1][DATA][1] ), .Z(n174) );
  HS65_LS_OAI212X5 U243 ( .A(n288), .B(n22), .C(n323), .D(n7), .E(n163), .Z(
        \chs_out_f[2][DATA][2] ) );
  HS65_LS_AOI222X2 U244 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][2] ), 
        .C(n39), .D(\chs_in_f[0][DATA][2] ), .E(n55), .F(
        \chs_in_f[1][DATA][2] ), .Z(n163) );
  HS65_LS_OAI212X5 U245 ( .A(n280), .B(n21), .C(n315), .D(n6), .E(n184), .Z(
        \chs_out_f[2][DATA][10] ) );
  HS65_LS_AOI222X2 U246 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][10] ), 
        .C(n38), .D(\chs_in_f[0][DATA][10] ), .E(n54), .F(
        \chs_in_f[1][DATA][10] ), .Z(n184) );
  HS65_LS_OAI212X5 U247 ( .A(n279), .B(n21), .C(n314), .D(n6), .E(n183), .Z(
        \chs_out_f[2][DATA][11] ) );
  HS65_LS_AOI222X2 U248 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][11] ), 
        .C(n38), .D(\chs_in_f[0][DATA][11] ), .E(n54), .F(
        \chs_in_f[1][DATA][11] ), .Z(n183) );
  HS65_LS_OAI212X5 U249 ( .A(n278), .B(n21), .C(n313), .D(n6), .E(n182), .Z(
        \chs_out_f[2][DATA][12] ) );
  HS65_LS_AOI222X2 U250 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][12] ), 
        .C(n38), .D(\chs_in_f[0][DATA][12] ), .E(n54), .F(
        \chs_in_f[1][DATA][12] ), .Z(n182) );
  HS65_LS_OAI212X5 U251 ( .A(n277), .B(n21), .C(n312), .D(n6), .E(n181), .Z(
        \chs_out_f[2][DATA][13] ) );
  HS65_LS_AOI222X2 U252 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][13] ), 
        .C(n38), .D(\chs_in_f[0][DATA][13] ), .E(n54), .F(
        \chs_in_f[1][DATA][13] ), .Z(n181) );
  HS65_LS_OAI212X5 U253 ( .A(n276), .B(n21), .C(n311), .D(n6), .E(n180), .Z(
        \chs_out_f[2][DATA][14] ) );
  HS65_LS_AOI222X2 U254 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][14] ), 
        .C(n38), .D(\chs_in_f[0][DATA][14] ), .E(n54), .F(
        \chs_in_f[1][DATA][14] ), .Z(n180) );
  HS65_LS_OAI212X5 U255 ( .A(n275), .B(n21), .C(n310), .D(n6), .E(n179), .Z(
        \chs_out_f[2][DATA][15] ) );
  HS65_LS_AOI222X2 U256 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][15] ), 
        .C(n38), .D(\chs_in_f[0][DATA][15] ), .E(n54), .F(
        \chs_in_f[1][DATA][15] ), .Z(n179) );
  HS65_LS_OAI212X5 U257 ( .A(n274), .B(n21), .C(n309), .D(n6), .E(n178), .Z(
        \chs_out_f[2][DATA][16] ) );
  HS65_LS_AOI222X2 U258 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][16] ), 
        .C(n38), .D(\chs_in_f[0][DATA][16] ), .E(n54), .F(
        \chs_in_f[1][DATA][16] ), .Z(n178) );
  HS65_LS_OAI212X5 U259 ( .A(n273), .B(n21), .C(n308), .D(n6), .E(n177), .Z(
        \chs_out_f[2][DATA][17] ) );
  HS65_LS_AOI222X2 U260 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][17] ), 
        .C(n38), .D(\chs_in_f[0][DATA][17] ), .E(n54), .F(
        \chs_in_f[1][DATA][17] ), .Z(n177) );
  HS65_LS_OAI212X5 U261 ( .A(n272), .B(n21), .C(n307), .D(n6), .E(n176), .Z(
        \chs_out_f[2][DATA][18] ) );
  HS65_LS_AOI222X2 U262 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][18] ), 
        .C(n38), .D(\chs_in_f[0][DATA][18] ), .E(n54), .F(
        \chs_in_f[1][DATA][18] ), .Z(n176) );
  HS65_LS_OAI212X5 U263 ( .A(n271), .B(n21), .C(n306), .D(n6), .E(n175), .Z(
        \chs_out_f[2][DATA][19] ) );
  HS65_LS_AOI222X2 U264 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][19] ), 
        .C(n38), .D(\chs_in_f[0][DATA][19] ), .E(n54), .F(
        \chs_in_f[1][DATA][19] ), .Z(n175) );
  HS65_LS_OAI212X5 U265 ( .A(n270), .B(n21), .C(n305), .D(n7), .E(n173), .Z(
        \chs_out_f[2][DATA][20] ) );
  HS65_LS_AOI222X2 U266 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][20] ), 
        .C(n39), .D(\chs_in_f[0][DATA][20] ), .E(n55), .F(
        \chs_in_f[1][DATA][20] ), .Z(n173) );
  HS65_LS_OAI212X5 U267 ( .A(n269), .B(n22), .C(n304), .D(n7), .E(n172), .Z(
        \chs_out_f[2][DATA][21] ) );
  HS65_LS_AOI222X2 U268 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][21] ), 
        .C(n39), .D(\chs_in_f[0][DATA][21] ), .E(n55), .F(
        \chs_in_f[1][DATA][21] ), .Z(n172) );
  HS65_LS_OAI212X5 U269 ( .A(n268), .B(n22), .C(n303), .D(n7), .E(n171), .Z(
        \chs_out_f[2][DATA][22] ) );
  HS65_LS_AOI222X2 U270 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][22] ), 
        .C(n39), .D(\chs_in_f[0][DATA][22] ), .E(n55), .F(
        \chs_in_f[1][DATA][22] ), .Z(n171) );
  HS65_LS_OAI212X5 U271 ( .A(n267), .B(n22), .C(n302), .D(n7), .E(n170), .Z(
        \chs_out_f[2][DATA][23] ) );
  HS65_LS_AOI222X2 U272 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][23] ), 
        .C(n39), .D(\chs_in_f[0][DATA][23] ), .E(n55), .F(
        \chs_in_f[1][DATA][23] ), .Z(n170) );
  HS65_LS_OAI212X5 U273 ( .A(n266), .B(n22), .C(n301), .D(n7), .E(n169), .Z(
        \chs_out_f[2][DATA][24] ) );
  HS65_LS_AOI222X2 U274 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][24] ), 
        .C(n39), .D(\chs_in_f[0][DATA][24] ), .E(n55), .F(
        \chs_in_f[1][DATA][24] ), .Z(n169) );
  HS65_LS_OAI212X5 U275 ( .A(n265), .B(n22), .C(n300), .D(n7), .E(n168), .Z(
        \chs_out_f[2][DATA][25] ) );
  HS65_LS_AOI222X2 U276 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][25] ), 
        .C(n39), .D(\chs_in_f[0][DATA][25] ), .E(n55), .F(
        \chs_in_f[1][DATA][25] ), .Z(n168) );
  HS65_LS_OAI212X5 U277 ( .A(n264), .B(n22), .C(n299), .D(n7), .E(n167), .Z(
        \chs_out_f[2][DATA][26] ) );
  HS65_LS_AOI222X2 U278 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][26] ), 
        .C(n39), .D(\chs_in_f[0][DATA][26] ), .E(n55), .F(
        \chs_in_f[1][DATA][26] ), .Z(n167) );
  HS65_LS_OAI212X5 U279 ( .A(n263), .B(n22), .C(n298), .D(n7), .E(n166), .Z(
        \chs_out_f[2][DATA][27] ) );
  HS65_LS_AOI222X2 U280 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][27] ), 
        .C(n39), .D(\chs_in_f[0][DATA][27] ), .E(n55), .F(
        \chs_in_f[1][DATA][27] ), .Z(n166) );
  HS65_LS_OAI212X5 U281 ( .A(n262), .B(n22), .C(n297), .D(n7), .E(n165), .Z(
        \chs_out_f[2][DATA][28] ) );
  HS65_LS_AOI222X2 U282 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][28] ), 
        .C(n39), .D(\chs_in_f[0][DATA][28] ), .E(n55), .F(
        \chs_in_f[1][DATA][28] ), .Z(n165) );
  HS65_LS_OAI212X5 U283 ( .A(n261), .B(n22), .C(n296), .D(n7), .E(n164), .Z(
        \chs_out_f[2][DATA][29] ) );
  HS65_LS_AOI222X2 U284 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][29] ), 
        .C(n39), .D(\chs_in_f[0][DATA][29] ), .E(n55), .F(
        \chs_in_f[1][DATA][29] ), .Z(n164) );
  HS65_LS_OAI212X5 U285 ( .A(n260), .B(n22), .C(n295), .D(n7), .E(n162), .Z(
        \chs_out_f[2][DATA][30] ) );
  HS65_LS_AOI222X2 U286 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][30] ), 
        .C(n39), .D(\chs_in_f[0][DATA][30] ), .E(n55), .F(
        \chs_in_f[1][DATA][30] ), .Z(n162) );
  HS65_LS_OAI212X5 U287 ( .A(n259), .B(n22), .C(n294), .D(n8), .E(n161), .Z(
        \chs_out_f[2][DATA][31] ) );
  HS65_LS_AOI222X2 U288 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][31] ), 
        .C(n40), .D(\chs_in_f[0][DATA][31] ), .E(n56), .F(
        \chs_in_f[1][DATA][31] ), .Z(n161) );
  HS65_LS_OAI212X5 U289 ( .A(n258), .B(n22), .C(n293), .D(n8), .E(n160), .Z(
        \chs_out_f[2][DATA][32] ) );
  HS65_LS_AOI222X2 U290 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][32] ), 
        .C(n40), .D(\chs_in_f[0][DATA][32] ), .E(n56), .F(
        \chs_in_f[1][DATA][32] ), .Z(n160) );
  HS65_LS_OAI212X5 U291 ( .A(n290), .B(n24), .C(n325), .D(n9), .E(n220), .Z(
        \chs_out_f[1][DATA][0] ) );
  HS65_LS_AOI222X2 U292 ( .A(n70), .B(\chs_in_f[2][DATA][0] ), .C(n34), .D(
        \chs_in_f[0][DATA][0] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][0] ), .Z(n220) );
  HS65_LS_OAI212X5 U293 ( .A(n289), .B(n24), .C(n324), .D(n9), .E(n209), .Z(
        \chs_out_f[1][DATA][1] ) );
  HS65_LS_AOI222X2 U294 ( .A(n70), .B(\chs_in_f[2][DATA][1] ), .C(n34), .D(
        \chs_in_f[0][DATA][1] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][1] ), .Z(n209) );
  HS65_LS_OAI212X5 U295 ( .A(n288), .B(n25), .C(n323), .D(n10), .E(n198), .Z(
        \chs_out_f[1][DATA][2] ) );
  HS65_LS_AOI222X2 U296 ( .A(n71), .B(\chs_in_f[2][DATA][2] ), .C(n35), .D(
        \chs_in_f[0][DATA][2] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][2] ), .Z(n198) );
  HS65_LS_OAI212X5 U297 ( .A(n280), .B(n24), .C(n315), .D(n9), .E(n219), .Z(
        \chs_out_f[1][DATA][10] ) );
  HS65_LS_AOI222X2 U298 ( .A(n70), .B(\chs_in_f[2][DATA][10] ), .C(n34), .D(
        \chs_in_f[0][DATA][10] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][10] ), .Z(n219) );
  HS65_LS_OAI212X5 U299 ( .A(n279), .B(n24), .C(n314), .D(n9), .E(n218), .Z(
        \chs_out_f[1][DATA][11] ) );
  HS65_LS_AOI222X2 U300 ( .A(n70), .B(\chs_in_f[2][DATA][11] ), .C(n34), .D(
        \chs_in_f[0][DATA][11] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][11] ), .Z(n218) );
  HS65_LS_OAI212X5 U301 ( .A(n278), .B(n24), .C(n313), .D(n9), .E(n217), .Z(
        \chs_out_f[1][DATA][12] ) );
  HS65_LS_AOI222X2 U302 ( .A(n70), .B(\chs_in_f[2][DATA][12] ), .C(n34), .D(
        \chs_in_f[0][DATA][12] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][12] ), .Z(n217) );
  HS65_LS_OAI212X5 U303 ( .A(n277), .B(n24), .C(n312), .D(n9), .E(n216), .Z(
        \chs_out_f[1][DATA][13] ) );
  HS65_LS_AOI222X2 U304 ( .A(n70), .B(\chs_in_f[2][DATA][13] ), .C(n34), .D(
        \chs_in_f[0][DATA][13] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][13] ), .Z(n216) );
  HS65_LS_OAI212X5 U305 ( .A(n276), .B(n24), .C(n311), .D(n9), .E(n215), .Z(
        \chs_out_f[1][DATA][14] ) );
  HS65_LS_AOI222X2 U306 ( .A(n70), .B(\chs_in_f[2][DATA][14] ), .C(n34), .D(
        \chs_in_f[0][DATA][14] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][14] ), .Z(n215) );
  HS65_LS_OAI212X5 U307 ( .A(n275), .B(n24), .C(n310), .D(n9), .E(n214), .Z(
        \chs_out_f[1][DATA][15] ) );
  HS65_LS_AOI222X2 U308 ( .A(n70), .B(\chs_in_f[2][DATA][15] ), .C(n34), .D(
        \chs_in_f[0][DATA][15] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][15] ), .Z(n214) );
  HS65_LS_OAI212X5 U309 ( .A(n274), .B(n24), .C(n309), .D(n9), .E(n213), .Z(
        \chs_out_f[1][DATA][16] ) );
  HS65_LS_AOI222X2 U310 ( .A(n70), .B(\chs_in_f[2][DATA][16] ), .C(n34), .D(
        \chs_in_f[0][DATA][16] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][16] ), .Z(n213) );
  HS65_LS_OAI212X5 U311 ( .A(n273), .B(n24), .C(n308), .D(n9), .E(n212), .Z(
        \chs_out_f[1][DATA][17] ) );
  HS65_LS_AOI222X2 U312 ( .A(n70), .B(\chs_in_f[2][DATA][17] ), .C(n34), .D(
        \chs_in_f[0][DATA][17] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][17] ), .Z(n212) );
  HS65_LS_OAI212X5 U313 ( .A(n272), .B(n24), .C(n307), .D(n9), .E(n211), .Z(
        \chs_out_f[1][DATA][18] ) );
  HS65_LS_AOI222X2 U314 ( .A(n70), .B(\chs_in_f[2][DATA][18] ), .C(n34), .D(
        \chs_in_f[0][DATA][18] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][18] ), .Z(n211) );
  HS65_LS_OAI212X5 U315 ( .A(n271), .B(n24), .C(n306), .D(n9), .E(n210), .Z(
        \chs_out_f[1][DATA][19] ) );
  HS65_LS_AOI222X2 U316 ( .A(n70), .B(\chs_in_f[2][DATA][19] ), .C(n34), .D(
        \chs_in_f[0][DATA][19] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][19] ), .Z(n210) );
  HS65_LS_OAI212X5 U317 ( .A(n270), .B(n24), .C(n305), .D(n10), .E(n208), .Z(
        \chs_out_f[1][DATA][20] ) );
  HS65_LS_AOI222X2 U318 ( .A(n71), .B(\chs_in_f[2][DATA][20] ), .C(n35), .D(
        \chs_in_f[0][DATA][20] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][20] ), .Z(n208) );
  HS65_LS_OAI212X5 U319 ( .A(n269), .B(n25), .C(n304), .D(n10), .E(n207), .Z(
        \chs_out_f[1][DATA][21] ) );
  HS65_LS_AOI222X2 U320 ( .A(n71), .B(\chs_in_f[2][DATA][21] ), .C(n35), .D(
        \chs_in_f[0][DATA][21] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][21] ), .Z(n207) );
  HS65_LS_OAI212X5 U321 ( .A(n268), .B(n25), .C(n303), .D(n10), .E(n206), .Z(
        \chs_out_f[1][DATA][22] ) );
  HS65_LS_AOI222X2 U322 ( .A(n71), .B(\chs_in_f[2][DATA][22] ), .C(n35), .D(
        \chs_in_f[0][DATA][22] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][22] ), .Z(n206) );
  HS65_LS_OAI212X5 U323 ( .A(n267), .B(n25), .C(n302), .D(n10), .E(n205), .Z(
        \chs_out_f[1][DATA][23] ) );
  HS65_LS_AOI222X2 U324 ( .A(n71), .B(\chs_in_f[2][DATA][23] ), .C(n35), .D(
        \chs_in_f[0][DATA][23] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][23] ), .Z(n205) );
  HS65_LS_OAI212X5 U325 ( .A(n266), .B(n25), .C(n301), .D(n10), .E(n204), .Z(
        \chs_out_f[1][DATA][24] ) );
  HS65_LS_AOI222X2 U326 ( .A(n71), .B(\chs_in_f[2][DATA][24] ), .C(n35), .D(
        \chs_in_f[0][DATA][24] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][24] ), .Z(n204) );
  HS65_LS_OAI212X5 U327 ( .A(n265), .B(n25), .C(n300), .D(n10), .E(n203), .Z(
        \chs_out_f[1][DATA][25] ) );
  HS65_LS_AOI222X2 U328 ( .A(n71), .B(\chs_in_f[2][DATA][25] ), .C(n35), .D(
        \chs_in_f[0][DATA][25] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][25] ), .Z(n203) );
  HS65_LS_OAI212X5 U329 ( .A(n264), .B(n25), .C(n299), .D(n10), .E(n202), .Z(
        \chs_out_f[1][DATA][26] ) );
  HS65_LS_AOI222X2 U330 ( .A(n71), .B(\chs_in_f[2][DATA][26] ), .C(n35), .D(
        \chs_in_f[0][DATA][26] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][26] ), .Z(n202) );
  HS65_LS_OAI212X5 U331 ( .A(n263), .B(n25), .C(n298), .D(n10), .E(n201), .Z(
        \chs_out_f[1][DATA][27] ) );
  HS65_LS_AOI222X2 U332 ( .A(n71), .B(\chs_in_f[2][DATA][27] ), .C(n35), .D(
        \chs_in_f[0][DATA][27] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][27] ), .Z(n201) );
  HS65_LS_OAI212X5 U333 ( .A(n262), .B(n25), .C(n297), .D(n10), .E(n200), .Z(
        \chs_out_f[1][DATA][28] ) );
  HS65_LS_AOI222X2 U334 ( .A(n71), .B(\chs_in_f[2][DATA][28] ), .C(n35), .D(
        \chs_in_f[0][DATA][28] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][28] ), .Z(n200) );
  HS65_LS_OAI212X5 U335 ( .A(n261), .B(n25), .C(n296), .D(n10), .E(n199), .Z(
        \chs_out_f[1][DATA][29] ) );
  HS65_LS_AOI222X2 U336 ( .A(n71), .B(\chs_in_f[2][DATA][29] ), .C(n35), .D(
        \chs_in_f[0][DATA][29] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][29] ), .Z(n199) );
  HS65_LS_OAI212X5 U337 ( .A(n260), .B(n25), .C(n295), .D(n10), .E(n197), .Z(
        \chs_out_f[1][DATA][30] ) );
  HS65_LS_AOI222X2 U338 ( .A(n71), .B(\chs_in_f[2][DATA][30] ), .C(n35), .D(
        \chs_in_f[0][DATA][30] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][30] ), .Z(n197) );
  HS65_LS_OAI212X5 U339 ( .A(n259), .B(n25), .C(n294), .D(n11), .E(n196), .Z(
        \chs_out_f[1][DATA][31] ) );
  HS65_LS_AOI222X2 U340 ( .A(n72), .B(\chs_in_f[2][DATA][31] ), .C(n36), .D(
        \chs_in_f[0][DATA][31] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][31] ), .Z(n196) );
  HS65_LS_OAI212X5 U341 ( .A(n258), .B(n25), .C(n293), .D(n11), .E(n195), .Z(
        \chs_out_f[1][DATA][32] ) );
  HS65_LS_AOI222X2 U342 ( .A(n72), .B(\chs_in_f[2][DATA][32] ), .C(n36), .D(
        \chs_in_f[0][DATA][32] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][32] ), .Z(n195) );
  HS65_LS_OAI212X5 U343 ( .A(n290), .B(n27), .C(n325), .D(n12), .E(n255), .Z(
        \chs_out_f[0][DATA][0] ) );
  HS65_LS_AOI222X2 U344 ( .A(n66), .B(\chs_in_f[2][DATA][0] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][0] ), .E(n50), .F(
        \chs_in_f[1][DATA][0] ), .Z(n255) );
  HS65_LS_OAI212X5 U345 ( .A(n289), .B(n27), .C(n324), .D(n12), .E(n244), .Z(
        \chs_out_f[0][DATA][1] ) );
  HS65_LS_AOI222X2 U346 ( .A(n66), .B(\chs_in_f[2][DATA][1] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][1] ), .E(n50), .F(
        \chs_in_f[1][DATA][1] ), .Z(n244) );
  HS65_LS_OAI212X5 U347 ( .A(n288), .B(n28), .C(n323), .D(n13), .E(n233), .Z(
        \chs_out_f[0][DATA][2] ) );
  HS65_LS_AOI222X2 U348 ( .A(n67), .B(\chs_in_f[2][DATA][2] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][2] ), .E(n51), .F(
        \chs_in_f[1][DATA][2] ), .Z(n233) );
  HS65_LS_OAI212X5 U349 ( .A(n280), .B(n27), .C(n315), .D(n12), .E(n254), .Z(
        \chs_out_f[0][DATA][10] ) );
  HS65_LS_AOI222X2 U350 ( .A(n66), .B(\chs_in_f[2][DATA][10] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][10] ), .E(n50), .F(
        \chs_in_f[1][DATA][10] ), .Z(n254) );
  HS65_LS_OAI212X5 U351 ( .A(n279), .B(n27), .C(n314), .D(n12), .E(n253), .Z(
        \chs_out_f[0][DATA][11] ) );
  HS65_LS_AOI222X2 U352 ( .A(n66), .B(\chs_in_f[2][DATA][11] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][11] ), .E(n50), .F(
        \chs_in_f[1][DATA][11] ), .Z(n253) );
  HS65_LS_OAI212X5 U353 ( .A(n278), .B(n27), .C(n313), .D(n12), .E(n252), .Z(
        \chs_out_f[0][DATA][12] ) );
  HS65_LS_AOI222X2 U354 ( .A(n66), .B(\chs_in_f[2][DATA][12] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][12] ), .E(n50), .F(
        \chs_in_f[1][DATA][12] ), .Z(n252) );
  HS65_LS_OAI212X5 U355 ( .A(n277), .B(n27), .C(n312), .D(n12), .E(n251), .Z(
        \chs_out_f[0][DATA][13] ) );
  HS65_LS_AOI222X2 U356 ( .A(n66), .B(\chs_in_f[2][DATA][13] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][13] ), .E(n50), .F(
        \chs_in_f[1][DATA][13] ), .Z(n251) );
  HS65_LS_OAI212X5 U357 ( .A(n276), .B(n27), .C(n311), .D(n12), .E(n250), .Z(
        \chs_out_f[0][DATA][14] ) );
  HS65_LS_AOI222X2 U358 ( .A(n66), .B(\chs_in_f[2][DATA][14] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][14] ), .E(n50), .F(
        \chs_in_f[1][DATA][14] ), .Z(n250) );
  HS65_LS_OAI212X5 U359 ( .A(n275), .B(n27), .C(n310), .D(n12), .E(n249), .Z(
        \chs_out_f[0][DATA][15] ) );
  HS65_LS_AOI222X2 U360 ( .A(n66), .B(\chs_in_f[2][DATA][15] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][15] ), .E(n50), .F(
        \chs_in_f[1][DATA][15] ), .Z(n249) );
  HS65_LS_OAI212X5 U361 ( .A(n274), .B(n27), .C(n309), .D(n12), .E(n248), .Z(
        \chs_out_f[0][DATA][16] ) );
  HS65_LS_AOI222X2 U362 ( .A(n66), .B(\chs_in_f[2][DATA][16] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][16] ), .E(n50), .F(
        \chs_in_f[1][DATA][16] ), .Z(n248) );
  HS65_LS_OAI212X5 U363 ( .A(n273), .B(n27), .C(n308), .D(n12), .E(n247), .Z(
        \chs_out_f[0][DATA][17] ) );
  HS65_LS_AOI222X2 U364 ( .A(n66), .B(\chs_in_f[2][DATA][17] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][17] ), .E(n50), .F(
        \chs_in_f[1][DATA][17] ), .Z(n247) );
  HS65_LS_OAI212X5 U365 ( .A(n272), .B(n27), .C(n307), .D(n12), .E(n246), .Z(
        \chs_out_f[0][DATA][18] ) );
  HS65_LS_AOI222X2 U366 ( .A(n66), .B(\chs_in_f[2][DATA][18] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][18] ), .E(n50), .F(
        \chs_in_f[1][DATA][18] ), .Z(n246) );
  HS65_LS_OAI212X5 U367 ( .A(n271), .B(n27), .C(n306), .D(n12), .E(n245), .Z(
        \chs_out_f[0][DATA][19] ) );
  HS65_LS_AOI222X2 U368 ( .A(n66), .B(\chs_in_f[2][DATA][19] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][19] ), .E(n50), .F(
        \chs_in_f[1][DATA][19] ), .Z(n245) );
  HS65_LS_OAI212X5 U369 ( .A(n270), .B(n27), .C(n305), .D(n13), .E(n243), .Z(
        \chs_out_f[0][DATA][20] ) );
  HS65_LS_AOI222X2 U370 ( .A(n67), .B(\chs_in_f[2][DATA][20] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][20] ), .E(n51), .F(
        \chs_in_f[1][DATA][20] ), .Z(n243) );
  HS65_LS_OAI212X5 U371 ( .A(n269), .B(n28), .C(n304), .D(n13), .E(n242), .Z(
        \chs_out_f[0][DATA][21] ) );
  HS65_LS_AOI222X2 U372 ( .A(n67), .B(\chs_in_f[2][DATA][21] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][21] ), .E(n51), .F(
        \chs_in_f[1][DATA][21] ), .Z(n242) );
  HS65_LS_OAI212X5 U373 ( .A(n268), .B(n28), .C(n303), .D(n13), .E(n241), .Z(
        \chs_out_f[0][DATA][22] ) );
  HS65_LS_AOI222X2 U374 ( .A(n67), .B(\chs_in_f[2][DATA][22] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][22] ), .E(n51), .F(
        \chs_in_f[1][DATA][22] ), .Z(n241) );
  HS65_LS_OAI212X5 U375 ( .A(n267), .B(n28), .C(n302), .D(n13), .E(n240), .Z(
        \chs_out_f[0][DATA][23] ) );
  HS65_LS_AOI222X2 U376 ( .A(n67), .B(\chs_in_f[2][DATA][23] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][23] ), .E(n51), .F(
        \chs_in_f[1][DATA][23] ), .Z(n240) );
  HS65_LS_OAI212X5 U377 ( .A(n266), .B(n28), .C(n301), .D(n13), .E(n239), .Z(
        \chs_out_f[0][DATA][24] ) );
  HS65_LS_AOI222X2 U378 ( .A(n67), .B(\chs_in_f[2][DATA][24] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][24] ), .E(n51), .F(
        \chs_in_f[1][DATA][24] ), .Z(n239) );
  HS65_LS_OAI212X5 U379 ( .A(n265), .B(n28), .C(n300), .D(n13), .E(n238), .Z(
        \chs_out_f[0][DATA][25] ) );
  HS65_LS_AOI222X2 U380 ( .A(n67), .B(\chs_in_f[2][DATA][25] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][25] ), .E(n51), .F(
        \chs_in_f[1][DATA][25] ), .Z(n238) );
  HS65_LS_OAI212X5 U381 ( .A(n264), .B(n28), .C(n299), .D(n13), .E(n237), .Z(
        \chs_out_f[0][DATA][26] ) );
  HS65_LS_AOI222X2 U382 ( .A(n67), .B(\chs_in_f[2][DATA][26] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][26] ), .E(n51), .F(
        \chs_in_f[1][DATA][26] ), .Z(n237) );
  HS65_LS_OAI212X5 U383 ( .A(n263), .B(n28), .C(n298), .D(n13), .E(n236), .Z(
        \chs_out_f[0][DATA][27] ) );
  HS65_LS_AOI222X2 U384 ( .A(n67), .B(\chs_in_f[2][DATA][27] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][27] ), .E(n51), .F(
        \chs_in_f[1][DATA][27] ), .Z(n236) );
  HS65_LS_OAI212X5 U385 ( .A(n262), .B(n28), .C(n297), .D(n13), .E(n235), .Z(
        \chs_out_f[0][DATA][28] ) );
  HS65_LS_AOI222X2 U386 ( .A(n67), .B(\chs_in_f[2][DATA][28] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][28] ), .E(n51), .F(
        \chs_in_f[1][DATA][28] ), .Z(n235) );
  HS65_LS_OAI212X5 U387 ( .A(n261), .B(n28), .C(n296), .D(n13), .E(n234), .Z(
        \chs_out_f[0][DATA][29] ) );
  HS65_LS_AOI222X2 U388 ( .A(n67), .B(\chs_in_f[2][DATA][29] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][29] ), .E(n51), .F(
        \chs_in_f[1][DATA][29] ), .Z(n234) );
  HS65_LS_OAI212X5 U389 ( .A(n260), .B(n28), .C(n295), .D(n13), .E(n232), .Z(
        \chs_out_f[0][DATA][30] ) );
  HS65_LS_AOI222X2 U390 ( .A(n67), .B(\chs_in_f[2][DATA][30] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][30] ), .E(n51), .F(
        \chs_in_f[1][DATA][30] ), .Z(n232) );
  HS65_LS_OAI212X5 U391 ( .A(n259), .B(n28), .C(n294), .D(n14), .E(n231), .Z(
        \chs_out_f[0][DATA][31] ) );
  HS65_LS_AOI222X2 U392 ( .A(n68), .B(\chs_in_f[2][DATA][31] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][31] ), .E(n52), .F(
        \chs_in_f[1][DATA][31] ), .Z(n231) );
  HS65_LS_OAI212X5 U393 ( .A(n258), .B(n28), .C(n293), .D(n14), .E(n230), .Z(
        \chs_out_f[0][DATA][32] ) );
  HS65_LS_AOI222X2 U394 ( .A(n68), .B(\chs_in_f[2][DATA][32] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][32] ), .E(n52), .F(
        \chs_in_f[1][DATA][32] ), .Z(n230) );
  HS65_LS_OAI212X5 U395 ( .A(n287), .B(n23), .C(n322), .D(n8), .E(n157), .Z(
        \chs_out_f[2][DATA][3] ) );
  HS65_LS_AOI222X2 U396 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][3] ), 
        .C(n40), .D(\chs_in_f[0][DATA][3] ), .E(n56), .F(
        \chs_in_f[1][DATA][3] ), .Z(n157) );
  HS65_LS_OAI212X5 U397 ( .A(n286), .B(n23), .C(n321), .D(n8), .E(n156), .Z(
        \chs_out_f[2][DATA][4] ) );
  HS65_LS_AOI222X2 U398 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][4] ), 
        .C(n40), .D(\chs_in_f[0][DATA][4] ), .E(n56), .F(
        \chs_in_f[1][DATA][4] ), .Z(n156) );
  HS65_LS_OAI212X5 U399 ( .A(n285), .B(n23), .C(n320), .D(n8), .E(n155), .Z(
        \chs_out_f[2][DATA][5] ) );
  HS65_LS_AOI222X2 U400 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][5] ), 
        .C(n40), .D(\chs_in_f[0][DATA][5] ), .E(n56), .F(
        \chs_in_f[1][DATA][5] ), .Z(n155) );
  HS65_LS_OAI212X5 U401 ( .A(n284), .B(n23), .C(n319), .D(n8), .E(n154), .Z(
        \chs_out_f[2][DATA][6] ) );
  HS65_LS_AOI222X2 U402 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][6] ), 
        .C(n40), .D(\chs_in_f[0][DATA][6] ), .E(n56), .F(
        \chs_in_f[1][DATA][6] ), .Z(n154) );
  HS65_LS_OAI212X5 U403 ( .A(n283), .B(n23), .C(n318), .D(n8), .E(n153), .Z(
        \chs_out_f[2][DATA][7] ) );
  HS65_LS_AOI222X2 U404 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][7] ), 
        .C(n40), .D(\chs_in_f[0][DATA][7] ), .E(n56), .F(
        \chs_in_f[1][DATA][7] ), .Z(n153) );
  HS65_LS_OAI212X5 U405 ( .A(n282), .B(n23), .C(n317), .D(n8), .E(n152), .Z(
        \chs_out_f[2][DATA][8] ) );
  HS65_LS_AOI222X2 U406 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][8] ), 
        .C(n40), .D(\chs_in_f[0][DATA][8] ), .E(n56), .F(
        \chs_in_f[1][DATA][8] ), .Z(n152) );
  HS65_LS_OAI212X5 U407 ( .A(n257), .B(n23), .C(n292), .D(n8), .E(n159), .Z(
        \chs_out_f[2][DATA][33] ) );
  HS65_LS_AOI222X2 U408 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][33] ), 
        .C(n40), .D(\chs_in_f[0][DATA][33] ), .E(n56), .F(
        \chs_in_f[1][DATA][33] ), .Z(n159) );
  HS65_LS_OAI212X5 U409 ( .A(n287), .B(n26), .C(n322), .D(n11), .E(n192), .Z(
        \chs_out_f[1][DATA][3] ) );
  HS65_LS_AOI222X2 U410 ( .A(n72), .B(\chs_in_f[2][DATA][3] ), .C(n36), .D(
        \chs_in_f[0][DATA][3] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][3] ), .Z(n192) );
  HS65_LS_OAI212X5 U411 ( .A(n286), .B(n26), .C(n321), .D(n11), .E(n191), .Z(
        \chs_out_f[1][DATA][4] ) );
  HS65_LS_AOI222X2 U412 ( .A(n72), .B(\chs_in_f[2][DATA][4] ), .C(n36), .D(
        \chs_in_f[0][DATA][4] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][4] ), .Z(n191) );
  HS65_LS_OAI212X5 U413 ( .A(n285), .B(n26), .C(n320), .D(n11), .E(n190), .Z(
        \chs_out_f[1][DATA][5] ) );
  HS65_LS_AOI222X2 U414 ( .A(n72), .B(\chs_in_f[2][DATA][5] ), .C(n36), .D(
        \chs_in_f[0][DATA][5] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][5] ), .Z(n190) );
  HS65_LS_OAI212X5 U415 ( .A(n284), .B(n26), .C(n319), .D(n11), .E(n189), .Z(
        \chs_out_f[1][DATA][6] ) );
  HS65_LS_AOI222X2 U416 ( .A(n72), .B(\chs_in_f[2][DATA][6] ), .C(n36), .D(
        \chs_in_f[0][DATA][6] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][6] ), .Z(n189) );
  HS65_LS_OAI212X5 U417 ( .A(n283), .B(n26), .C(n318), .D(n11), .E(n188), .Z(
        \chs_out_f[1][DATA][7] ) );
  HS65_LS_AOI222X2 U418 ( .A(n72), .B(\chs_in_f[2][DATA][7] ), .C(n36), .D(
        \chs_in_f[0][DATA][7] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][7] ), .Z(n188) );
  HS65_LS_OAI212X5 U419 ( .A(n282), .B(n26), .C(n317), .D(n11), .E(n187), .Z(
        \chs_out_f[1][DATA][8] ) );
  HS65_LS_AOI222X2 U420 ( .A(n72), .B(\chs_in_f[2][DATA][8] ), .C(n36), .D(
        \chs_in_f[0][DATA][8] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][8] ), .Z(n187) );
  HS65_LS_OAI212X5 U421 ( .A(n257), .B(n26), .C(n292), .D(n11), .E(n194), .Z(
        \chs_out_f[1][DATA][33] ) );
  HS65_LS_AOI222X2 U422 ( .A(n72), .B(\chs_in_f[2][DATA][33] ), .C(n36), .D(
        \chs_in_f[0][DATA][33] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][33] ), .Z(n194) );
  HS65_LS_OAI212X5 U423 ( .A(n287), .B(n29), .C(n322), .D(n14), .E(n227), .Z(
        \chs_out_f[0][DATA][3] ) );
  HS65_LS_AOI222X2 U424 ( .A(n68), .B(\chs_in_f[2][DATA][3] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][3] ), .E(n52), .F(
        \chs_in_f[1][DATA][3] ), .Z(n227) );
  HS65_LS_OAI212X5 U425 ( .A(n286), .B(n29), .C(n321), .D(n14), .E(n226), .Z(
        \chs_out_f[0][DATA][4] ) );
  HS65_LS_AOI222X2 U426 ( .A(n68), .B(\chs_in_f[2][DATA][4] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][4] ), .E(n52), .F(
        \chs_in_f[1][DATA][4] ), .Z(n226) );
  HS65_LS_OAI212X5 U427 ( .A(n285), .B(n29), .C(n320), .D(n14), .E(n225), .Z(
        \chs_out_f[0][DATA][5] ) );
  HS65_LS_AOI222X2 U428 ( .A(n68), .B(\chs_in_f[2][DATA][5] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][5] ), .E(n52), .F(
        \chs_in_f[1][DATA][5] ), .Z(n225) );
  HS65_LS_OAI212X5 U429 ( .A(n284), .B(n29), .C(n319), .D(n14), .E(n224), .Z(
        \chs_out_f[0][DATA][6] ) );
  HS65_LS_AOI222X2 U430 ( .A(n68), .B(\chs_in_f[2][DATA][6] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][6] ), .E(n52), .F(
        \chs_in_f[1][DATA][6] ), .Z(n224) );
  HS65_LS_OAI212X5 U431 ( .A(n283), .B(n29), .C(n318), .D(n14), .E(n223), .Z(
        \chs_out_f[0][DATA][7] ) );
  HS65_LS_AOI222X2 U432 ( .A(n68), .B(\chs_in_f[2][DATA][7] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][7] ), .E(n52), .F(
        \chs_in_f[1][DATA][7] ), .Z(n223) );
  HS65_LS_OAI212X5 U433 ( .A(n282), .B(n29), .C(n317), .D(n14), .E(n222), .Z(
        \chs_out_f[0][DATA][8] ) );
  HS65_LS_AOI222X2 U434 ( .A(n68), .B(\chs_in_f[2][DATA][8] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][8] ), .E(n52), .F(
        \chs_in_f[1][DATA][8] ), .Z(n222) );
  HS65_LS_OAI212X5 U435 ( .A(n257), .B(n29), .C(n292), .D(n14), .E(n229), .Z(
        \chs_out_f[0][DATA][33] ) );
  HS65_LS_AOI222X2 U436 ( .A(n68), .B(\chs_in_f[2][DATA][33] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][33] ), .E(n52), .F(
        \chs_in_f[1][DATA][33] ), .Z(n229) );
  HS65_LS_OAI212X5 U437 ( .A(n281), .B(n32), .C(n316), .D(n5), .E(n116), .Z(
        \chs_out_f[3][DATA][9] ) );
  HS65_LS_AOI222X2 U438 ( .A(n76), .B(\chs_in_f[2][DATA][9] ), .C(n44), .D(
        \chs_in_f[0][DATA][9] ), .E(n60), .F(\chs_in_f[1][DATA][9] ), .Z(n116)
         );
  HS65_LS_OAI212X5 U439 ( .A(n290), .B(n30), .C(n325), .D(n3), .E(n150), .Z(
        \chs_out_f[3][DATA][0] ) );
  HS65_LS_AOI222X2 U440 ( .A(n74), .B(\chs_in_f[2][DATA][0] ), .C(n42), .D(
        \chs_in_f[0][DATA][0] ), .E(n58), .F(\chs_in_f[1][DATA][0] ), .Z(n150)
         );
  HS65_LS_OAI212X5 U441 ( .A(n289), .B(n30), .C(n324), .D(n3), .E(n139), .Z(
        \chs_out_f[3][DATA][1] ) );
  HS65_LS_AOI222X2 U442 ( .A(n74), .B(\chs_in_f[2][DATA][1] ), .C(n42), .D(
        \chs_in_f[0][DATA][1] ), .E(n58), .F(\chs_in_f[1][DATA][1] ), .Z(n139)
         );
  HS65_LS_OAI212X5 U443 ( .A(n288), .B(n31), .C(n323), .D(n4), .E(n128), .Z(
        \chs_out_f[3][DATA][2] ) );
  HS65_LS_AOI222X2 U444 ( .A(n75), .B(\chs_in_f[2][DATA][2] ), .C(n43), .D(
        \chs_in_f[0][DATA][2] ), .E(n59), .F(\chs_in_f[1][DATA][2] ), .Z(n128)
         );
  HS65_LS_OAI212X5 U445 ( .A(n287), .B(n32), .C(n322), .D(n5), .E(n122), .Z(
        \chs_out_f[3][DATA][3] ) );
  HS65_LS_AOI222X2 U446 ( .A(n76), .B(\chs_in_f[2][DATA][3] ), .C(n44), .D(
        \chs_in_f[0][DATA][3] ), .E(n60), .F(\chs_in_f[1][DATA][3] ), .Z(n122)
         );
  HS65_LS_OAI212X5 U447 ( .A(n286), .B(n32), .C(n321), .D(n5), .E(n121), .Z(
        \chs_out_f[3][DATA][4] ) );
  HS65_LS_AOI222X2 U448 ( .A(n76), .B(\chs_in_f[2][DATA][4] ), .C(n44), .D(
        \chs_in_f[0][DATA][4] ), .E(n60), .F(\chs_in_f[1][DATA][4] ), .Z(n121)
         );
  HS65_LS_OAI212X5 U449 ( .A(n285), .B(n32), .C(n320), .D(n5), .E(n120), .Z(
        \chs_out_f[3][DATA][5] ) );
  HS65_LS_AOI222X2 U450 ( .A(n76), .B(\chs_in_f[2][DATA][5] ), .C(n44), .D(
        \chs_in_f[0][DATA][5] ), .E(n60), .F(\chs_in_f[1][DATA][5] ), .Z(n120)
         );
  HS65_LS_OAI212X5 U451 ( .A(n284), .B(n32), .C(n319), .D(n5), .E(n119), .Z(
        \chs_out_f[3][DATA][6] ) );
  HS65_LS_AOI222X2 U452 ( .A(n76), .B(\chs_in_f[2][DATA][6] ), .C(n44), .D(
        \chs_in_f[0][DATA][6] ), .E(n60), .F(\chs_in_f[1][DATA][6] ), .Z(n119)
         );
  HS65_LS_OAI212X5 U453 ( .A(n283), .B(n32), .C(n318), .D(n5), .E(n118), .Z(
        \chs_out_f[3][DATA][7] ) );
  HS65_LS_AOI222X2 U454 ( .A(n76), .B(\chs_in_f[2][DATA][7] ), .C(n44), .D(
        \chs_in_f[0][DATA][7] ), .E(n60), .F(\chs_in_f[1][DATA][7] ), .Z(n118)
         );
  HS65_LS_OAI212X5 U455 ( .A(n282), .B(n32), .C(n317), .D(n5), .E(n117), .Z(
        \chs_out_f[3][DATA][8] ) );
  HS65_LS_AOI222X2 U456 ( .A(n76), .B(\chs_in_f[2][DATA][8] ), .C(n44), .D(
        \chs_in_f[0][DATA][8] ), .E(n60), .F(\chs_in_f[1][DATA][8] ), .Z(n117)
         );
  HS65_LS_OAI212X5 U457 ( .A(n280), .B(n30), .C(n315), .D(n3), .E(n149), .Z(
        \chs_out_f[3][DATA][10] ) );
  HS65_LS_AOI222X2 U458 ( .A(n74), .B(\chs_in_f[2][DATA][10] ), .C(n42), .D(
        \chs_in_f[0][DATA][10] ), .E(n58), .F(\chs_in_f[1][DATA][10] ), .Z(
        n149) );
  HS65_LS_OAI212X5 U459 ( .A(n279), .B(n30), .C(n314), .D(n3), .E(n148), .Z(
        \chs_out_f[3][DATA][11] ) );
  HS65_LS_AOI222X2 U460 ( .A(n74), .B(\chs_in_f[2][DATA][11] ), .C(n42), .D(
        \chs_in_f[0][DATA][11] ), .E(n58), .F(\chs_in_f[1][DATA][11] ), .Z(
        n148) );
  HS65_LS_OAI212X5 U461 ( .A(n278), .B(n30), .C(n313), .D(n3), .E(n147), .Z(
        \chs_out_f[3][DATA][12] ) );
  HS65_LS_AOI222X2 U462 ( .A(n74), .B(\chs_in_f[2][DATA][12] ), .C(n42), .D(
        \chs_in_f[0][DATA][12] ), .E(n58), .F(\chs_in_f[1][DATA][12] ), .Z(
        n147) );
  HS65_LS_OAI212X5 U463 ( .A(n277), .B(n30), .C(n312), .D(n3), .E(n146), .Z(
        \chs_out_f[3][DATA][13] ) );
  HS65_LS_AOI222X2 U464 ( .A(n74), .B(\chs_in_f[2][DATA][13] ), .C(n42), .D(
        \chs_in_f[0][DATA][13] ), .E(n58), .F(\chs_in_f[1][DATA][13] ), .Z(
        n146) );
  HS65_LS_OAI212X5 U465 ( .A(n276), .B(n30), .C(n311), .D(n3), .E(n145), .Z(
        \chs_out_f[3][DATA][14] ) );
  HS65_LS_AOI222X2 U466 ( .A(n74), .B(\chs_in_f[2][DATA][14] ), .C(n42), .D(
        \chs_in_f[0][DATA][14] ), .E(n58), .F(\chs_in_f[1][DATA][14] ), .Z(
        n145) );
  HS65_LS_OAI212X5 U467 ( .A(n275), .B(n30), .C(n310), .D(n3), .E(n144), .Z(
        \chs_out_f[3][DATA][15] ) );
  HS65_LS_AOI222X2 U468 ( .A(n74), .B(\chs_in_f[2][DATA][15] ), .C(n42), .D(
        \chs_in_f[0][DATA][15] ), .E(n58), .F(\chs_in_f[1][DATA][15] ), .Z(
        n144) );
  HS65_LS_OAI212X5 U469 ( .A(n274), .B(n30), .C(n309), .D(n3), .E(n143), .Z(
        \chs_out_f[3][DATA][16] ) );
  HS65_LS_AOI222X2 U470 ( .A(n74), .B(\chs_in_f[2][DATA][16] ), .C(n42), .D(
        \chs_in_f[0][DATA][16] ), .E(n58), .F(\chs_in_f[1][DATA][16] ), .Z(
        n143) );
  HS65_LS_OAI212X5 U471 ( .A(n273), .B(n30), .C(n308), .D(n3), .E(n142), .Z(
        \chs_out_f[3][DATA][17] ) );
  HS65_LS_AOI222X2 U472 ( .A(n74), .B(\chs_in_f[2][DATA][17] ), .C(n42), .D(
        \chs_in_f[0][DATA][17] ), .E(n58), .F(\chs_in_f[1][DATA][17] ), .Z(
        n142) );
  HS65_LS_OAI212X5 U473 ( .A(n272), .B(n30), .C(n307), .D(n3), .E(n141), .Z(
        \chs_out_f[3][DATA][18] ) );
  HS65_LS_AOI222X2 U474 ( .A(n74), .B(\chs_in_f[2][DATA][18] ), .C(n42), .D(
        \chs_in_f[0][DATA][18] ), .E(n58), .F(\chs_in_f[1][DATA][18] ), .Z(
        n141) );
  HS65_LS_OAI212X5 U475 ( .A(n271), .B(n30), .C(n306), .D(n3), .E(n140), .Z(
        \chs_out_f[3][DATA][19] ) );
  HS65_LS_AOI222X2 U476 ( .A(n74), .B(\chs_in_f[2][DATA][19] ), .C(n42), .D(
        \chs_in_f[0][DATA][19] ), .E(n58), .F(\chs_in_f[1][DATA][19] ), .Z(
        n140) );
  HS65_LS_OAI212X5 U477 ( .A(n270), .B(n30), .C(n305), .D(n4), .E(n138), .Z(
        \chs_out_f[3][DATA][20] ) );
  HS65_LS_AOI222X2 U478 ( .A(n75), .B(\chs_in_f[2][DATA][20] ), .C(n43), .D(
        \chs_in_f[0][DATA][20] ), .E(n59), .F(\chs_in_f[1][DATA][20] ), .Z(
        n138) );
  HS65_LS_OAI212X5 U479 ( .A(n269), .B(n31), .C(n304), .D(n4), .E(n137), .Z(
        \chs_out_f[3][DATA][21] ) );
  HS65_LS_AOI222X2 U480 ( .A(n75), .B(\chs_in_f[2][DATA][21] ), .C(n43), .D(
        \chs_in_f[0][DATA][21] ), .E(n59), .F(\chs_in_f[1][DATA][21] ), .Z(
        n137) );
  HS65_LS_OAI212X5 U481 ( .A(n268), .B(n31), .C(n303), .D(n4), .E(n136), .Z(
        \chs_out_f[3][DATA][22] ) );
  HS65_LS_AOI222X2 U482 ( .A(n75), .B(\chs_in_f[2][DATA][22] ), .C(n43), .D(
        \chs_in_f[0][DATA][22] ), .E(n59), .F(\chs_in_f[1][DATA][22] ), .Z(
        n136) );
  HS65_LS_OAI212X5 U483 ( .A(n267), .B(n31), .C(n302), .D(n4), .E(n135), .Z(
        \chs_out_f[3][DATA][23] ) );
  HS65_LS_AOI222X2 U484 ( .A(n75), .B(\chs_in_f[2][DATA][23] ), .C(n43), .D(
        \chs_in_f[0][DATA][23] ), .E(n59), .F(\chs_in_f[1][DATA][23] ), .Z(
        n135) );
  HS65_LS_OAI212X5 U485 ( .A(n266), .B(n31), .C(n301), .D(n4), .E(n134), .Z(
        \chs_out_f[3][DATA][24] ) );
  HS65_LS_AOI222X2 U486 ( .A(n75), .B(\chs_in_f[2][DATA][24] ), .C(n43), .D(
        \chs_in_f[0][DATA][24] ), .E(n59), .F(\chs_in_f[1][DATA][24] ), .Z(
        n134) );
  HS65_LS_OAI212X5 U487 ( .A(n265), .B(n31), .C(n300), .D(n4), .E(n133), .Z(
        \chs_out_f[3][DATA][25] ) );
  HS65_LS_AOI222X2 U488 ( .A(n75), .B(\chs_in_f[2][DATA][25] ), .C(n43), .D(
        \chs_in_f[0][DATA][25] ), .E(n59), .F(\chs_in_f[1][DATA][25] ), .Z(
        n133) );
  HS65_LS_OAI212X5 U489 ( .A(n264), .B(n31), .C(n299), .D(n4), .E(n132), .Z(
        \chs_out_f[3][DATA][26] ) );
  HS65_LS_AOI222X2 U490 ( .A(n75), .B(\chs_in_f[2][DATA][26] ), .C(n43), .D(
        \chs_in_f[0][DATA][26] ), .E(n59), .F(\chs_in_f[1][DATA][26] ), .Z(
        n132) );
  HS65_LS_OAI212X5 U491 ( .A(n263), .B(n31), .C(n298), .D(n4), .E(n131), .Z(
        \chs_out_f[3][DATA][27] ) );
  HS65_LS_AOI222X2 U492 ( .A(n75), .B(\chs_in_f[2][DATA][27] ), .C(n43), .D(
        \chs_in_f[0][DATA][27] ), .E(n59), .F(\chs_in_f[1][DATA][27] ), .Z(
        n131) );
  HS65_LS_OAI212X5 U493 ( .A(n262), .B(n31), .C(n297), .D(n4), .E(n130), .Z(
        \chs_out_f[3][DATA][28] ) );
  HS65_LS_AOI222X2 U494 ( .A(n75), .B(\chs_in_f[2][DATA][28] ), .C(n43), .D(
        \chs_in_f[0][DATA][28] ), .E(n59), .F(\chs_in_f[1][DATA][28] ), .Z(
        n130) );
  HS65_LS_OAI212X5 U495 ( .A(n261), .B(n31), .C(n296), .D(n4), .E(n129), .Z(
        \chs_out_f[3][DATA][29] ) );
  HS65_LS_AOI222X2 U496 ( .A(n75), .B(\chs_in_f[2][DATA][29] ), .C(n43), .D(
        \chs_in_f[0][DATA][29] ), .E(n59), .F(\chs_in_f[1][DATA][29] ), .Z(
        n129) );
  HS65_LS_OAI212X5 U497 ( .A(n260), .B(n31), .C(n295), .D(n4), .E(n127), .Z(
        \chs_out_f[3][DATA][30] ) );
  HS65_LS_AOI222X2 U498 ( .A(n75), .B(\chs_in_f[2][DATA][30] ), .C(n43), .D(
        \chs_in_f[0][DATA][30] ), .E(n59), .F(\chs_in_f[1][DATA][30] ), .Z(
        n127) );
  HS65_LS_OAI212X5 U499 ( .A(n259), .B(n31), .C(n294), .D(n5), .E(n126), .Z(
        \chs_out_f[3][DATA][31] ) );
  HS65_LS_AOI222X2 U500 ( .A(n76), .B(\chs_in_f[2][DATA][31] ), .C(n44), .D(
        \chs_in_f[0][DATA][31] ), .E(n60), .F(\chs_in_f[1][DATA][31] ), .Z(
        n126) );
  HS65_LS_OAI212X5 U501 ( .A(n258), .B(n31), .C(n293), .D(n5), .E(n125), .Z(
        \chs_out_f[3][DATA][32] ) );
  HS65_LS_AOI222X2 U502 ( .A(n76), .B(\chs_in_f[2][DATA][32] ), .C(n44), .D(
        \chs_in_f[0][DATA][32] ), .E(n60), .F(\chs_in_f[1][DATA][32] ), .Z(
        n125) );
  HS65_LS_OAI212X5 U503 ( .A(n257), .B(n32), .C(n292), .D(n5), .E(n124), .Z(
        \chs_out_f[3][DATA][33] ) );
  HS65_LS_AOI222X2 U504 ( .A(n76), .B(\chs_in_f[2][DATA][33] ), .C(n44), .D(
        \chs_in_f[0][DATA][33] ), .E(n60), .F(\chs_in_f[1][DATA][33] ), .Z(
        n124) );
  HS65_LS_OAI212X5 U505 ( .A(n256), .B(n32), .C(n291), .D(n5), .E(n123), .Z(
        \chs_out_f[3][DATA][34] ) );
  HS65_LS_OAI212X5 U506 ( .A(n256), .B(n23), .C(n291), .D(n8), .E(n158), .Z(
        \chs_out_f[2][DATA][34] ) );
  HS65_LS_OAI212X5 U507 ( .A(n256), .B(n26), .C(n291), .D(n11), .E(n193), .Z(
        \chs_out_f[1][DATA][34] ) );
  HS65_LS_OAI212X5 U508 ( .A(n256), .B(n29), .C(n291), .D(n14), .E(n228), .Z(
        \chs_out_f[0][DATA][34] ) );
  HS65_LS_OAI212X5 U509 ( .A(n20), .B(n256), .C(n17), .D(n291), .E(n88), .Z(
        \chs_out_f[4][DATA][34] ) );
  HS65_LS_IVX9 U510 ( .A(\switch_sel[3][3] ), .Z(n335) );
  HS65_LS_IVX9 U511 ( .A(\switch_sel[4][4] ), .Z(n330) );
endmodule


module latch_controller_0_0 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_0_000000000_0 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, n1, n2, n4, n3, n5, n6, n7;
  assign N0 = preset;

  latch_controller_0_0 controller ( .preset(n6), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLQX9 type_out_reg ( .D(N4), .GN(n4), .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U8 ( .A(\left_in[DATA][34] ), .B(n3), .Z(n2) );
  HS65_LS_AND2X4 U7 ( .A(1'b0), .B(n7), .Z(n1) );
  HS65_LS_OR2X9 U9 ( .A(n1), .B(n2), .Z(N4) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(N39), .Q(\right_out[DATA][33] )
         );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(N38), .Q(\right_out[DATA][32] )
         );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(N37), .Q(\right_out[DATA][31] )
         );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(N36), .Q(\right_out[DATA][30] )
         );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(N35), .Q(\right_out[DATA][29] )
         );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(N34), .Q(\right_out[DATA][28] )
         );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(N33), .Q(\right_out[DATA][27] )
         );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(N32), .Q(\right_out[DATA][26] )
         );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(N31), .Q(\right_out[DATA][25] )
         );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(N30), .Q(\right_out[DATA][24] )
         );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(N29), .Q(\right_out[DATA][23] )
         );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(N28), .Q(\right_out[DATA][22] )
         );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(N27), .Q(\right_out[DATA][21] )
         );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(N26), .Q(\right_out[DATA][20] )
         );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(N25), .Q(\right_out[DATA][19] )
         );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(N24), .Q(\right_out[DATA][18] )
         );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(N23), .Q(\right_out[DATA][17] )
         );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(N22), .Q(\right_out[DATA][16] )
         );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(N21), .Q(\right_out[DATA][15] )
         );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(N20), .Q(\right_out[DATA][14] )
         );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(N19), .Q(\right_out[DATA][13] )
         );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(N18), .Q(\right_out[DATA][12] )
         );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(N17), .Q(\right_out[DATA][11] )
         );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(N16), .Q(\right_out[DATA][10] )
         );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(N15), .Q(\right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(N14), .Q(\right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(N13), .Q(\right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(N12), .Q(\right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(N11), .Q(\right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(N10), .Q(\right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(N9), .Q(\right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(N8), .Q(\right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(N7), .Q(\right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(N6), .Q(\right_out[DATA][0] ) );
  HS65_LS_BFX9 U3 ( .A(N0), .Z(n6) );
  HS65_LS_IVX9 U4 ( .A(n6), .Z(n3) );
  HS65_LS_IVX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_NOR2X6 U6 ( .A(lt_enable), .B(n7), .Z(n4) );
  HS65_LS_AND2X4 U10 ( .A(\left_in[DATA][9] ), .B(n3), .Z(N15) );
  HS65_LS_AND2X4 U11 ( .A(\left_in[DATA][0] ), .B(n3), .Z(N6) );
  HS65_LS_AND2X4 U12 ( .A(\left_in[DATA][1] ), .B(n5), .Z(N7) );
  HS65_LS_AND2X4 U13 ( .A(\left_in[DATA][2] ), .B(n3), .Z(N8) );
  HS65_LS_AND2X4 U14 ( .A(\left_in[DATA][3] ), .B(n5), .Z(N9) );
  HS65_LS_AND2X4 U15 ( .A(\left_in[DATA][4] ), .B(n3), .Z(N10) );
  HS65_LS_AND2X4 U16 ( .A(\left_in[DATA][5] ), .B(n3), .Z(N11) );
  HS65_LS_AND2X4 U17 ( .A(\left_in[DATA][6] ), .B(n3), .Z(N12) );
  HS65_LS_AND2X4 U18 ( .A(\left_in[DATA][7] ), .B(n3), .Z(N13) );
  HS65_LS_AND2X4 U19 ( .A(\left_in[DATA][8] ), .B(n3), .Z(N14) );
  HS65_LS_AND2X4 U20 ( .A(\left_in[DATA][10] ), .B(n3), .Z(N16) );
  HS65_LS_AND2X4 U21 ( .A(\left_in[DATA][11] ), .B(n3), .Z(N17) );
  HS65_LS_AND2X4 U22 ( .A(\left_in[DATA][12] ), .B(n3), .Z(N18) );
  HS65_LS_AND2X4 U23 ( .A(\left_in[DATA][13] ), .B(n3), .Z(N19) );
  HS65_LS_AND2X4 U24 ( .A(\left_in[DATA][14] ), .B(n3), .Z(N20) );
  HS65_LS_AND2X4 U25 ( .A(\left_in[DATA][15] ), .B(n3), .Z(N21) );
  HS65_LS_AND2X4 U26 ( .A(\left_in[DATA][16] ), .B(n3), .Z(N22) );
  HS65_LS_AND2X4 U27 ( .A(\left_in[DATA][17] ), .B(n5), .Z(N23) );
  HS65_LS_AND2X4 U28 ( .A(\left_in[DATA][18] ), .B(n5), .Z(N24) );
  HS65_LS_AND2X4 U29 ( .A(\left_in[DATA][19] ), .B(n5), .Z(N25) );
  HS65_LS_AND2X4 U30 ( .A(\left_in[DATA][20] ), .B(n5), .Z(N26) );
  HS65_LS_AND2X4 U31 ( .A(\left_in[DATA][21] ), .B(n5), .Z(N27) );
  HS65_LS_AND2X4 U32 ( .A(\left_in[DATA][22] ), .B(n5), .Z(N28) );
  HS65_LS_AND2X4 U33 ( .A(\left_in[DATA][23] ), .B(n5), .Z(N29) );
  HS65_LS_AND2X4 U34 ( .A(\left_in[DATA][24] ), .B(n5), .Z(N30) );
  HS65_LS_AND2X4 U35 ( .A(\left_in[DATA][25] ), .B(n5), .Z(N31) );
  HS65_LS_AND2X4 U36 ( .A(\left_in[DATA][26] ), .B(n5), .Z(N32) );
  HS65_LS_AND2X4 U37 ( .A(\left_in[DATA][27] ), .B(n5), .Z(N33) );
  HS65_LS_AND2X4 U38 ( .A(\left_in[DATA][28] ), .B(n5), .Z(N34) );
  HS65_LS_AND2X4 U39 ( .A(\left_in[DATA][29] ), .B(n5), .Z(N35) );
  HS65_LS_AND2X4 U40 ( .A(\left_in[DATA][30] ), .B(n3), .Z(N36) );
  HS65_LS_AND2X4 U41 ( .A(\left_in[DATA][31] ), .B(n5), .Z(N37) );
  HS65_LS_AND2X4 U42 ( .A(\left_in[DATA][32] ), .B(n3), .Z(N38) );
  HS65_LS_AND2X4 U43 ( .A(\left_in[DATA][33] ), .B(n5), .Z(N39) );
  HS65_LS_BFX9 U44 ( .A(N0), .Z(n7) );
  HS65_LS_NAND2X7 U45 ( .A(\right_out[DATA][34] ), .B(n4), .Z(N5) );
endmodule


module latch_controller_0_19 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_0_000000000_19 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, n3, n5, n6, n7, n8, n9, n10;
  assign N0 = preset;

  latch_controller_0_19 controller ( .preset(n6), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLQX9 type_out_reg ( .D(N4), .GN(n8), .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(1'b0), .B(n7), .Z(n10) );
  HS65_LS_OR2X9 U9 ( .A(n10), .B(n9), .Z(N4) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(N39), .Q(\right_out[DATA][33] )
         );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(N38), .Q(\right_out[DATA][32] )
         );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(N37), .Q(\right_out[DATA][31] )
         );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(N36), .Q(\right_out[DATA][30] )
         );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(N35), .Q(\right_out[DATA][29] )
         );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(N34), .Q(\right_out[DATA][28] )
         );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(N33), .Q(\right_out[DATA][27] )
         );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(N32), .Q(\right_out[DATA][26] )
         );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(N31), .Q(\right_out[DATA][25] )
         );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(N30), .Q(\right_out[DATA][24] )
         );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(N29), .Q(\right_out[DATA][23] )
         );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(N28), .Q(\right_out[DATA][22] )
         );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(N27), .Q(\right_out[DATA][21] )
         );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(N26), .Q(\right_out[DATA][20] )
         );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(N25), .Q(\right_out[DATA][19] )
         );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(N24), .Q(\right_out[DATA][18] )
         );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(N23), .Q(\right_out[DATA][17] )
         );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(N22), .Q(\right_out[DATA][16] )
         );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(N21), .Q(\right_out[DATA][15] )
         );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(N20), .Q(\right_out[DATA][14] )
         );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(N19), .Q(\right_out[DATA][13] )
         );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(N18), .Q(\right_out[DATA][12] )
         );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(N17), .Q(\right_out[DATA][11] )
         );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(N16), .Q(\right_out[DATA][10] )
         );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(N15), .Q(\right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(N14), .Q(\right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(N13), .Q(\right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(N12), .Q(\right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(N11), .Q(\right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(N10), .Q(\right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(N9), .Q(\right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(N8), .Q(\right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(N7), .Q(\right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(N6), .Q(\right_out[DATA][0] ) );
  HS65_LS_AND2X4 U8 ( .A(\left_in[DATA][34] ), .B(n3), .Z(n9) );
  HS65_LS_AND2X4 U3 ( .A(\left_in[DATA][0] ), .B(n3), .Z(N6) );
  HS65_LS_AND2X4 U4 ( .A(\left_in[DATA][1] ), .B(n5), .Z(N7) );
  HS65_LS_AND2X4 U5 ( .A(\left_in[DATA][2] ), .B(n3), .Z(N8) );
  HS65_LS_AND2X4 U6 ( .A(\left_in[DATA][10] ), .B(n3), .Z(N16) );
  HS65_LS_AND2X4 U10 ( .A(\left_in[DATA][11] ), .B(n3), .Z(N17) );
  HS65_LS_AND2X4 U11 ( .A(\left_in[DATA][12] ), .B(n3), .Z(N18) );
  HS65_LS_AND2X4 U12 ( .A(\left_in[DATA][13] ), .B(n3), .Z(N19) );
  HS65_LS_AND2X4 U13 ( .A(\left_in[DATA][14] ), .B(n3), .Z(N20) );
  HS65_LS_AND2X4 U14 ( .A(\left_in[DATA][15] ), .B(n3), .Z(N21) );
  HS65_LS_AND2X4 U15 ( .A(\left_in[DATA][16] ), .B(n3), .Z(N22) );
  HS65_LS_AND2X4 U16 ( .A(\left_in[DATA][17] ), .B(n5), .Z(N23) );
  HS65_LS_AND2X4 U17 ( .A(\left_in[DATA][18] ), .B(n5), .Z(N24) );
  HS65_LS_AND2X4 U18 ( .A(\left_in[DATA][19] ), .B(n5), .Z(N25) );
  HS65_LS_AND2X4 U19 ( .A(\left_in[DATA][20] ), .B(n5), .Z(N26) );
  HS65_LS_AND2X4 U20 ( .A(\left_in[DATA][21] ), .B(n5), .Z(N27) );
  HS65_LS_AND2X4 U21 ( .A(\left_in[DATA][22] ), .B(n5), .Z(N28) );
  HS65_LS_AND2X4 U22 ( .A(\left_in[DATA][23] ), .B(n5), .Z(N29) );
  HS65_LS_AND2X4 U23 ( .A(\left_in[DATA][24] ), .B(n5), .Z(N30) );
  HS65_LS_AND2X4 U24 ( .A(\left_in[DATA][25] ), .B(n5), .Z(N31) );
  HS65_LS_AND2X4 U25 ( .A(\left_in[DATA][26] ), .B(n5), .Z(N32) );
  HS65_LS_AND2X4 U26 ( .A(\left_in[DATA][27] ), .B(n5), .Z(N33) );
  HS65_LS_AND2X4 U27 ( .A(\left_in[DATA][28] ), .B(n5), .Z(N34) );
  HS65_LS_AND2X4 U28 ( .A(\left_in[DATA][29] ), .B(n5), .Z(N35) );
  HS65_LS_AND2X4 U29 ( .A(\left_in[DATA][30] ), .B(n5), .Z(N36) );
  HS65_LS_AND2X4 U30 ( .A(\left_in[DATA][3] ), .B(n3), .Z(N9) );
  HS65_LS_AND2X4 U31 ( .A(\left_in[DATA][4] ), .B(n3), .Z(N10) );
  HS65_LS_AND2X4 U32 ( .A(\left_in[DATA][5] ), .B(n3), .Z(N11) );
  HS65_LS_AND2X4 U33 ( .A(\left_in[DATA][6] ), .B(n3), .Z(N12) );
  HS65_LS_AND2X4 U34 ( .A(\left_in[DATA][7] ), .B(n3), .Z(N13) );
  HS65_LS_AND2X4 U35 ( .A(\left_in[DATA][8] ), .B(n3), .Z(N14) );
  HS65_LS_AND2X4 U36 ( .A(\left_in[DATA][9] ), .B(n3), .Z(N15) );
  HS65_LS_AND2X4 U37 ( .A(\left_in[DATA][31] ), .B(n5), .Z(N37) );
  HS65_LS_AND2X4 U38 ( .A(\left_in[DATA][32] ), .B(n3), .Z(N38) );
  HS65_LS_AND2X4 U39 ( .A(\left_in[DATA][33] ), .B(n5), .Z(N39) );
  HS65_LS_BFX9 U40 ( .A(N0), .Z(n6) );
  HS65_LS_IVX9 U41 ( .A(n6), .Z(n3) );
  HS65_LS_IVX9 U42 ( .A(n6), .Z(n5) );
  HS65_LS_NOR2X6 U43 ( .A(lt_enable), .B(n7), .Z(n8) );
  HS65_LS_BFX9 U44 ( .A(N0), .Z(n7) );
  HS65_LS_NAND2X7 U45 ( .A(\right_out[DATA][34] ), .B(n8), .Z(N5) );
endmodule


module latch_controller_0_18 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_0_000000000_18 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, n3, n5, n6, n7, n8, n9, n10;
  assign N0 = preset;

  latch_controller_0_18 controller ( .preset(n6), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLQX9 type_out_reg ( .D(N4), .GN(n8), .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U8 ( .A(\left_in[DATA][34] ), .B(n3), .Z(n9) );
  HS65_LS_AND2X4 U7 ( .A(1'b0), .B(n7), .Z(n10) );
  HS65_LS_OR2X9 U9 ( .A(n10), .B(n9), .Z(N4) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(N39), .Q(\right_out[DATA][33] )
         );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(N38), .Q(\right_out[DATA][32] )
         );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(N37), .Q(\right_out[DATA][31] )
         );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(N36), .Q(\right_out[DATA][30] )
         );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(N35), .Q(\right_out[DATA][29] )
         );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(N34), .Q(\right_out[DATA][28] )
         );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(N33), .Q(\right_out[DATA][27] )
         );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(N32), .Q(\right_out[DATA][26] )
         );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(N31), .Q(\right_out[DATA][25] )
         );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(N30), .Q(\right_out[DATA][24] )
         );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(N29), .Q(\right_out[DATA][23] )
         );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(N28), .Q(\right_out[DATA][22] )
         );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(N27), .Q(\right_out[DATA][21] )
         );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(N26), .Q(\right_out[DATA][20] )
         );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(N25), .Q(\right_out[DATA][19] )
         );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(N24), .Q(\right_out[DATA][18] )
         );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(N23), .Q(\right_out[DATA][17] )
         );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(N22), .Q(\right_out[DATA][16] )
         );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(N21), .Q(\right_out[DATA][15] )
         );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(N20), .Q(\right_out[DATA][14] )
         );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(N19), .Q(\right_out[DATA][13] )
         );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(N18), .Q(\right_out[DATA][12] )
         );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(N17), .Q(\right_out[DATA][11] )
         );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(N16), .Q(\right_out[DATA][10] )
         );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(N15), .Q(\right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(N14), .Q(\right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(N13), .Q(\right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(N12), .Q(\right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(N11), .Q(\right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(N10), .Q(\right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(N9), .Q(\right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(N8), .Q(\right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(N7), .Q(\right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(N6), .Q(\right_out[DATA][0] ) );
  HS65_LS_AND2X4 U3 ( .A(\left_in[DATA][0] ), .B(n3), .Z(N6) );
  HS65_LS_AND2X4 U4 ( .A(\left_in[DATA][1] ), .B(n5), .Z(N7) );
  HS65_LS_AND2X4 U5 ( .A(\left_in[DATA][2] ), .B(n3), .Z(N8) );
  HS65_LS_AND2X4 U6 ( .A(\left_in[DATA][10] ), .B(n3), .Z(N16) );
  HS65_LS_AND2X4 U10 ( .A(\left_in[DATA][11] ), .B(n3), .Z(N17) );
  HS65_LS_AND2X4 U11 ( .A(\left_in[DATA][12] ), .B(n3), .Z(N18) );
  HS65_LS_AND2X4 U12 ( .A(\left_in[DATA][13] ), .B(n3), .Z(N19) );
  HS65_LS_AND2X4 U13 ( .A(\left_in[DATA][14] ), .B(n3), .Z(N20) );
  HS65_LS_AND2X4 U14 ( .A(\left_in[DATA][15] ), .B(n3), .Z(N21) );
  HS65_LS_AND2X4 U15 ( .A(\left_in[DATA][16] ), .B(n3), .Z(N22) );
  HS65_LS_AND2X4 U16 ( .A(\left_in[DATA][17] ), .B(n5), .Z(N23) );
  HS65_LS_AND2X4 U17 ( .A(\left_in[DATA][18] ), .B(n5), .Z(N24) );
  HS65_LS_AND2X4 U18 ( .A(\left_in[DATA][19] ), .B(n5), .Z(N25) );
  HS65_LS_AND2X4 U19 ( .A(\left_in[DATA][20] ), .B(n5), .Z(N26) );
  HS65_LS_AND2X4 U20 ( .A(\left_in[DATA][21] ), .B(n5), .Z(N27) );
  HS65_LS_AND2X4 U21 ( .A(\left_in[DATA][22] ), .B(n5), .Z(N28) );
  HS65_LS_AND2X4 U22 ( .A(\left_in[DATA][23] ), .B(n5), .Z(N29) );
  HS65_LS_AND2X4 U23 ( .A(\left_in[DATA][24] ), .B(n5), .Z(N30) );
  HS65_LS_AND2X4 U24 ( .A(\left_in[DATA][25] ), .B(n5), .Z(N31) );
  HS65_LS_AND2X4 U25 ( .A(\left_in[DATA][26] ), .B(n5), .Z(N32) );
  HS65_LS_AND2X4 U26 ( .A(\left_in[DATA][27] ), .B(n5), .Z(N33) );
  HS65_LS_AND2X4 U27 ( .A(\left_in[DATA][28] ), .B(n5), .Z(N34) );
  HS65_LS_AND2X4 U28 ( .A(\left_in[DATA][29] ), .B(n5), .Z(N35) );
  HS65_LS_AND2X4 U29 ( .A(\left_in[DATA][30] ), .B(n5), .Z(N36) );
  HS65_LS_AND2X4 U30 ( .A(\left_in[DATA][31] ), .B(n3), .Z(N37) );
  HS65_LS_AND2X4 U31 ( .A(\left_in[DATA][32] ), .B(n5), .Z(N38) );
  HS65_LS_AND2X4 U32 ( .A(\left_in[DATA][4] ), .B(n3), .Z(N10) );
  HS65_LS_AND2X4 U33 ( .A(\left_in[DATA][5] ), .B(n3), .Z(N11) );
  HS65_LS_AND2X4 U34 ( .A(\left_in[DATA][6] ), .B(n3), .Z(N12) );
  HS65_LS_AND2X4 U35 ( .A(\left_in[DATA][7] ), .B(n3), .Z(N13) );
  HS65_LS_AND2X4 U36 ( .A(\left_in[DATA][8] ), .B(n3), .Z(N14) );
  HS65_LS_AND2X4 U37 ( .A(\left_in[DATA][9] ), .B(n3), .Z(N15) );
  HS65_LS_AND2X4 U38 ( .A(\left_in[DATA][3] ), .B(n3), .Z(N9) );
  HS65_LS_AND2X4 U39 ( .A(\left_in[DATA][33] ), .B(n5), .Z(N39) );
  HS65_LS_BFX9 U40 ( .A(N0), .Z(n6) );
  HS65_LS_IVX9 U41 ( .A(n6), .Z(n3) );
  HS65_LS_IVX9 U42 ( .A(n6), .Z(n5) );
  HS65_LS_NOR2X6 U43 ( .A(lt_enable), .B(n7), .Z(n8) );
  HS65_LS_BFX9 U44 ( .A(N0), .Z(n7) );
  HS65_LS_NAND2X7 U45 ( .A(\right_out[DATA][34] ), .B(n8), .Z(N5) );
endmodule


module latch_controller_0_17 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_0_000000000_17 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, n3, n5, n6, n7, n8, n9, n10;
  assign N0 = preset;

  latch_controller_0_17 controller ( .preset(n6), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLQX9 type_out_reg ( .D(N4), .GN(n8), .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U8 ( .A(\left_in[DATA][34] ), .B(n3), .Z(n9) );
  HS65_LS_AND2X4 U7 ( .A(1'b0), .B(n7), .Z(n10) );
  HS65_LS_OR2X9 U9 ( .A(n10), .B(n9), .Z(N4) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(N39), .Q(\right_out[DATA][33] )
         );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(N38), .Q(\right_out[DATA][32] )
         );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(N37), .Q(\right_out[DATA][31] )
         );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(N36), .Q(\right_out[DATA][30] )
         );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(N35), .Q(\right_out[DATA][29] )
         );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(N34), .Q(\right_out[DATA][28] )
         );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(N33), .Q(\right_out[DATA][27] )
         );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(N32), .Q(\right_out[DATA][26] )
         );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(N31), .Q(\right_out[DATA][25] )
         );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(N30), .Q(\right_out[DATA][24] )
         );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(N29), .Q(\right_out[DATA][23] )
         );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(N28), .Q(\right_out[DATA][22] )
         );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(N27), .Q(\right_out[DATA][21] )
         );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(N26), .Q(\right_out[DATA][20] )
         );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(N25), .Q(\right_out[DATA][19] )
         );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(N24), .Q(\right_out[DATA][18] )
         );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(N23), .Q(\right_out[DATA][17] )
         );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(N22), .Q(\right_out[DATA][16] )
         );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(N21), .Q(\right_out[DATA][15] )
         );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(N20), .Q(\right_out[DATA][14] )
         );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(N19), .Q(\right_out[DATA][13] )
         );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(N18), .Q(\right_out[DATA][12] )
         );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(N17), .Q(\right_out[DATA][11] )
         );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(N16), .Q(\right_out[DATA][10] )
         );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(N15), .Q(\right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(N14), .Q(\right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(N13), .Q(\right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(N12), .Q(\right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(N11), .Q(\right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(N10), .Q(\right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(N9), .Q(\right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(N8), .Q(\right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(N7), .Q(\right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(N6), .Q(\right_out[DATA][0] ) );
  HS65_LS_AND2X4 U3 ( .A(\left_in[DATA][0] ), .B(n3), .Z(N6) );
  HS65_LS_AND2X4 U4 ( .A(\left_in[DATA][1] ), .B(n5), .Z(N7) );
  HS65_LS_AND2X4 U5 ( .A(\left_in[DATA][2] ), .B(n3), .Z(N8) );
  HS65_LS_AND2X4 U6 ( .A(\left_in[DATA][10] ), .B(n3), .Z(N16) );
  HS65_LS_AND2X4 U10 ( .A(\left_in[DATA][11] ), .B(n3), .Z(N17) );
  HS65_LS_AND2X4 U11 ( .A(\left_in[DATA][12] ), .B(n3), .Z(N18) );
  HS65_LS_AND2X4 U12 ( .A(\left_in[DATA][13] ), .B(n3), .Z(N19) );
  HS65_LS_AND2X4 U13 ( .A(\left_in[DATA][14] ), .B(n3), .Z(N20) );
  HS65_LS_AND2X4 U14 ( .A(\left_in[DATA][15] ), .B(n3), .Z(N21) );
  HS65_LS_AND2X4 U15 ( .A(\left_in[DATA][16] ), .B(n3), .Z(N22) );
  HS65_LS_AND2X4 U16 ( .A(\left_in[DATA][17] ), .B(n5), .Z(N23) );
  HS65_LS_AND2X4 U17 ( .A(\left_in[DATA][18] ), .B(n5), .Z(N24) );
  HS65_LS_AND2X4 U18 ( .A(\left_in[DATA][19] ), .B(n5), .Z(N25) );
  HS65_LS_AND2X4 U19 ( .A(\left_in[DATA][20] ), .B(n5), .Z(N26) );
  HS65_LS_AND2X4 U20 ( .A(\left_in[DATA][21] ), .B(n5), .Z(N27) );
  HS65_LS_AND2X4 U21 ( .A(\left_in[DATA][22] ), .B(n5), .Z(N28) );
  HS65_LS_AND2X4 U22 ( .A(\left_in[DATA][23] ), .B(n5), .Z(N29) );
  HS65_LS_AND2X4 U23 ( .A(\left_in[DATA][24] ), .B(n5), .Z(N30) );
  HS65_LS_AND2X4 U24 ( .A(\left_in[DATA][25] ), .B(n5), .Z(N31) );
  HS65_LS_AND2X4 U25 ( .A(\left_in[DATA][26] ), .B(n5), .Z(N32) );
  HS65_LS_AND2X4 U26 ( .A(\left_in[DATA][27] ), .B(n5), .Z(N33) );
  HS65_LS_AND2X4 U27 ( .A(\left_in[DATA][28] ), .B(n5), .Z(N34) );
  HS65_LS_AND2X4 U28 ( .A(\left_in[DATA][29] ), .B(n5), .Z(N35) );
  HS65_LS_AND2X4 U29 ( .A(\left_in[DATA][30] ), .B(n5), .Z(N36) );
  HS65_LS_AND2X4 U30 ( .A(\left_in[DATA][31] ), .B(n3), .Z(N37) );
  HS65_LS_AND2X4 U31 ( .A(\left_in[DATA][32] ), .B(n5), .Z(N38) );
  HS65_LS_AND2X4 U32 ( .A(\left_in[DATA][4] ), .B(n3), .Z(N10) );
  HS65_LS_AND2X4 U33 ( .A(\left_in[DATA][5] ), .B(n3), .Z(N11) );
  HS65_LS_AND2X4 U34 ( .A(\left_in[DATA][6] ), .B(n3), .Z(N12) );
  HS65_LS_AND2X4 U35 ( .A(\left_in[DATA][7] ), .B(n3), .Z(N13) );
  HS65_LS_AND2X4 U36 ( .A(\left_in[DATA][8] ), .B(n3), .Z(N14) );
  HS65_LS_AND2X4 U37 ( .A(\left_in[DATA][9] ), .B(n3), .Z(N15) );
  HS65_LS_AND2X4 U38 ( .A(\left_in[DATA][3] ), .B(n3), .Z(N9) );
  HS65_LS_AND2X4 U39 ( .A(\left_in[DATA][33] ), .B(n5), .Z(N39) );
  HS65_LS_BFX9 U40 ( .A(N0), .Z(n6) );
  HS65_LS_IVX9 U41 ( .A(n6), .Z(n3) );
  HS65_LS_IVX9 U42 ( .A(n6), .Z(n5) );
  HS65_LS_NOR2X6 U43 ( .A(lt_enable), .B(n7), .Z(n8) );
  HS65_LS_BFX9 U44 ( .A(N0), .Z(n7) );
  HS65_LS_NAND2X7 U45 ( .A(\right_out[DATA][34] ), .B(n8), .Z(N5) );
endmodule


module latch_controller_0_16 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_0_000000000_16 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, n3, n5, n6, n7, n8, n9, n10;
  assign N0 = preset;

  latch_controller_0_16 controller ( .preset(n6), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLQX9 type_out_reg ( .D(N4), .GN(n8), .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U8 ( .A(\left_in[DATA][34] ), .B(n3), .Z(n9) );
  HS65_LS_AND2X4 U7 ( .A(1'b0), .B(n7), .Z(n10) );
  HS65_LS_OR2X9 U9 ( .A(n10), .B(n9), .Z(N4) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(N39), .Q(\right_out[DATA][33] )
         );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(N38), .Q(\right_out[DATA][32] )
         );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(N37), .Q(\right_out[DATA][31] )
         );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(N36), .Q(\right_out[DATA][30] )
         );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(N35), .Q(\right_out[DATA][29] )
         );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(N34), .Q(\right_out[DATA][28] )
         );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(N33), .Q(\right_out[DATA][27] )
         );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(N32), .Q(\right_out[DATA][26] )
         );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(N31), .Q(\right_out[DATA][25] )
         );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(N30), .Q(\right_out[DATA][24] )
         );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(N29), .Q(\right_out[DATA][23] )
         );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(N28), .Q(\right_out[DATA][22] )
         );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(N27), .Q(\right_out[DATA][21] )
         );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(N26), .Q(\right_out[DATA][20] )
         );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(N25), .Q(\right_out[DATA][19] )
         );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(N24), .Q(\right_out[DATA][18] )
         );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(N23), .Q(\right_out[DATA][17] )
         );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(N22), .Q(\right_out[DATA][16] )
         );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(N21), .Q(\right_out[DATA][15] )
         );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(N20), .Q(\right_out[DATA][14] )
         );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(N19), .Q(\right_out[DATA][13] )
         );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(N18), .Q(\right_out[DATA][12] )
         );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(N17), .Q(\right_out[DATA][11] )
         );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(N16), .Q(\right_out[DATA][10] )
         );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(N15), .Q(\right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(N14), .Q(\right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(N13), .Q(\right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(N12), .Q(\right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(N11), .Q(\right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(N10), .Q(\right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(N9), .Q(\right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(N8), .Q(\right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(N7), .Q(\right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(N6), .Q(\right_out[DATA][0] ) );
  HS65_LS_AND2X4 U3 ( .A(\left_in[DATA][16] ), .B(n3), .Z(N22) );
  HS65_LS_AND2X4 U4 ( .A(\left_in[DATA][17] ), .B(n5), .Z(N23) );
  HS65_LS_AND2X4 U5 ( .A(\left_in[DATA][18] ), .B(n5), .Z(N24) );
  HS65_LS_AND2X4 U6 ( .A(\left_in[DATA][19] ), .B(n5), .Z(N25) );
  HS65_LS_AND2X4 U10 ( .A(\left_in[DATA][20] ), .B(n5), .Z(N26) );
  HS65_LS_AND2X4 U11 ( .A(\left_in[DATA][21] ), .B(n5), .Z(N27) );
  HS65_LS_AND2X4 U12 ( .A(\left_in[DATA][22] ), .B(n5), .Z(N28) );
  HS65_LS_AND2X4 U13 ( .A(\left_in[DATA][23] ), .B(n5), .Z(N29) );
  HS65_LS_AND2X4 U14 ( .A(\left_in[DATA][24] ), .B(n5), .Z(N30) );
  HS65_LS_AND2X4 U15 ( .A(\left_in[DATA][25] ), .B(n5), .Z(N31) );
  HS65_LS_AND2X4 U16 ( .A(\left_in[DATA][26] ), .B(n5), .Z(N32) );
  HS65_LS_AND2X4 U17 ( .A(\left_in[DATA][27] ), .B(n5), .Z(N33) );
  HS65_LS_AND2X4 U18 ( .A(\left_in[DATA][28] ), .B(n5), .Z(N34) );
  HS65_LS_AND2X4 U19 ( .A(\left_in[DATA][29] ), .B(n5), .Z(N35) );
  HS65_LS_AND2X4 U20 ( .A(\left_in[DATA][4] ), .B(n3), .Z(N10) );
  HS65_LS_AND2X4 U21 ( .A(\left_in[DATA][5] ), .B(n3), .Z(N11) );
  HS65_LS_AND2X4 U22 ( .A(\left_in[DATA][6] ), .B(n3), .Z(N12) );
  HS65_LS_AND2X4 U23 ( .A(\left_in[DATA][7] ), .B(n3), .Z(N13) );
  HS65_LS_AND2X4 U24 ( .A(\left_in[DATA][8] ), .B(n3), .Z(N14) );
  HS65_LS_AND2X4 U25 ( .A(\left_in[DATA][9] ), .B(n3), .Z(N15) );
  HS65_LS_AND2X4 U26 ( .A(\left_in[DATA][10] ), .B(n3), .Z(N16) );
  HS65_LS_AND2X4 U27 ( .A(\left_in[DATA][11] ), .B(n3), .Z(N17) );
  HS65_LS_AND2X4 U28 ( .A(\left_in[DATA][12] ), .B(n3), .Z(N18) );
  HS65_LS_AND2X4 U29 ( .A(\left_in[DATA][13] ), .B(n3), .Z(N19) );
  HS65_LS_AND2X4 U30 ( .A(\left_in[DATA][14] ), .B(n3), .Z(N20) );
  HS65_LS_AND2X4 U31 ( .A(\left_in[DATA][15] ), .B(n3), .Z(N21) );
  HS65_LS_AND2X4 U32 ( .A(\left_in[DATA][30] ), .B(n3), .Z(N36) );
  HS65_LS_AND2X4 U33 ( .A(\left_in[DATA][31] ), .B(n5), .Z(N37) );
  HS65_LS_AND2X4 U34 ( .A(\left_in[DATA][32] ), .B(n3), .Z(N38) );
  HS65_LS_AND2X4 U35 ( .A(\left_in[DATA][33] ), .B(n5), .Z(N39) );
  HS65_LS_AND2X4 U36 ( .A(\left_in[DATA][0] ), .B(n3), .Z(N6) );
  HS65_LS_AND2X4 U37 ( .A(\left_in[DATA][1] ), .B(n5), .Z(N7) );
  HS65_LS_AND2X4 U38 ( .A(\left_in[DATA][2] ), .B(n3), .Z(N8) );
  HS65_LS_AND2X4 U39 ( .A(\left_in[DATA][3] ), .B(n5), .Z(N9) );
  HS65_LS_BFX9 U40 ( .A(N0), .Z(n6) );
  HS65_LS_IVX9 U41 ( .A(n6), .Z(n3) );
  HS65_LS_IVX9 U42 ( .A(n6), .Z(n5) );
  HS65_LS_NOR2X6 U43 ( .A(lt_enable), .B(n7), .Z(n8) );
  HS65_LS_BFX9 U44 ( .A(N0), .Z(n7) );
  HS65_LS_NAND2X7 U45 ( .A(\right_out[DATA][34] ), .B(n8), .Z(N5) );
endmodule


module crossbar_stage_0 ( preset, .switch_sel({\switch_sel[4][4] , 
        \switch_sel[4][3] , \switch_sel[4][2] , \switch_sel[4][1] , 
        \switch_sel[4][0] , \switch_sel[3][4] , \switch_sel[3][3] , 
        \switch_sel[3][2] , \switch_sel[3][1] , \switch_sel[3][0] , 
        \switch_sel[2][4] , \switch_sel[2][3] , \switch_sel[2][2] , 
        \switch_sel[2][1] , \switch_sel[2][0] , \switch_sel[1][4] , 
        \switch_sel[1][3] , \switch_sel[1][2] , \switch_sel[1][1] , 
        \switch_sel[1][0] , \switch_sel[0][4] , \switch_sel[0][3] , 
        \switch_sel[0][2] , \switch_sel[0][1] , \switch_sel[0][0] }), 
    .chs_in_f({\chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] , 
        \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] , 
        \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] , 
        \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] , 
        \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] , 
        \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] , 
        \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] , 
        \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] , 
        \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] , 
        \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] , 
        \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] , 
        \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] , 
        \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] , 
        \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] , \chs_in_f[4][DATA][7] , 
        \chs_in_f[4][DATA][6] , \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] , 
        \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] , \chs_in_f[4][DATA][1] , 
        \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] , \chs_in_f[3][DATA][34] , 
        \chs_in_f[3][DATA][33] , \chs_in_f[3][DATA][32] , 
        \chs_in_f[3][DATA][31] , \chs_in_f[3][DATA][30] , 
        \chs_in_f[3][DATA][29] , \chs_in_f[3][DATA][28] , 
        \chs_in_f[3][DATA][27] , \chs_in_f[3][DATA][26] , 
        \chs_in_f[3][DATA][25] , \chs_in_f[3][DATA][24] , 
        \chs_in_f[3][DATA][23] , \chs_in_f[3][DATA][22] , 
        \chs_in_f[3][DATA][21] , \chs_in_f[3][DATA][20] , 
        \chs_in_f[3][DATA][19] , \chs_in_f[3][DATA][18] , 
        \chs_in_f[3][DATA][17] , \chs_in_f[3][DATA][16] , 
        \chs_in_f[3][DATA][15] , \chs_in_f[3][DATA][14] , 
        \chs_in_f[3][DATA][13] , \chs_in_f[3][DATA][12] , 
        \chs_in_f[3][DATA][11] , \chs_in_f[3][DATA][10] , 
        \chs_in_f[3][DATA][9] , \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] , 
        \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] , \chs_in_f[3][DATA][4] , 
        \chs_in_f[3][DATA][3] , \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] , 
        \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] , 
        \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] , 
        \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] , 
        \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] , 
        \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] , 
        \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] , 
        \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] , 
        \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] , 
        \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] , 
        \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] , 
        \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] , 
        \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] , 
        \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] , 
        \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] , \chs_in_f[2][DATA][7] , 
        \chs_in_f[2][DATA][6] , \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] , 
        \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] , \chs_in_f[2][DATA][1] , 
        \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] , \chs_in_f[1][DATA][34] , 
        \chs_in_f[1][DATA][33] , \chs_in_f[1][DATA][32] , 
        \chs_in_f[1][DATA][31] , \chs_in_f[1][DATA][30] , 
        \chs_in_f[1][DATA][29] , \chs_in_f[1][DATA][28] , 
        \chs_in_f[1][DATA][27] , \chs_in_f[1][DATA][26] , 
        \chs_in_f[1][DATA][25] , \chs_in_f[1][DATA][24] , 
        \chs_in_f[1][DATA][23] , \chs_in_f[1][DATA][22] , 
        \chs_in_f[1][DATA][21] , \chs_in_f[1][DATA][20] , 
        \chs_in_f[1][DATA][19] , \chs_in_f[1][DATA][18] , 
        \chs_in_f[1][DATA][17] , \chs_in_f[1][DATA][16] , 
        \chs_in_f[1][DATA][15] , \chs_in_f[1][DATA][14] , 
        \chs_in_f[1][DATA][13] , \chs_in_f[1][DATA][12] , 
        \chs_in_f[1][DATA][11] , \chs_in_f[1][DATA][10] , 
        \chs_in_f[1][DATA][9] , \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] , 
        \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] , \chs_in_f[1][DATA][4] , 
        \chs_in_f[1][DATA][3] , \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] , 
        \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] , 
        \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] , 
        \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] , 
        \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] , 
        \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] , 
        \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] , 
        \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] , 
        \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] , 
        \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] , 
        \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] , 
        \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] , 
        \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] , 
        \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] , 
        \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] , \chs_in_f[0][DATA][7] , 
        \chs_in_f[0][DATA][6] , \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] , 
        \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] , \chs_in_f[0][DATA][1] , 
        \chs_in_f[0][DATA][0] }), .chs_in_b({\chs_in_b[4][ACK] , 
        \chs_in_b[3][ACK] , \chs_in_b[2][ACK] , \chs_in_b[1][ACK] , 
        \chs_in_b[0][ACK] }), .latches_out_f({\latches_out_f[4][REQ] , 
        \latches_out_f[4][DATA][34] , \latches_out_f[4][DATA][33] , 
        \latches_out_f[4][DATA][32] , \latches_out_f[4][DATA][31] , 
        \latches_out_f[4][DATA][30] , \latches_out_f[4][DATA][29] , 
        \latches_out_f[4][DATA][28] , \latches_out_f[4][DATA][27] , 
        \latches_out_f[4][DATA][26] , \latches_out_f[4][DATA][25] , 
        \latches_out_f[4][DATA][24] , \latches_out_f[4][DATA][23] , 
        \latches_out_f[4][DATA][22] , \latches_out_f[4][DATA][21] , 
        \latches_out_f[4][DATA][20] , \latches_out_f[4][DATA][19] , 
        \latches_out_f[4][DATA][18] , \latches_out_f[4][DATA][17] , 
        \latches_out_f[4][DATA][16] , \latches_out_f[4][DATA][15] , 
        \latches_out_f[4][DATA][14] , \latches_out_f[4][DATA][13] , 
        \latches_out_f[4][DATA][12] , \latches_out_f[4][DATA][11] , 
        \latches_out_f[4][DATA][10] , \latches_out_f[4][DATA][9] , 
        \latches_out_f[4][DATA][8] , \latches_out_f[4][DATA][7] , 
        \latches_out_f[4][DATA][6] , \latches_out_f[4][DATA][5] , 
        \latches_out_f[4][DATA][4] , \latches_out_f[4][DATA][3] , 
        \latches_out_f[4][DATA][2] , \latches_out_f[4][DATA][1] , 
        \latches_out_f[4][DATA][0] , \latches_out_f[3][REQ] , 
        \latches_out_f[3][DATA][34] , \latches_out_f[3][DATA][33] , 
        \latches_out_f[3][DATA][32] , \latches_out_f[3][DATA][31] , 
        \latches_out_f[3][DATA][30] , \latches_out_f[3][DATA][29] , 
        \latches_out_f[3][DATA][28] , \latches_out_f[3][DATA][27] , 
        \latches_out_f[3][DATA][26] , \latches_out_f[3][DATA][25] , 
        \latches_out_f[3][DATA][24] , \latches_out_f[3][DATA][23] , 
        \latches_out_f[3][DATA][22] , \latches_out_f[3][DATA][21] , 
        \latches_out_f[3][DATA][20] , \latches_out_f[3][DATA][19] , 
        \latches_out_f[3][DATA][18] , \latches_out_f[3][DATA][17] , 
        \latches_out_f[3][DATA][16] , \latches_out_f[3][DATA][15] , 
        \latches_out_f[3][DATA][14] , \latches_out_f[3][DATA][13] , 
        \latches_out_f[3][DATA][12] , \latches_out_f[3][DATA][11] , 
        \latches_out_f[3][DATA][10] , \latches_out_f[3][DATA][9] , 
        \latches_out_f[3][DATA][8] , \latches_out_f[3][DATA][7] , 
        \latches_out_f[3][DATA][6] , \latches_out_f[3][DATA][5] , 
        \latches_out_f[3][DATA][4] , \latches_out_f[3][DATA][3] , 
        \latches_out_f[3][DATA][2] , \latches_out_f[3][DATA][1] , 
        \latches_out_f[3][DATA][0] , \latches_out_f[2][REQ] , 
        \latches_out_f[2][DATA][34] , \latches_out_f[2][DATA][33] , 
        \latches_out_f[2][DATA][32] , \latches_out_f[2][DATA][31] , 
        \latches_out_f[2][DATA][30] , \latches_out_f[2][DATA][29] , 
        \latches_out_f[2][DATA][28] , \latches_out_f[2][DATA][27] , 
        \latches_out_f[2][DATA][26] , \latches_out_f[2][DATA][25] , 
        \latches_out_f[2][DATA][24] , \latches_out_f[2][DATA][23] , 
        \latches_out_f[2][DATA][22] , \latches_out_f[2][DATA][21] , 
        \latches_out_f[2][DATA][20] , \latches_out_f[2][DATA][19] , 
        \latches_out_f[2][DATA][18] , \latches_out_f[2][DATA][17] , 
        \latches_out_f[2][DATA][16] , \latches_out_f[2][DATA][15] , 
        \latches_out_f[2][DATA][14] , \latches_out_f[2][DATA][13] , 
        \latches_out_f[2][DATA][12] , \latches_out_f[2][DATA][11] , 
        \latches_out_f[2][DATA][10] , \latches_out_f[2][DATA][9] , 
        \latches_out_f[2][DATA][8] , \latches_out_f[2][DATA][7] , 
        \latches_out_f[2][DATA][6] , \latches_out_f[2][DATA][5] , 
        \latches_out_f[2][DATA][4] , \latches_out_f[2][DATA][3] , 
        \latches_out_f[2][DATA][2] , \latches_out_f[2][DATA][1] , 
        \latches_out_f[2][DATA][0] , \latches_out_f[1][REQ] , 
        \latches_out_f[1][DATA][34] , \latches_out_f[1][DATA][33] , 
        \latches_out_f[1][DATA][32] , \latches_out_f[1][DATA][31] , 
        \latches_out_f[1][DATA][30] , \latches_out_f[1][DATA][29] , 
        \latches_out_f[1][DATA][28] , \latches_out_f[1][DATA][27] , 
        \latches_out_f[1][DATA][26] , \latches_out_f[1][DATA][25] , 
        \latches_out_f[1][DATA][24] , \latches_out_f[1][DATA][23] , 
        \latches_out_f[1][DATA][22] , \latches_out_f[1][DATA][21] , 
        \latches_out_f[1][DATA][20] , \latches_out_f[1][DATA][19] , 
        \latches_out_f[1][DATA][18] , \latches_out_f[1][DATA][17] , 
        \latches_out_f[1][DATA][16] , \latches_out_f[1][DATA][15] , 
        \latches_out_f[1][DATA][14] , \latches_out_f[1][DATA][13] , 
        \latches_out_f[1][DATA][12] , \latches_out_f[1][DATA][11] , 
        \latches_out_f[1][DATA][10] , \latches_out_f[1][DATA][9] , 
        \latches_out_f[1][DATA][8] , \latches_out_f[1][DATA][7] , 
        \latches_out_f[1][DATA][6] , \latches_out_f[1][DATA][5] , 
        \latches_out_f[1][DATA][4] , \latches_out_f[1][DATA][3] , 
        \latches_out_f[1][DATA][2] , \latches_out_f[1][DATA][1] , 
        \latches_out_f[1][DATA][0] , \latches_out_f[0][REQ] , 
        \latches_out_f[0][DATA][34] , \latches_out_f[0][DATA][33] , 
        \latches_out_f[0][DATA][32] , \latches_out_f[0][DATA][31] , 
        \latches_out_f[0][DATA][30] , \latches_out_f[0][DATA][29] , 
        \latches_out_f[0][DATA][28] , \latches_out_f[0][DATA][27] , 
        \latches_out_f[0][DATA][26] , \latches_out_f[0][DATA][25] , 
        \latches_out_f[0][DATA][24] , \latches_out_f[0][DATA][23] , 
        \latches_out_f[0][DATA][22] , \latches_out_f[0][DATA][21] , 
        \latches_out_f[0][DATA][20] , \latches_out_f[0][DATA][19] , 
        \latches_out_f[0][DATA][18] , \latches_out_f[0][DATA][17] , 
        \latches_out_f[0][DATA][16] , \latches_out_f[0][DATA][15] , 
        \latches_out_f[0][DATA][14] , \latches_out_f[0][DATA][13] , 
        \latches_out_f[0][DATA][12] , \latches_out_f[0][DATA][11] , 
        \latches_out_f[0][DATA][10] , \latches_out_f[0][DATA][9] , 
        \latches_out_f[0][DATA][8] , \latches_out_f[0][DATA][7] , 
        \latches_out_f[0][DATA][6] , \latches_out_f[0][DATA][5] , 
        \latches_out_f[0][DATA][4] , \latches_out_f[0][DATA][3] , 
        \latches_out_f[0][DATA][2] , \latches_out_f[0][DATA][1] , 
        \latches_out_f[0][DATA][0] }), .latches_out_b({\latches_out_b[4][ACK] , 
        \latches_out_b[3][ACK] , \latches_out_b[2][ACK] , 
        \latches_out_b[1][ACK] , \latches_out_b[0][ACK] }) );
  input preset, \switch_sel[4][4] , \switch_sel[4][3] , \switch_sel[4][2] ,
         \switch_sel[4][1] , \switch_sel[4][0] , \switch_sel[3][4] ,
         \switch_sel[3][3] , \switch_sel[3][2] , \switch_sel[3][1] ,
         \switch_sel[3][0] , \switch_sel[2][4] , \switch_sel[2][3] ,
         \switch_sel[2][2] , \switch_sel[2][1] , \switch_sel[2][0] ,
         \switch_sel[1][4] , \switch_sel[1][3] , \switch_sel[1][2] ,
         \switch_sel[1][1] , \switch_sel[1][0] , \switch_sel[0][4] ,
         \switch_sel[0][3] , \switch_sel[0][2] , \switch_sel[0][1] ,
         \switch_sel[0][0] , \chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] ,
         \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] ,
         \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] ,
         \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] ,
         \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] ,
         \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] ,
         \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] ,
         \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] ,
         \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] ,
         \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] ,
         \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] ,
         \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] ,
         \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] ,
         \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] ,
         \chs_in_f[4][DATA][7] , \chs_in_f[4][DATA][6] ,
         \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] ,
         \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] ,
         \chs_in_f[4][DATA][1] , \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] ,
         \chs_in_f[3][DATA][34] , \chs_in_f[3][DATA][33] ,
         \chs_in_f[3][DATA][32] , \chs_in_f[3][DATA][31] ,
         \chs_in_f[3][DATA][30] , \chs_in_f[3][DATA][29] ,
         \chs_in_f[3][DATA][28] , \chs_in_f[3][DATA][27] ,
         \chs_in_f[3][DATA][26] , \chs_in_f[3][DATA][25] ,
         \chs_in_f[3][DATA][24] , \chs_in_f[3][DATA][23] ,
         \chs_in_f[3][DATA][22] , \chs_in_f[3][DATA][21] ,
         \chs_in_f[3][DATA][20] , \chs_in_f[3][DATA][19] ,
         \chs_in_f[3][DATA][18] , \chs_in_f[3][DATA][17] ,
         \chs_in_f[3][DATA][16] , \chs_in_f[3][DATA][15] ,
         \chs_in_f[3][DATA][14] , \chs_in_f[3][DATA][13] ,
         \chs_in_f[3][DATA][12] , \chs_in_f[3][DATA][11] ,
         \chs_in_f[3][DATA][10] , \chs_in_f[3][DATA][9] ,
         \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] ,
         \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] ,
         \chs_in_f[3][DATA][4] , \chs_in_f[3][DATA][3] ,
         \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] ,
         \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] ,
         \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] ,
         \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] ,
         \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] ,
         \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] ,
         \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] ,
         \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] ,
         \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] ,
         \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] ,
         \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] ,
         \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] ,
         \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] ,
         \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] ,
         \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] ,
         \chs_in_f[2][DATA][7] , \chs_in_f[2][DATA][6] ,
         \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] ,
         \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] ,
         \chs_in_f[2][DATA][1] , \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] ,
         \chs_in_f[1][DATA][34] , \chs_in_f[1][DATA][33] ,
         \chs_in_f[1][DATA][32] , \chs_in_f[1][DATA][31] ,
         \chs_in_f[1][DATA][30] , \chs_in_f[1][DATA][29] ,
         \chs_in_f[1][DATA][28] , \chs_in_f[1][DATA][27] ,
         \chs_in_f[1][DATA][26] , \chs_in_f[1][DATA][25] ,
         \chs_in_f[1][DATA][24] , \chs_in_f[1][DATA][23] ,
         \chs_in_f[1][DATA][22] , \chs_in_f[1][DATA][21] ,
         \chs_in_f[1][DATA][20] , \chs_in_f[1][DATA][19] ,
         \chs_in_f[1][DATA][18] , \chs_in_f[1][DATA][17] ,
         \chs_in_f[1][DATA][16] , \chs_in_f[1][DATA][15] ,
         \chs_in_f[1][DATA][14] , \chs_in_f[1][DATA][13] ,
         \chs_in_f[1][DATA][12] , \chs_in_f[1][DATA][11] ,
         \chs_in_f[1][DATA][10] , \chs_in_f[1][DATA][9] ,
         \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] ,
         \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] ,
         \chs_in_f[1][DATA][4] , \chs_in_f[1][DATA][3] ,
         \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] ,
         \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] ,
         \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] ,
         \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] ,
         \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] ,
         \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] ,
         \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] ,
         \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] ,
         \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] ,
         \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] ,
         \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] ,
         \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] ,
         \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] ,
         \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] ,
         \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] ,
         \chs_in_f[0][DATA][7] , \chs_in_f[0][DATA][6] ,
         \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] ,
         \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] ,
         \chs_in_f[0][DATA][1] , \chs_in_f[0][DATA][0] ,
         \latches_out_b[4][ACK] , \latches_out_b[3][ACK] ,
         \latches_out_b[2][ACK] , \latches_out_b[1][ACK] ,
         \latches_out_b[0][ACK] ;
  output \chs_in_b[4][ACK] , \chs_in_b[3][ACK] , \chs_in_b[2][ACK] ,
         \chs_in_b[1][ACK] , \chs_in_b[0][ACK] , \latches_out_f[4][REQ] ,
         \latches_out_f[4][DATA][34] , \latches_out_f[4][DATA][33] ,
         \latches_out_f[4][DATA][32] , \latches_out_f[4][DATA][31] ,
         \latches_out_f[4][DATA][30] , \latches_out_f[4][DATA][29] ,
         \latches_out_f[4][DATA][28] , \latches_out_f[4][DATA][27] ,
         \latches_out_f[4][DATA][26] , \latches_out_f[4][DATA][25] ,
         \latches_out_f[4][DATA][24] , \latches_out_f[4][DATA][23] ,
         \latches_out_f[4][DATA][22] , \latches_out_f[4][DATA][21] ,
         \latches_out_f[4][DATA][20] , \latches_out_f[4][DATA][19] ,
         \latches_out_f[4][DATA][18] , \latches_out_f[4][DATA][17] ,
         \latches_out_f[4][DATA][16] , \latches_out_f[4][DATA][15] ,
         \latches_out_f[4][DATA][14] , \latches_out_f[4][DATA][13] ,
         \latches_out_f[4][DATA][12] , \latches_out_f[4][DATA][11] ,
         \latches_out_f[4][DATA][10] , \latches_out_f[4][DATA][9] ,
         \latches_out_f[4][DATA][8] , \latches_out_f[4][DATA][7] ,
         \latches_out_f[4][DATA][6] , \latches_out_f[4][DATA][5] ,
         \latches_out_f[4][DATA][4] , \latches_out_f[4][DATA][3] ,
         \latches_out_f[4][DATA][2] , \latches_out_f[4][DATA][1] ,
         \latches_out_f[4][DATA][0] , \latches_out_f[3][REQ] ,
         \latches_out_f[3][DATA][34] , \latches_out_f[3][DATA][33] ,
         \latches_out_f[3][DATA][32] , \latches_out_f[3][DATA][31] ,
         \latches_out_f[3][DATA][30] , \latches_out_f[3][DATA][29] ,
         \latches_out_f[3][DATA][28] , \latches_out_f[3][DATA][27] ,
         \latches_out_f[3][DATA][26] , \latches_out_f[3][DATA][25] ,
         \latches_out_f[3][DATA][24] , \latches_out_f[3][DATA][23] ,
         \latches_out_f[3][DATA][22] , \latches_out_f[3][DATA][21] ,
         \latches_out_f[3][DATA][20] , \latches_out_f[3][DATA][19] ,
         \latches_out_f[3][DATA][18] , \latches_out_f[3][DATA][17] ,
         \latches_out_f[3][DATA][16] , \latches_out_f[3][DATA][15] ,
         \latches_out_f[3][DATA][14] , \latches_out_f[3][DATA][13] ,
         \latches_out_f[3][DATA][12] , \latches_out_f[3][DATA][11] ,
         \latches_out_f[3][DATA][10] , \latches_out_f[3][DATA][9] ,
         \latches_out_f[3][DATA][8] , \latches_out_f[3][DATA][7] ,
         \latches_out_f[3][DATA][6] , \latches_out_f[3][DATA][5] ,
         \latches_out_f[3][DATA][4] , \latches_out_f[3][DATA][3] ,
         \latches_out_f[3][DATA][2] , \latches_out_f[3][DATA][1] ,
         \latches_out_f[3][DATA][0] , \latches_out_f[2][REQ] ,
         \latches_out_f[2][DATA][34] , \latches_out_f[2][DATA][33] ,
         \latches_out_f[2][DATA][32] , \latches_out_f[2][DATA][31] ,
         \latches_out_f[2][DATA][30] , \latches_out_f[2][DATA][29] ,
         \latches_out_f[2][DATA][28] , \latches_out_f[2][DATA][27] ,
         \latches_out_f[2][DATA][26] , \latches_out_f[2][DATA][25] ,
         \latches_out_f[2][DATA][24] , \latches_out_f[2][DATA][23] ,
         \latches_out_f[2][DATA][22] , \latches_out_f[2][DATA][21] ,
         \latches_out_f[2][DATA][20] , \latches_out_f[2][DATA][19] ,
         \latches_out_f[2][DATA][18] , \latches_out_f[2][DATA][17] ,
         \latches_out_f[2][DATA][16] , \latches_out_f[2][DATA][15] ,
         \latches_out_f[2][DATA][14] , \latches_out_f[2][DATA][13] ,
         \latches_out_f[2][DATA][12] , \latches_out_f[2][DATA][11] ,
         \latches_out_f[2][DATA][10] , \latches_out_f[2][DATA][9] ,
         \latches_out_f[2][DATA][8] , \latches_out_f[2][DATA][7] ,
         \latches_out_f[2][DATA][6] , \latches_out_f[2][DATA][5] ,
         \latches_out_f[2][DATA][4] , \latches_out_f[2][DATA][3] ,
         \latches_out_f[2][DATA][2] , \latches_out_f[2][DATA][1] ,
         \latches_out_f[2][DATA][0] , \latches_out_f[1][REQ] ,
         \latches_out_f[1][DATA][34] , \latches_out_f[1][DATA][33] ,
         \latches_out_f[1][DATA][32] , \latches_out_f[1][DATA][31] ,
         \latches_out_f[1][DATA][30] , \latches_out_f[1][DATA][29] ,
         \latches_out_f[1][DATA][28] , \latches_out_f[1][DATA][27] ,
         \latches_out_f[1][DATA][26] , \latches_out_f[1][DATA][25] ,
         \latches_out_f[1][DATA][24] , \latches_out_f[1][DATA][23] ,
         \latches_out_f[1][DATA][22] , \latches_out_f[1][DATA][21] ,
         \latches_out_f[1][DATA][20] , \latches_out_f[1][DATA][19] ,
         \latches_out_f[1][DATA][18] , \latches_out_f[1][DATA][17] ,
         \latches_out_f[1][DATA][16] , \latches_out_f[1][DATA][15] ,
         \latches_out_f[1][DATA][14] , \latches_out_f[1][DATA][13] ,
         \latches_out_f[1][DATA][12] , \latches_out_f[1][DATA][11] ,
         \latches_out_f[1][DATA][10] , \latches_out_f[1][DATA][9] ,
         \latches_out_f[1][DATA][8] , \latches_out_f[1][DATA][7] ,
         \latches_out_f[1][DATA][6] , \latches_out_f[1][DATA][5] ,
         \latches_out_f[1][DATA][4] , \latches_out_f[1][DATA][3] ,
         \latches_out_f[1][DATA][2] , \latches_out_f[1][DATA][1] ,
         \latches_out_f[1][DATA][0] , \latches_out_f[0][REQ] ,
         \latches_out_f[0][DATA][34] , \latches_out_f[0][DATA][33] ,
         \latches_out_f[0][DATA][32] , \latches_out_f[0][DATA][31] ,
         \latches_out_f[0][DATA][30] , \latches_out_f[0][DATA][29] ,
         \latches_out_f[0][DATA][28] , \latches_out_f[0][DATA][27] ,
         \latches_out_f[0][DATA][26] , \latches_out_f[0][DATA][25] ,
         \latches_out_f[0][DATA][24] , \latches_out_f[0][DATA][23] ,
         \latches_out_f[0][DATA][22] , \latches_out_f[0][DATA][21] ,
         \latches_out_f[0][DATA][20] , \latches_out_f[0][DATA][19] ,
         \latches_out_f[0][DATA][18] , \latches_out_f[0][DATA][17] ,
         \latches_out_f[0][DATA][16] , \latches_out_f[0][DATA][15] ,
         \latches_out_f[0][DATA][14] , \latches_out_f[0][DATA][13] ,
         \latches_out_f[0][DATA][12] , \latches_out_f[0][DATA][11] ,
         \latches_out_f[0][DATA][10] , \latches_out_f[0][DATA][9] ,
         \latches_out_f[0][DATA][8] , \latches_out_f[0][DATA][7] ,
         \latches_out_f[0][DATA][6] , \latches_out_f[0][DATA][5] ,
         \latches_out_f[0][DATA][4] , \latches_out_f[0][DATA][3] ,
         \latches_out_f[0][DATA][2] , \latches_out_f[0][DATA][1] ,
         \latches_out_f[0][DATA][0] ;
  wire   \latches_in_f[4][REQ] , \latches_in_f[4][DATA][34] ,
         \latches_in_f[4][DATA][33] , \latches_in_f[4][DATA][32] ,
         \latches_in_f[4][DATA][31] , \latches_in_f[4][DATA][30] ,
         \latches_in_f[4][DATA][29] , \latches_in_f[4][DATA][28] ,
         \latches_in_f[4][DATA][27] , \latches_in_f[4][DATA][26] ,
         \latches_in_f[4][DATA][25] , \latches_in_f[4][DATA][24] ,
         \latches_in_f[4][DATA][23] , \latches_in_f[4][DATA][22] ,
         \latches_in_f[4][DATA][21] , \latches_in_f[4][DATA][20] ,
         \latches_in_f[4][DATA][19] , \latches_in_f[4][DATA][18] ,
         \latches_in_f[4][DATA][17] , \latches_in_f[4][DATA][16] ,
         \latches_in_f[4][DATA][15] , \latches_in_f[4][DATA][14] ,
         \latches_in_f[4][DATA][13] , \latches_in_f[4][DATA][12] ,
         \latches_in_f[4][DATA][11] , \latches_in_f[4][DATA][10] ,
         \latches_in_f[4][DATA][9] , \latches_in_f[4][DATA][8] ,
         \latches_in_f[4][DATA][7] , \latches_in_f[4][DATA][6] ,
         \latches_in_f[4][DATA][5] , \latches_in_f[4][DATA][4] ,
         \latches_in_f[4][DATA][3] , \latches_in_f[4][DATA][2] ,
         \latches_in_f[4][DATA][1] , \latches_in_f[4][DATA][0] ,
         \latches_in_f[3][REQ] , \latches_in_f[3][DATA][34] ,
         \latches_in_f[3][DATA][33] , \latches_in_f[3][DATA][32] ,
         \latches_in_f[3][DATA][31] , \latches_in_f[3][DATA][30] ,
         \latches_in_f[3][DATA][29] , \latches_in_f[3][DATA][28] ,
         \latches_in_f[3][DATA][27] , \latches_in_f[3][DATA][26] ,
         \latches_in_f[3][DATA][25] , \latches_in_f[3][DATA][24] ,
         \latches_in_f[3][DATA][23] , \latches_in_f[3][DATA][22] ,
         \latches_in_f[3][DATA][21] , \latches_in_f[3][DATA][20] ,
         \latches_in_f[3][DATA][19] , \latches_in_f[3][DATA][18] ,
         \latches_in_f[3][DATA][17] , \latches_in_f[3][DATA][16] ,
         \latches_in_f[3][DATA][15] , \latches_in_f[3][DATA][14] ,
         \latches_in_f[3][DATA][13] , \latches_in_f[3][DATA][12] ,
         \latches_in_f[3][DATA][11] , \latches_in_f[3][DATA][10] ,
         \latches_in_f[3][DATA][9] , \latches_in_f[3][DATA][8] ,
         \latches_in_f[3][DATA][7] , \latches_in_f[3][DATA][6] ,
         \latches_in_f[3][DATA][5] , \latches_in_f[3][DATA][4] ,
         \latches_in_f[3][DATA][3] , \latches_in_f[3][DATA][2] ,
         \latches_in_f[3][DATA][1] , \latches_in_f[3][DATA][0] ,
         \latches_in_f[2][REQ] , \latches_in_f[2][DATA][34] ,
         \latches_in_f[2][DATA][33] , \latches_in_f[2][DATA][32] ,
         \latches_in_f[2][DATA][31] , \latches_in_f[2][DATA][30] ,
         \latches_in_f[2][DATA][29] , \latches_in_f[2][DATA][28] ,
         \latches_in_f[2][DATA][27] , \latches_in_f[2][DATA][26] ,
         \latches_in_f[2][DATA][25] , \latches_in_f[2][DATA][24] ,
         \latches_in_f[2][DATA][23] , \latches_in_f[2][DATA][22] ,
         \latches_in_f[2][DATA][21] , \latches_in_f[2][DATA][20] ,
         \latches_in_f[2][DATA][19] , \latches_in_f[2][DATA][18] ,
         \latches_in_f[2][DATA][17] , \latches_in_f[2][DATA][16] ,
         \latches_in_f[2][DATA][15] , \latches_in_f[2][DATA][14] ,
         \latches_in_f[2][DATA][13] , \latches_in_f[2][DATA][12] ,
         \latches_in_f[2][DATA][11] , \latches_in_f[2][DATA][10] ,
         \latches_in_f[2][DATA][9] , \latches_in_f[2][DATA][8] ,
         \latches_in_f[2][DATA][7] , \latches_in_f[2][DATA][6] ,
         \latches_in_f[2][DATA][5] , \latches_in_f[2][DATA][4] ,
         \latches_in_f[2][DATA][3] , \latches_in_f[2][DATA][2] ,
         \latches_in_f[2][DATA][1] , \latches_in_f[2][DATA][0] ,
         \latches_in_f[1][REQ] , \latches_in_f[1][DATA][34] ,
         \latches_in_f[1][DATA][33] , \latches_in_f[1][DATA][32] ,
         \latches_in_f[1][DATA][31] , \latches_in_f[1][DATA][30] ,
         \latches_in_f[1][DATA][29] , \latches_in_f[1][DATA][28] ,
         \latches_in_f[1][DATA][27] , \latches_in_f[1][DATA][26] ,
         \latches_in_f[1][DATA][25] , \latches_in_f[1][DATA][24] ,
         \latches_in_f[1][DATA][23] , \latches_in_f[1][DATA][22] ,
         \latches_in_f[1][DATA][21] , \latches_in_f[1][DATA][20] ,
         \latches_in_f[1][DATA][19] , \latches_in_f[1][DATA][18] ,
         \latches_in_f[1][DATA][17] , \latches_in_f[1][DATA][16] ,
         \latches_in_f[1][DATA][15] , \latches_in_f[1][DATA][14] ,
         \latches_in_f[1][DATA][13] , \latches_in_f[1][DATA][12] ,
         \latches_in_f[1][DATA][11] , \latches_in_f[1][DATA][10] ,
         \latches_in_f[1][DATA][9] , \latches_in_f[1][DATA][8] ,
         \latches_in_f[1][DATA][7] , \latches_in_f[1][DATA][6] ,
         \latches_in_f[1][DATA][5] , \latches_in_f[1][DATA][4] ,
         \latches_in_f[1][DATA][3] , \latches_in_f[1][DATA][2] ,
         \latches_in_f[1][DATA][1] , \latches_in_f[1][DATA][0] ,
         \latches_in_f[0][REQ] , \latches_in_f[0][DATA][34] ,
         \latches_in_f[0][DATA][33] , \latches_in_f[0][DATA][32] ,
         \latches_in_f[0][DATA][31] , \latches_in_f[0][DATA][30] ,
         \latches_in_f[0][DATA][29] , \latches_in_f[0][DATA][28] ,
         \latches_in_f[0][DATA][27] , \latches_in_f[0][DATA][26] ,
         \latches_in_f[0][DATA][25] , \latches_in_f[0][DATA][24] ,
         \latches_in_f[0][DATA][23] , \latches_in_f[0][DATA][22] ,
         \latches_in_f[0][DATA][21] , \latches_in_f[0][DATA][20] ,
         \latches_in_f[0][DATA][19] , \latches_in_f[0][DATA][18] ,
         \latches_in_f[0][DATA][17] , \latches_in_f[0][DATA][16] ,
         \latches_in_f[0][DATA][15] , \latches_in_f[0][DATA][14] ,
         \latches_in_f[0][DATA][13] , \latches_in_f[0][DATA][12] ,
         \latches_in_f[0][DATA][11] , \latches_in_f[0][DATA][10] ,
         \latches_in_f[0][DATA][9] , \latches_in_f[0][DATA][8] ,
         \latches_in_f[0][DATA][7] , \latches_in_f[0][DATA][6] ,
         \latches_in_f[0][DATA][5] , \latches_in_f[0][DATA][4] ,
         \latches_in_f[0][DATA][3] , \latches_in_f[0][DATA][2] ,
         \latches_in_f[0][DATA][1] , \latches_in_f[0][DATA][0] ,
         \latches_in_b[4][ACK] , \latches_in_b[3][ACK] ,
         \latches_in_b[2][ACK] , \latches_in_b[1][ACK] ,
         \latches_in_b[0][ACK] , n1;

  crossbar_0 crossbar ( .preset(n1), .switch_sel({\switch_sel[4][4] , 
        \switch_sel[4][3] , \switch_sel[4][2] , \switch_sel[4][1] , 
        \switch_sel[4][0] , \switch_sel[3][4] , \switch_sel[3][3] , 
        \switch_sel[3][2] , \switch_sel[3][1] , \switch_sel[3][0] , 
        \switch_sel[2][4] , \switch_sel[2][3] , \switch_sel[2][2] , 
        \switch_sel[2][1] , \switch_sel[2][0] , \switch_sel[1][4] , 
        \switch_sel[1][3] , \switch_sel[1][2] , \switch_sel[1][1] , 
        \switch_sel[1][0] , \switch_sel[0][4] , \switch_sel[0][3] , 
        \switch_sel[0][2] , \switch_sel[0][1] , \switch_sel[0][0] }), 
        .chs_in_f({\chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] , 
        \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] , 
        \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] , 
        \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] , 
        \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] , 
        \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] , 
        \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] , 
        \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] , 
        \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] , 
        \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] , 
        \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] , 
        \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] , 
        \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] , 
        \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] , \chs_in_f[4][DATA][7] , 
        \chs_in_f[4][DATA][6] , \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] , 
        \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] , \chs_in_f[4][DATA][1] , 
        \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] , \chs_in_f[3][DATA][34] , 
        \chs_in_f[3][DATA][33] , \chs_in_f[3][DATA][32] , 
        \chs_in_f[3][DATA][31] , \chs_in_f[3][DATA][30] , 
        \chs_in_f[3][DATA][29] , \chs_in_f[3][DATA][28] , 
        \chs_in_f[3][DATA][27] , \chs_in_f[3][DATA][26] , 
        \chs_in_f[3][DATA][25] , \chs_in_f[3][DATA][24] , 
        \chs_in_f[3][DATA][23] , \chs_in_f[3][DATA][22] , 
        \chs_in_f[3][DATA][21] , \chs_in_f[3][DATA][20] , 
        \chs_in_f[3][DATA][19] , \chs_in_f[3][DATA][18] , 
        \chs_in_f[3][DATA][17] , \chs_in_f[3][DATA][16] , 
        \chs_in_f[3][DATA][15] , \chs_in_f[3][DATA][14] , 
        \chs_in_f[3][DATA][13] , \chs_in_f[3][DATA][12] , 
        \chs_in_f[3][DATA][11] , \chs_in_f[3][DATA][10] , 
        \chs_in_f[3][DATA][9] , \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] , 
        \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] , \chs_in_f[3][DATA][4] , 
        \chs_in_f[3][DATA][3] , \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] , 
        \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] , 
        \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] , 
        \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] , 
        \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] , 
        \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] , 
        \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] , 
        \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] , 
        \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] , 
        \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] , 
        \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] , 
        \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] , 
        \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] , 
        \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] , 
        \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] , \chs_in_f[2][DATA][7] , 
        \chs_in_f[2][DATA][6] , \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] , 
        \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] , \chs_in_f[2][DATA][1] , 
        \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] , \chs_in_f[1][DATA][34] , 
        \chs_in_f[1][DATA][33] , \chs_in_f[1][DATA][32] , 
        \chs_in_f[1][DATA][31] , \chs_in_f[1][DATA][30] , 
        \chs_in_f[1][DATA][29] , \chs_in_f[1][DATA][28] , 
        \chs_in_f[1][DATA][27] , \chs_in_f[1][DATA][26] , 
        \chs_in_f[1][DATA][25] , \chs_in_f[1][DATA][24] , 
        \chs_in_f[1][DATA][23] , \chs_in_f[1][DATA][22] , 
        \chs_in_f[1][DATA][21] , \chs_in_f[1][DATA][20] , 
        \chs_in_f[1][DATA][19] , \chs_in_f[1][DATA][18] , 
        \chs_in_f[1][DATA][17] , \chs_in_f[1][DATA][16] , 
        \chs_in_f[1][DATA][15] , \chs_in_f[1][DATA][14] , 
        \chs_in_f[1][DATA][13] , \chs_in_f[1][DATA][12] , 
        \chs_in_f[1][DATA][11] , \chs_in_f[1][DATA][10] , 
        \chs_in_f[1][DATA][9] , \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] , 
        \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] , \chs_in_f[1][DATA][4] , 
        \chs_in_f[1][DATA][3] , \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] , 
        \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] , 
        \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] , 
        \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] , 
        \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] , 
        \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] , 
        \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] , 
        \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] , 
        \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] , 
        \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] , 
        \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] , 
        \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] , 
        \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] , 
        \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] , 
        \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] , \chs_in_f[0][DATA][7] , 
        \chs_in_f[0][DATA][6] , \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] , 
        \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] , \chs_in_f[0][DATA][1] , 
        \chs_in_f[0][DATA][0] }), .chs_in_b({\chs_in_b[4][ACK] , 
        \chs_in_b[3][ACK] , \chs_in_b[2][ACK] , \chs_in_b[1][ACK] , 
        \chs_in_b[0][ACK] }), .chs_out_f({\latches_in_f[4][REQ] , 
        \latches_in_f[4][DATA][34] , \latches_in_f[4][DATA][33] , 
        \latches_in_f[4][DATA][32] , \latches_in_f[4][DATA][31] , 
        \latches_in_f[4][DATA][30] , \latches_in_f[4][DATA][29] , 
        \latches_in_f[4][DATA][28] , \latches_in_f[4][DATA][27] , 
        \latches_in_f[4][DATA][26] , \latches_in_f[4][DATA][25] , 
        \latches_in_f[4][DATA][24] , \latches_in_f[4][DATA][23] , 
        \latches_in_f[4][DATA][22] , \latches_in_f[4][DATA][21] , 
        \latches_in_f[4][DATA][20] , \latches_in_f[4][DATA][19] , 
        \latches_in_f[4][DATA][18] , \latches_in_f[4][DATA][17] , 
        \latches_in_f[4][DATA][16] , \latches_in_f[4][DATA][15] , 
        \latches_in_f[4][DATA][14] , \latches_in_f[4][DATA][13] , 
        \latches_in_f[4][DATA][12] , \latches_in_f[4][DATA][11] , 
        \latches_in_f[4][DATA][10] , \latches_in_f[4][DATA][9] , 
        \latches_in_f[4][DATA][8] , \latches_in_f[4][DATA][7] , 
        \latches_in_f[4][DATA][6] , \latches_in_f[4][DATA][5] , 
        \latches_in_f[4][DATA][4] , \latches_in_f[4][DATA][3] , 
        \latches_in_f[4][DATA][2] , \latches_in_f[4][DATA][1] , 
        \latches_in_f[4][DATA][0] , \latches_in_f[3][REQ] , 
        \latches_in_f[3][DATA][34] , \latches_in_f[3][DATA][33] , 
        \latches_in_f[3][DATA][32] , \latches_in_f[3][DATA][31] , 
        \latches_in_f[3][DATA][30] , \latches_in_f[3][DATA][29] , 
        \latches_in_f[3][DATA][28] , \latches_in_f[3][DATA][27] , 
        \latches_in_f[3][DATA][26] , \latches_in_f[3][DATA][25] , 
        \latches_in_f[3][DATA][24] , \latches_in_f[3][DATA][23] , 
        \latches_in_f[3][DATA][22] , \latches_in_f[3][DATA][21] , 
        \latches_in_f[3][DATA][20] , \latches_in_f[3][DATA][19] , 
        \latches_in_f[3][DATA][18] , \latches_in_f[3][DATA][17] , 
        \latches_in_f[3][DATA][16] , \latches_in_f[3][DATA][15] , 
        \latches_in_f[3][DATA][14] , \latches_in_f[3][DATA][13] , 
        \latches_in_f[3][DATA][12] , \latches_in_f[3][DATA][11] , 
        \latches_in_f[3][DATA][10] , \latches_in_f[3][DATA][9] , 
        \latches_in_f[3][DATA][8] , \latches_in_f[3][DATA][7] , 
        \latches_in_f[3][DATA][6] , \latches_in_f[3][DATA][5] , 
        \latches_in_f[3][DATA][4] , \latches_in_f[3][DATA][3] , 
        \latches_in_f[3][DATA][2] , \latches_in_f[3][DATA][1] , 
        \latches_in_f[3][DATA][0] , \latches_in_f[2][REQ] , 
        \latches_in_f[2][DATA][34] , \latches_in_f[2][DATA][33] , 
        \latches_in_f[2][DATA][32] , \latches_in_f[2][DATA][31] , 
        \latches_in_f[2][DATA][30] , \latches_in_f[2][DATA][29] , 
        \latches_in_f[2][DATA][28] , \latches_in_f[2][DATA][27] , 
        \latches_in_f[2][DATA][26] , \latches_in_f[2][DATA][25] , 
        \latches_in_f[2][DATA][24] , \latches_in_f[2][DATA][23] , 
        \latches_in_f[2][DATA][22] , \latches_in_f[2][DATA][21] , 
        \latches_in_f[2][DATA][20] , \latches_in_f[2][DATA][19] , 
        \latches_in_f[2][DATA][18] , \latches_in_f[2][DATA][17] , 
        \latches_in_f[2][DATA][16] , \latches_in_f[2][DATA][15] , 
        \latches_in_f[2][DATA][14] , \latches_in_f[2][DATA][13] , 
        \latches_in_f[2][DATA][12] , \latches_in_f[2][DATA][11] , 
        \latches_in_f[2][DATA][10] , \latches_in_f[2][DATA][9] , 
        \latches_in_f[2][DATA][8] , \latches_in_f[2][DATA][7] , 
        \latches_in_f[2][DATA][6] , \latches_in_f[2][DATA][5] , 
        \latches_in_f[2][DATA][4] , \latches_in_f[2][DATA][3] , 
        \latches_in_f[2][DATA][2] , \latches_in_f[2][DATA][1] , 
        \latches_in_f[2][DATA][0] , \latches_in_f[1][REQ] , 
        \latches_in_f[1][DATA][34] , \latches_in_f[1][DATA][33] , 
        \latches_in_f[1][DATA][32] , \latches_in_f[1][DATA][31] , 
        \latches_in_f[1][DATA][30] , \latches_in_f[1][DATA][29] , 
        \latches_in_f[1][DATA][28] , \latches_in_f[1][DATA][27] , 
        \latches_in_f[1][DATA][26] , \latches_in_f[1][DATA][25] , 
        \latches_in_f[1][DATA][24] , \latches_in_f[1][DATA][23] , 
        \latches_in_f[1][DATA][22] , \latches_in_f[1][DATA][21] , 
        \latches_in_f[1][DATA][20] , \latches_in_f[1][DATA][19] , 
        \latches_in_f[1][DATA][18] , \latches_in_f[1][DATA][17] , 
        \latches_in_f[1][DATA][16] , \latches_in_f[1][DATA][15] , 
        \latches_in_f[1][DATA][14] , \latches_in_f[1][DATA][13] , 
        \latches_in_f[1][DATA][12] , \latches_in_f[1][DATA][11] , 
        \latches_in_f[1][DATA][10] , \latches_in_f[1][DATA][9] , 
        \latches_in_f[1][DATA][8] , \latches_in_f[1][DATA][7] , 
        \latches_in_f[1][DATA][6] , \latches_in_f[1][DATA][5] , 
        \latches_in_f[1][DATA][4] , \latches_in_f[1][DATA][3] , 
        \latches_in_f[1][DATA][2] , \latches_in_f[1][DATA][1] , 
        \latches_in_f[1][DATA][0] , \latches_in_f[0][REQ] , 
        \latches_in_f[0][DATA][34] , \latches_in_f[0][DATA][33] , 
        \latches_in_f[0][DATA][32] , \latches_in_f[0][DATA][31] , 
        \latches_in_f[0][DATA][30] , \latches_in_f[0][DATA][29] , 
        \latches_in_f[0][DATA][28] , \latches_in_f[0][DATA][27] , 
        \latches_in_f[0][DATA][26] , \latches_in_f[0][DATA][25] , 
        \latches_in_f[0][DATA][24] , \latches_in_f[0][DATA][23] , 
        \latches_in_f[0][DATA][22] , \latches_in_f[0][DATA][21] , 
        \latches_in_f[0][DATA][20] , \latches_in_f[0][DATA][19] , 
        \latches_in_f[0][DATA][18] , \latches_in_f[0][DATA][17] , 
        \latches_in_f[0][DATA][16] , \latches_in_f[0][DATA][15] , 
        \latches_in_f[0][DATA][14] , \latches_in_f[0][DATA][13] , 
        \latches_in_f[0][DATA][12] , \latches_in_f[0][DATA][11] , 
        \latches_in_f[0][DATA][10] , \latches_in_f[0][DATA][9] , 
        \latches_in_f[0][DATA][8] , \latches_in_f[0][DATA][7] , 
        \latches_in_f[0][DATA][6] , \latches_in_f[0][DATA][5] , 
        \latches_in_f[0][DATA][4] , \latches_in_f[0][DATA][3] , 
        \latches_in_f[0][DATA][2] , \latches_in_f[0][DATA][1] , 
        \latches_in_f[0][DATA][0] }), .chs_out_b({\latches_in_b[4][ACK] , 
        \latches_in_b[3][ACK] , \latches_in_b[2][ACK] , \latches_in_b[1][ACK] , 
        \latches_in_b[0][ACK] }) );
  channel_latch_0_000000000_0 ch_latch_4 ( .preset(n1), .left_in({
        \latches_in_f[4][REQ] , \latches_in_f[4][DATA][34] , 
        \latches_in_f[4][DATA][33] , \latches_in_f[4][DATA][32] , 
        \latches_in_f[4][DATA][31] , \latches_in_f[4][DATA][30] , 
        \latches_in_f[4][DATA][29] , \latches_in_f[4][DATA][28] , 
        \latches_in_f[4][DATA][27] , \latches_in_f[4][DATA][26] , 
        \latches_in_f[4][DATA][25] , \latches_in_f[4][DATA][24] , 
        \latches_in_f[4][DATA][23] , \latches_in_f[4][DATA][22] , 
        \latches_in_f[4][DATA][21] , \latches_in_f[4][DATA][20] , 
        \latches_in_f[4][DATA][19] , \latches_in_f[4][DATA][18] , 
        \latches_in_f[4][DATA][17] , \latches_in_f[4][DATA][16] , 
        \latches_in_f[4][DATA][15] , \latches_in_f[4][DATA][14] , 
        \latches_in_f[4][DATA][13] , \latches_in_f[4][DATA][12] , 
        \latches_in_f[4][DATA][11] , \latches_in_f[4][DATA][10] , 
        \latches_in_f[4][DATA][9] , \latches_in_f[4][DATA][8] , 
        \latches_in_f[4][DATA][7] , \latches_in_f[4][DATA][6] , 
        \latches_in_f[4][DATA][5] , \latches_in_f[4][DATA][4] , 
        \latches_in_f[4][DATA][3] , \latches_in_f[4][DATA][2] , 
        \latches_in_f[4][DATA][1] , \latches_in_f[4][DATA][0] }), .left_out(
        \latches_in_b[4][ACK] ), .right_out({\latches_out_f[4][REQ] , 
        \latches_out_f[4][DATA][34] , \latches_out_f[4][DATA][33] , 
        \latches_out_f[4][DATA][32] , \latches_out_f[4][DATA][31] , 
        \latches_out_f[4][DATA][30] , \latches_out_f[4][DATA][29] , 
        \latches_out_f[4][DATA][28] , \latches_out_f[4][DATA][27] , 
        \latches_out_f[4][DATA][26] , \latches_out_f[4][DATA][25] , 
        \latches_out_f[4][DATA][24] , \latches_out_f[4][DATA][23] , 
        \latches_out_f[4][DATA][22] , \latches_out_f[4][DATA][21] , 
        \latches_out_f[4][DATA][20] , \latches_out_f[4][DATA][19] , 
        \latches_out_f[4][DATA][18] , \latches_out_f[4][DATA][17] , 
        \latches_out_f[4][DATA][16] , \latches_out_f[4][DATA][15] , 
        \latches_out_f[4][DATA][14] , \latches_out_f[4][DATA][13] , 
        \latches_out_f[4][DATA][12] , \latches_out_f[4][DATA][11] , 
        \latches_out_f[4][DATA][10] , \latches_out_f[4][DATA][9] , 
        \latches_out_f[4][DATA][8] , \latches_out_f[4][DATA][7] , 
        \latches_out_f[4][DATA][6] , \latches_out_f[4][DATA][5] , 
        \latches_out_f[4][DATA][4] , \latches_out_f[4][DATA][3] , 
        \latches_out_f[4][DATA][2] , \latches_out_f[4][DATA][1] , 
        \latches_out_f[4][DATA][0] }), .right_in(\latches_out_b[4][ACK] ) );
  channel_latch_0_000000000_19 ch_latch_3 ( .preset(n1), .left_in({
        \latches_in_f[3][REQ] , \latches_in_f[3][DATA][34] , 
        \latches_in_f[3][DATA][33] , \latches_in_f[3][DATA][32] , 
        \latches_in_f[3][DATA][31] , \latches_in_f[3][DATA][30] , 
        \latches_in_f[3][DATA][29] , \latches_in_f[3][DATA][28] , 
        \latches_in_f[3][DATA][27] , \latches_in_f[3][DATA][26] , 
        \latches_in_f[3][DATA][25] , \latches_in_f[3][DATA][24] , 
        \latches_in_f[3][DATA][23] , \latches_in_f[3][DATA][22] , 
        \latches_in_f[3][DATA][21] , \latches_in_f[3][DATA][20] , 
        \latches_in_f[3][DATA][19] , \latches_in_f[3][DATA][18] , 
        \latches_in_f[3][DATA][17] , \latches_in_f[3][DATA][16] , 
        \latches_in_f[3][DATA][15] , \latches_in_f[3][DATA][14] , 
        \latches_in_f[3][DATA][13] , \latches_in_f[3][DATA][12] , 
        \latches_in_f[3][DATA][11] , \latches_in_f[3][DATA][10] , 
        \latches_in_f[3][DATA][9] , \latches_in_f[3][DATA][8] , 
        \latches_in_f[3][DATA][7] , \latches_in_f[3][DATA][6] , 
        \latches_in_f[3][DATA][5] , \latches_in_f[3][DATA][4] , 
        \latches_in_f[3][DATA][3] , \latches_in_f[3][DATA][2] , 
        \latches_in_f[3][DATA][1] , \latches_in_f[3][DATA][0] }), .left_out(
        \latches_in_b[3][ACK] ), .right_out({\latches_out_f[3][REQ] , 
        \latches_out_f[3][DATA][34] , \latches_out_f[3][DATA][33] , 
        \latches_out_f[3][DATA][32] , \latches_out_f[3][DATA][31] , 
        \latches_out_f[3][DATA][30] , \latches_out_f[3][DATA][29] , 
        \latches_out_f[3][DATA][28] , \latches_out_f[3][DATA][27] , 
        \latches_out_f[3][DATA][26] , \latches_out_f[3][DATA][25] , 
        \latches_out_f[3][DATA][24] , \latches_out_f[3][DATA][23] , 
        \latches_out_f[3][DATA][22] , \latches_out_f[3][DATA][21] , 
        \latches_out_f[3][DATA][20] , \latches_out_f[3][DATA][19] , 
        \latches_out_f[3][DATA][18] , \latches_out_f[3][DATA][17] , 
        \latches_out_f[3][DATA][16] , \latches_out_f[3][DATA][15] , 
        \latches_out_f[3][DATA][14] , \latches_out_f[3][DATA][13] , 
        \latches_out_f[3][DATA][12] , \latches_out_f[3][DATA][11] , 
        \latches_out_f[3][DATA][10] , \latches_out_f[3][DATA][9] , 
        \latches_out_f[3][DATA][8] , \latches_out_f[3][DATA][7] , 
        \latches_out_f[3][DATA][6] , \latches_out_f[3][DATA][5] , 
        \latches_out_f[3][DATA][4] , \latches_out_f[3][DATA][3] , 
        \latches_out_f[3][DATA][2] , \latches_out_f[3][DATA][1] , 
        \latches_out_f[3][DATA][0] }), .right_in(\latches_out_b[3][ACK] ) );
  channel_latch_0_000000000_18 ch_latch_2 ( .preset(n1), .left_in({
        \latches_in_f[2][REQ] , \latches_in_f[2][DATA][34] , 
        \latches_in_f[2][DATA][33] , \latches_in_f[2][DATA][32] , 
        \latches_in_f[2][DATA][31] , \latches_in_f[2][DATA][30] , 
        \latches_in_f[2][DATA][29] , \latches_in_f[2][DATA][28] , 
        \latches_in_f[2][DATA][27] , \latches_in_f[2][DATA][26] , 
        \latches_in_f[2][DATA][25] , \latches_in_f[2][DATA][24] , 
        \latches_in_f[2][DATA][23] , \latches_in_f[2][DATA][22] , 
        \latches_in_f[2][DATA][21] , \latches_in_f[2][DATA][20] , 
        \latches_in_f[2][DATA][19] , \latches_in_f[2][DATA][18] , 
        \latches_in_f[2][DATA][17] , \latches_in_f[2][DATA][16] , 
        \latches_in_f[2][DATA][15] , \latches_in_f[2][DATA][14] , 
        \latches_in_f[2][DATA][13] , \latches_in_f[2][DATA][12] , 
        \latches_in_f[2][DATA][11] , \latches_in_f[2][DATA][10] , 
        \latches_in_f[2][DATA][9] , \latches_in_f[2][DATA][8] , 
        \latches_in_f[2][DATA][7] , \latches_in_f[2][DATA][6] , 
        \latches_in_f[2][DATA][5] , \latches_in_f[2][DATA][4] , 
        \latches_in_f[2][DATA][3] , \latches_in_f[2][DATA][2] , 
        \latches_in_f[2][DATA][1] , \latches_in_f[2][DATA][0] }), .left_out(
        \latches_in_b[2][ACK] ), .right_out({\latches_out_f[2][REQ] , 
        \latches_out_f[2][DATA][34] , \latches_out_f[2][DATA][33] , 
        \latches_out_f[2][DATA][32] , \latches_out_f[2][DATA][31] , 
        \latches_out_f[2][DATA][30] , \latches_out_f[2][DATA][29] , 
        \latches_out_f[2][DATA][28] , \latches_out_f[2][DATA][27] , 
        \latches_out_f[2][DATA][26] , \latches_out_f[2][DATA][25] , 
        \latches_out_f[2][DATA][24] , \latches_out_f[2][DATA][23] , 
        \latches_out_f[2][DATA][22] , \latches_out_f[2][DATA][21] , 
        \latches_out_f[2][DATA][20] , \latches_out_f[2][DATA][19] , 
        \latches_out_f[2][DATA][18] , \latches_out_f[2][DATA][17] , 
        \latches_out_f[2][DATA][16] , \latches_out_f[2][DATA][15] , 
        \latches_out_f[2][DATA][14] , \latches_out_f[2][DATA][13] , 
        \latches_out_f[2][DATA][12] , \latches_out_f[2][DATA][11] , 
        \latches_out_f[2][DATA][10] , \latches_out_f[2][DATA][9] , 
        \latches_out_f[2][DATA][8] , \latches_out_f[2][DATA][7] , 
        \latches_out_f[2][DATA][6] , \latches_out_f[2][DATA][5] , 
        \latches_out_f[2][DATA][4] , \latches_out_f[2][DATA][3] , 
        \latches_out_f[2][DATA][2] , \latches_out_f[2][DATA][1] , 
        \latches_out_f[2][DATA][0] }), .right_in(\latches_out_b[2][ACK] ) );
  channel_latch_0_000000000_17 ch_latch_1 ( .preset(n1), .left_in({
        \latches_in_f[1][REQ] , \latches_in_f[1][DATA][34] , 
        \latches_in_f[1][DATA][33] , \latches_in_f[1][DATA][32] , 
        \latches_in_f[1][DATA][31] , \latches_in_f[1][DATA][30] , 
        \latches_in_f[1][DATA][29] , \latches_in_f[1][DATA][28] , 
        \latches_in_f[1][DATA][27] , \latches_in_f[1][DATA][26] , 
        \latches_in_f[1][DATA][25] , \latches_in_f[1][DATA][24] , 
        \latches_in_f[1][DATA][23] , \latches_in_f[1][DATA][22] , 
        \latches_in_f[1][DATA][21] , \latches_in_f[1][DATA][20] , 
        \latches_in_f[1][DATA][19] , \latches_in_f[1][DATA][18] , 
        \latches_in_f[1][DATA][17] , \latches_in_f[1][DATA][16] , 
        \latches_in_f[1][DATA][15] , \latches_in_f[1][DATA][14] , 
        \latches_in_f[1][DATA][13] , \latches_in_f[1][DATA][12] , 
        \latches_in_f[1][DATA][11] , \latches_in_f[1][DATA][10] , 
        \latches_in_f[1][DATA][9] , \latches_in_f[1][DATA][8] , 
        \latches_in_f[1][DATA][7] , \latches_in_f[1][DATA][6] , 
        \latches_in_f[1][DATA][5] , \latches_in_f[1][DATA][4] , 
        \latches_in_f[1][DATA][3] , \latches_in_f[1][DATA][2] , 
        \latches_in_f[1][DATA][1] , \latches_in_f[1][DATA][0] }), .left_out(
        \latches_in_b[1][ACK] ), .right_out({\latches_out_f[1][REQ] , 
        \latches_out_f[1][DATA][34] , \latches_out_f[1][DATA][33] , 
        \latches_out_f[1][DATA][32] , \latches_out_f[1][DATA][31] , 
        \latches_out_f[1][DATA][30] , \latches_out_f[1][DATA][29] , 
        \latches_out_f[1][DATA][28] , \latches_out_f[1][DATA][27] , 
        \latches_out_f[1][DATA][26] , \latches_out_f[1][DATA][25] , 
        \latches_out_f[1][DATA][24] , \latches_out_f[1][DATA][23] , 
        \latches_out_f[1][DATA][22] , \latches_out_f[1][DATA][21] , 
        \latches_out_f[1][DATA][20] , \latches_out_f[1][DATA][19] , 
        \latches_out_f[1][DATA][18] , \latches_out_f[1][DATA][17] , 
        \latches_out_f[1][DATA][16] , \latches_out_f[1][DATA][15] , 
        \latches_out_f[1][DATA][14] , \latches_out_f[1][DATA][13] , 
        \latches_out_f[1][DATA][12] , \latches_out_f[1][DATA][11] , 
        \latches_out_f[1][DATA][10] , \latches_out_f[1][DATA][9] , 
        \latches_out_f[1][DATA][8] , \latches_out_f[1][DATA][7] , 
        \latches_out_f[1][DATA][6] , \latches_out_f[1][DATA][5] , 
        \latches_out_f[1][DATA][4] , \latches_out_f[1][DATA][3] , 
        \latches_out_f[1][DATA][2] , \latches_out_f[1][DATA][1] , 
        \latches_out_f[1][DATA][0] }), .right_in(\latches_out_b[1][ACK] ) );
  channel_latch_0_000000000_16 ch_latch_0 ( .preset(n1), .left_in({
        \latches_in_f[0][REQ] , \latches_in_f[0][DATA][34] , 
        \latches_in_f[0][DATA][33] , \latches_in_f[0][DATA][32] , 
        \latches_in_f[0][DATA][31] , \latches_in_f[0][DATA][30] , 
        \latches_in_f[0][DATA][29] , \latches_in_f[0][DATA][28] , 
        \latches_in_f[0][DATA][27] , \latches_in_f[0][DATA][26] , 
        \latches_in_f[0][DATA][25] , \latches_in_f[0][DATA][24] , 
        \latches_in_f[0][DATA][23] , \latches_in_f[0][DATA][22] , 
        \latches_in_f[0][DATA][21] , \latches_in_f[0][DATA][20] , 
        \latches_in_f[0][DATA][19] , \latches_in_f[0][DATA][18] , 
        \latches_in_f[0][DATA][17] , \latches_in_f[0][DATA][16] , 
        \latches_in_f[0][DATA][15] , \latches_in_f[0][DATA][14] , 
        \latches_in_f[0][DATA][13] , \latches_in_f[0][DATA][12] , 
        \latches_in_f[0][DATA][11] , \latches_in_f[0][DATA][10] , 
        \latches_in_f[0][DATA][9] , \latches_in_f[0][DATA][8] , 
        \latches_in_f[0][DATA][7] , \latches_in_f[0][DATA][6] , 
        \latches_in_f[0][DATA][5] , \latches_in_f[0][DATA][4] , 
        \latches_in_f[0][DATA][3] , \latches_in_f[0][DATA][2] , 
        \latches_in_f[0][DATA][1] , \latches_in_f[0][DATA][0] }), .left_out(
        \latches_in_b[0][ACK] ), .right_out({\latches_out_f[0][REQ] , 
        \latches_out_f[0][DATA][34] , \latches_out_f[0][DATA][33] , 
        \latches_out_f[0][DATA][32] , \latches_out_f[0][DATA][31] , 
        \latches_out_f[0][DATA][30] , \latches_out_f[0][DATA][29] , 
        \latches_out_f[0][DATA][28] , \latches_out_f[0][DATA][27] , 
        \latches_out_f[0][DATA][26] , \latches_out_f[0][DATA][25] , 
        \latches_out_f[0][DATA][24] , \latches_out_f[0][DATA][23] , 
        \latches_out_f[0][DATA][22] , \latches_out_f[0][DATA][21] , 
        \latches_out_f[0][DATA][20] , \latches_out_f[0][DATA][19] , 
        \latches_out_f[0][DATA][18] , \latches_out_f[0][DATA][17] , 
        \latches_out_f[0][DATA][16] , \latches_out_f[0][DATA][15] , 
        \latches_out_f[0][DATA][14] , \latches_out_f[0][DATA][13] , 
        \latches_out_f[0][DATA][12] , \latches_out_f[0][DATA][11] , 
        \latches_out_f[0][DATA][10] , \latches_out_f[0][DATA][9] , 
        \latches_out_f[0][DATA][8] , \latches_out_f[0][DATA][7] , 
        \latches_out_f[0][DATA][6] , \latches_out_f[0][DATA][5] , 
        \latches_out_f[0][DATA][4] , \latches_out_f[0][DATA][3] , 
        \latches_out_f[0][DATA][2] , \latches_out_f[0][DATA][1] , 
        \latches_out_f[0][DATA][0] }), .right_in(\latches_out_b[0][ACK] ) );
  HS65_LS_BFX9 U1 ( .A(preset), .Z(n1) );
endmodule


module noc_switch_0 ( preset, .north_in_f({\north_in_f[REQ] , 
        \north_in_f[DATA][34] , \north_in_f[DATA][33] , \north_in_f[DATA][32] , 
        \north_in_f[DATA][31] , \north_in_f[DATA][30] , \north_in_f[DATA][29] , 
        \north_in_f[DATA][28] , \north_in_f[DATA][27] , \north_in_f[DATA][26] , 
        \north_in_f[DATA][25] , \north_in_f[DATA][24] , \north_in_f[DATA][23] , 
        \north_in_f[DATA][22] , \north_in_f[DATA][21] , \north_in_f[DATA][20] , 
        \north_in_f[DATA][19] , \north_in_f[DATA][18] , \north_in_f[DATA][17] , 
        \north_in_f[DATA][16] , \north_in_f[DATA][15] , \north_in_f[DATA][14] , 
        \north_in_f[DATA][13] , \north_in_f[DATA][12] , \north_in_f[DATA][11] , 
        \north_in_f[DATA][10] , \north_in_f[DATA][9] , \north_in_f[DATA][8] , 
        \north_in_f[DATA][7] , \north_in_f[DATA][6] , \north_in_f[DATA][5] , 
        \north_in_f[DATA][4] , \north_in_f[DATA][3] , \north_in_f[DATA][2] , 
        \north_in_f[DATA][1] , \north_in_f[DATA][0] }), .north_in_b(
        \north_in_b[ACK] ), .east_in_f({\east_in_f[REQ] , 
        \east_in_f[DATA][34] , \east_in_f[DATA][33] , \east_in_f[DATA][32] , 
        \east_in_f[DATA][31] , \east_in_f[DATA][30] , \east_in_f[DATA][29] , 
        \east_in_f[DATA][28] , \east_in_f[DATA][27] , \east_in_f[DATA][26] , 
        \east_in_f[DATA][25] , \east_in_f[DATA][24] , \east_in_f[DATA][23] , 
        \east_in_f[DATA][22] , \east_in_f[DATA][21] , \east_in_f[DATA][20] , 
        \east_in_f[DATA][19] , \east_in_f[DATA][18] , \east_in_f[DATA][17] , 
        \east_in_f[DATA][16] , \east_in_f[DATA][15] , \east_in_f[DATA][14] , 
        \east_in_f[DATA][13] , \east_in_f[DATA][12] , \east_in_f[DATA][11] , 
        \east_in_f[DATA][10] , \east_in_f[DATA][9] , \east_in_f[DATA][8] , 
        \east_in_f[DATA][7] , \east_in_f[DATA][6] , \east_in_f[DATA][5] , 
        \east_in_f[DATA][4] , \east_in_f[DATA][3] , \east_in_f[DATA][2] , 
        \east_in_f[DATA][1] , \east_in_f[DATA][0] }), .east_in_b(
        \east_in_b[ACK] ), .south_in_f({\south_in_f[REQ] , 
        \south_in_f[DATA][34] , \south_in_f[DATA][33] , \south_in_f[DATA][32] , 
        \south_in_f[DATA][31] , \south_in_f[DATA][30] , \south_in_f[DATA][29] , 
        \south_in_f[DATA][28] , \south_in_f[DATA][27] , \south_in_f[DATA][26] , 
        \south_in_f[DATA][25] , \south_in_f[DATA][24] , \south_in_f[DATA][23] , 
        \south_in_f[DATA][22] , \south_in_f[DATA][21] , \south_in_f[DATA][20] , 
        \south_in_f[DATA][19] , \south_in_f[DATA][18] , \south_in_f[DATA][17] , 
        \south_in_f[DATA][16] , \south_in_f[DATA][15] , \south_in_f[DATA][14] , 
        \south_in_f[DATA][13] , \south_in_f[DATA][12] , \south_in_f[DATA][11] , 
        \south_in_f[DATA][10] , \south_in_f[DATA][9] , \south_in_f[DATA][8] , 
        \south_in_f[DATA][7] , \south_in_f[DATA][6] , \south_in_f[DATA][5] , 
        \south_in_f[DATA][4] , \south_in_f[DATA][3] , \south_in_f[DATA][2] , 
        \south_in_f[DATA][1] , \south_in_f[DATA][0] }), .south_in_b(
        \south_in_b[ACK] ), .west_in_f({\west_in_f[REQ] , 
        \west_in_f[DATA][34] , \west_in_f[DATA][33] , \west_in_f[DATA][32] , 
        \west_in_f[DATA][31] , \west_in_f[DATA][30] , \west_in_f[DATA][29] , 
        \west_in_f[DATA][28] , \west_in_f[DATA][27] , \west_in_f[DATA][26] , 
        \west_in_f[DATA][25] , \west_in_f[DATA][24] , \west_in_f[DATA][23] , 
        \west_in_f[DATA][22] , \west_in_f[DATA][21] , \west_in_f[DATA][20] , 
        \west_in_f[DATA][19] , \west_in_f[DATA][18] , \west_in_f[DATA][17] , 
        \west_in_f[DATA][16] , \west_in_f[DATA][15] , \west_in_f[DATA][14] , 
        \west_in_f[DATA][13] , \west_in_f[DATA][12] , \west_in_f[DATA][11] , 
        \west_in_f[DATA][10] , \west_in_f[DATA][9] , \west_in_f[DATA][8] , 
        \west_in_f[DATA][7] , \west_in_f[DATA][6] , \west_in_f[DATA][5] , 
        \west_in_f[DATA][4] , \west_in_f[DATA][3] , \west_in_f[DATA][2] , 
        \west_in_f[DATA][1] , \west_in_f[DATA][0] }), .west_in_b(
        \west_in_b[ACK] ), .resource_in_f({\resource_in_f[REQ] , 
        \resource_in_f[DATA][34] , \resource_in_f[DATA][33] , 
        \resource_in_f[DATA][32] , \resource_in_f[DATA][31] , 
        \resource_in_f[DATA][30] , \resource_in_f[DATA][29] , 
        \resource_in_f[DATA][28] , \resource_in_f[DATA][27] , 
        \resource_in_f[DATA][26] , \resource_in_f[DATA][25] , 
        \resource_in_f[DATA][24] , \resource_in_f[DATA][23] , 
        \resource_in_f[DATA][22] , \resource_in_f[DATA][21] , 
        \resource_in_f[DATA][20] , \resource_in_f[DATA][19] , 
        \resource_in_f[DATA][18] , \resource_in_f[DATA][17] , 
        \resource_in_f[DATA][16] , \resource_in_f[DATA][15] , 
        \resource_in_f[DATA][14] , \resource_in_f[DATA][13] , 
        \resource_in_f[DATA][12] , \resource_in_f[DATA][11] , 
        \resource_in_f[DATA][10] , \resource_in_f[DATA][9] , 
        \resource_in_f[DATA][8] , \resource_in_f[DATA][7] , 
        \resource_in_f[DATA][6] , \resource_in_f[DATA][5] , 
        \resource_in_f[DATA][4] , \resource_in_f[DATA][3] , 
        \resource_in_f[DATA][2] , \resource_in_f[DATA][1] , 
        \resource_in_f[DATA][0] }), .resource_in_b(\resource_in_b[ACK] ), 
    .north_out_f({\north_out_f[REQ] , \north_out_f[DATA][34] , 
        \north_out_f[DATA][33] , \north_out_f[DATA][32] , 
        \north_out_f[DATA][31] , \north_out_f[DATA][30] , 
        \north_out_f[DATA][29] , \north_out_f[DATA][28] , 
        \north_out_f[DATA][27] , \north_out_f[DATA][26] , 
        \north_out_f[DATA][25] , \north_out_f[DATA][24] , 
        \north_out_f[DATA][23] , \north_out_f[DATA][22] , 
        \north_out_f[DATA][21] , \north_out_f[DATA][20] , 
        \north_out_f[DATA][19] , \north_out_f[DATA][18] , 
        \north_out_f[DATA][17] , \north_out_f[DATA][16] , 
        \north_out_f[DATA][15] , \north_out_f[DATA][14] , 
        \north_out_f[DATA][13] , \north_out_f[DATA][12] , 
        \north_out_f[DATA][11] , \north_out_f[DATA][10] , 
        \north_out_f[DATA][9] , \north_out_f[DATA][8] , \north_out_f[DATA][7] , 
        \north_out_f[DATA][6] , \north_out_f[DATA][5] , \north_out_f[DATA][4] , 
        \north_out_f[DATA][3] , \north_out_f[DATA][2] , \north_out_f[DATA][1] , 
        \north_out_f[DATA][0] }), .north_out_b(\north_out_b[ACK] ), 
    .east_out_f({\east_out_f[REQ] , \east_out_f[DATA][34] , 
        \east_out_f[DATA][33] , \east_out_f[DATA][32] , \east_out_f[DATA][31] , 
        \east_out_f[DATA][30] , \east_out_f[DATA][29] , \east_out_f[DATA][28] , 
        \east_out_f[DATA][27] , \east_out_f[DATA][26] , \east_out_f[DATA][25] , 
        \east_out_f[DATA][24] , \east_out_f[DATA][23] , \east_out_f[DATA][22] , 
        \east_out_f[DATA][21] , \east_out_f[DATA][20] , \east_out_f[DATA][19] , 
        \east_out_f[DATA][18] , \east_out_f[DATA][17] , \east_out_f[DATA][16] , 
        \east_out_f[DATA][15] , \east_out_f[DATA][14] , \east_out_f[DATA][13] , 
        \east_out_f[DATA][12] , \east_out_f[DATA][11] , \east_out_f[DATA][10] , 
        \east_out_f[DATA][9] , \east_out_f[DATA][8] , \east_out_f[DATA][7] , 
        \east_out_f[DATA][6] , \east_out_f[DATA][5] , \east_out_f[DATA][4] , 
        \east_out_f[DATA][3] , \east_out_f[DATA][2] , \east_out_f[DATA][1] , 
        \east_out_f[DATA][0] }), .east_out_b(\east_out_b[ACK] ), 
    .south_out_f({\south_out_f[REQ] , \south_out_f[DATA][34] , 
        \south_out_f[DATA][33] , \south_out_f[DATA][32] , 
        \south_out_f[DATA][31] , \south_out_f[DATA][30] , 
        \south_out_f[DATA][29] , \south_out_f[DATA][28] , 
        \south_out_f[DATA][27] , \south_out_f[DATA][26] , 
        \south_out_f[DATA][25] , \south_out_f[DATA][24] , 
        \south_out_f[DATA][23] , \south_out_f[DATA][22] , 
        \south_out_f[DATA][21] , \south_out_f[DATA][20] , 
        \south_out_f[DATA][19] , \south_out_f[DATA][18] , 
        \south_out_f[DATA][17] , \south_out_f[DATA][16] , 
        \south_out_f[DATA][15] , \south_out_f[DATA][14] , 
        \south_out_f[DATA][13] , \south_out_f[DATA][12] , 
        \south_out_f[DATA][11] , \south_out_f[DATA][10] , 
        \south_out_f[DATA][9] , \south_out_f[DATA][8] , \south_out_f[DATA][7] , 
        \south_out_f[DATA][6] , \south_out_f[DATA][5] , \south_out_f[DATA][4] , 
        \south_out_f[DATA][3] , \south_out_f[DATA][2] , \south_out_f[DATA][1] , 
        \south_out_f[DATA][0] }), .south_out_b(\south_out_b[ACK] ), 
    .west_out_f({\west_out_f[REQ] , \west_out_f[DATA][34] , 
        \west_out_f[DATA][33] , \west_out_f[DATA][32] , \west_out_f[DATA][31] , 
        \west_out_f[DATA][30] , \west_out_f[DATA][29] , \west_out_f[DATA][28] , 
        \west_out_f[DATA][27] , \west_out_f[DATA][26] , \west_out_f[DATA][25] , 
        \west_out_f[DATA][24] , \west_out_f[DATA][23] , \west_out_f[DATA][22] , 
        \west_out_f[DATA][21] , \west_out_f[DATA][20] , \west_out_f[DATA][19] , 
        \west_out_f[DATA][18] , \west_out_f[DATA][17] , \west_out_f[DATA][16] , 
        \west_out_f[DATA][15] , \west_out_f[DATA][14] , \west_out_f[DATA][13] , 
        \west_out_f[DATA][12] , \west_out_f[DATA][11] , \west_out_f[DATA][10] , 
        \west_out_f[DATA][9] , \west_out_f[DATA][8] , \west_out_f[DATA][7] , 
        \west_out_f[DATA][6] , \west_out_f[DATA][5] , \west_out_f[DATA][4] , 
        \west_out_f[DATA][3] , \west_out_f[DATA][2] , \west_out_f[DATA][1] , 
        \west_out_f[DATA][0] }), .west_out_b(\west_out_b[ACK] ), 
    .resource_out_f({\resource_out_f[REQ] , \resource_out_f[DATA][34] , 
        \resource_out_f[DATA][33] , \resource_out_f[DATA][32] , 
        \resource_out_f[DATA][31] , \resource_out_f[DATA][30] , 
        \resource_out_f[DATA][29] , \resource_out_f[DATA][28] , 
        \resource_out_f[DATA][27] , \resource_out_f[DATA][26] , 
        \resource_out_f[DATA][25] , \resource_out_f[DATA][24] , 
        \resource_out_f[DATA][23] , \resource_out_f[DATA][22] , 
        \resource_out_f[DATA][21] , \resource_out_f[DATA][20] , 
        \resource_out_f[DATA][19] , \resource_out_f[DATA][18] , 
        \resource_out_f[DATA][17] , \resource_out_f[DATA][16] , 
        \resource_out_f[DATA][15] , \resource_out_f[DATA][14] , 
        \resource_out_f[DATA][13] , \resource_out_f[DATA][12] , 
        \resource_out_f[DATA][11] , \resource_out_f[DATA][10] , 
        \resource_out_f[DATA][9] , \resource_out_f[DATA][8] , 
        \resource_out_f[DATA][7] , \resource_out_f[DATA][6] , 
        \resource_out_f[DATA][5] , \resource_out_f[DATA][4] , 
        \resource_out_f[DATA][3] , \resource_out_f[DATA][2] , 
        \resource_out_f[DATA][1] , \resource_out_f[DATA][0] }), 
    .resource_out_b(\resource_out_b[ACK] ) );
  input preset, \north_in_f[REQ] , \north_in_f[DATA][34] ,
         \north_in_f[DATA][33] , \north_in_f[DATA][32] ,
         \north_in_f[DATA][31] , \north_in_f[DATA][30] ,
         \north_in_f[DATA][29] , \north_in_f[DATA][28] ,
         \north_in_f[DATA][27] , \north_in_f[DATA][26] ,
         \north_in_f[DATA][25] , \north_in_f[DATA][24] ,
         \north_in_f[DATA][23] , \north_in_f[DATA][22] ,
         \north_in_f[DATA][21] , \north_in_f[DATA][20] ,
         \north_in_f[DATA][19] , \north_in_f[DATA][18] ,
         \north_in_f[DATA][17] , \north_in_f[DATA][16] ,
         \north_in_f[DATA][15] , \north_in_f[DATA][14] ,
         \north_in_f[DATA][13] , \north_in_f[DATA][12] ,
         \north_in_f[DATA][11] , \north_in_f[DATA][10] , \north_in_f[DATA][9] ,
         \north_in_f[DATA][8] , \north_in_f[DATA][7] , \north_in_f[DATA][6] ,
         \north_in_f[DATA][5] , \north_in_f[DATA][4] , \north_in_f[DATA][3] ,
         \north_in_f[DATA][2] , \north_in_f[DATA][1] , \north_in_f[DATA][0] ,
         \east_in_f[REQ] , \east_in_f[DATA][34] , \east_in_f[DATA][33] ,
         \east_in_f[DATA][32] , \east_in_f[DATA][31] , \east_in_f[DATA][30] ,
         \east_in_f[DATA][29] , \east_in_f[DATA][28] , \east_in_f[DATA][27] ,
         \east_in_f[DATA][26] , \east_in_f[DATA][25] , \east_in_f[DATA][24] ,
         \east_in_f[DATA][23] , \east_in_f[DATA][22] , \east_in_f[DATA][21] ,
         \east_in_f[DATA][20] , \east_in_f[DATA][19] , \east_in_f[DATA][18] ,
         \east_in_f[DATA][17] , \east_in_f[DATA][16] , \east_in_f[DATA][15] ,
         \east_in_f[DATA][14] , \east_in_f[DATA][13] , \east_in_f[DATA][12] ,
         \east_in_f[DATA][11] , \east_in_f[DATA][10] , \east_in_f[DATA][9] ,
         \east_in_f[DATA][8] , \east_in_f[DATA][7] , \east_in_f[DATA][6] ,
         \east_in_f[DATA][5] , \east_in_f[DATA][4] , \east_in_f[DATA][3] ,
         \east_in_f[DATA][2] , \east_in_f[DATA][1] , \east_in_f[DATA][0] ,
         \south_in_f[REQ] , \south_in_f[DATA][34] , \south_in_f[DATA][33] ,
         \south_in_f[DATA][32] , \south_in_f[DATA][31] ,
         \south_in_f[DATA][30] , \south_in_f[DATA][29] ,
         \south_in_f[DATA][28] , \south_in_f[DATA][27] ,
         \south_in_f[DATA][26] , \south_in_f[DATA][25] ,
         \south_in_f[DATA][24] , \south_in_f[DATA][23] ,
         \south_in_f[DATA][22] , \south_in_f[DATA][21] ,
         \south_in_f[DATA][20] , \south_in_f[DATA][19] ,
         \south_in_f[DATA][18] , \south_in_f[DATA][17] ,
         \south_in_f[DATA][16] , \south_in_f[DATA][15] ,
         \south_in_f[DATA][14] , \south_in_f[DATA][13] ,
         \south_in_f[DATA][12] , \south_in_f[DATA][11] ,
         \south_in_f[DATA][10] , \south_in_f[DATA][9] , \south_in_f[DATA][8] ,
         \south_in_f[DATA][7] , \south_in_f[DATA][6] , \south_in_f[DATA][5] ,
         \south_in_f[DATA][4] , \south_in_f[DATA][3] , \south_in_f[DATA][2] ,
         \south_in_f[DATA][1] , \south_in_f[DATA][0] , \west_in_f[REQ] ,
         \west_in_f[DATA][34] , \west_in_f[DATA][33] , \west_in_f[DATA][32] ,
         \west_in_f[DATA][31] , \west_in_f[DATA][30] , \west_in_f[DATA][29] ,
         \west_in_f[DATA][28] , \west_in_f[DATA][27] , \west_in_f[DATA][26] ,
         \west_in_f[DATA][25] , \west_in_f[DATA][24] , \west_in_f[DATA][23] ,
         \west_in_f[DATA][22] , \west_in_f[DATA][21] , \west_in_f[DATA][20] ,
         \west_in_f[DATA][19] , \west_in_f[DATA][18] , \west_in_f[DATA][17] ,
         \west_in_f[DATA][16] , \west_in_f[DATA][15] , \west_in_f[DATA][14] ,
         \west_in_f[DATA][13] , \west_in_f[DATA][12] , \west_in_f[DATA][11] ,
         \west_in_f[DATA][10] , \west_in_f[DATA][9] , \west_in_f[DATA][8] ,
         \west_in_f[DATA][7] , \west_in_f[DATA][6] , \west_in_f[DATA][5] ,
         \west_in_f[DATA][4] , \west_in_f[DATA][3] , \west_in_f[DATA][2] ,
         \west_in_f[DATA][1] , \west_in_f[DATA][0] , \resource_in_f[REQ] ,
         \resource_in_f[DATA][34] , \resource_in_f[DATA][33] ,
         \resource_in_f[DATA][32] , \resource_in_f[DATA][31] ,
         \resource_in_f[DATA][30] , \resource_in_f[DATA][29] ,
         \resource_in_f[DATA][28] , \resource_in_f[DATA][27] ,
         \resource_in_f[DATA][26] , \resource_in_f[DATA][25] ,
         \resource_in_f[DATA][24] , \resource_in_f[DATA][23] ,
         \resource_in_f[DATA][22] , \resource_in_f[DATA][21] ,
         \resource_in_f[DATA][20] , \resource_in_f[DATA][19] ,
         \resource_in_f[DATA][18] , \resource_in_f[DATA][17] ,
         \resource_in_f[DATA][16] , \resource_in_f[DATA][15] ,
         \resource_in_f[DATA][14] , \resource_in_f[DATA][13] ,
         \resource_in_f[DATA][12] , \resource_in_f[DATA][11] ,
         \resource_in_f[DATA][10] , \resource_in_f[DATA][9] ,
         \resource_in_f[DATA][8] , \resource_in_f[DATA][7] ,
         \resource_in_f[DATA][6] , \resource_in_f[DATA][5] ,
         \resource_in_f[DATA][4] , \resource_in_f[DATA][3] ,
         \resource_in_f[DATA][2] , \resource_in_f[DATA][1] ,
         \resource_in_f[DATA][0] , \north_out_b[ACK] , \east_out_b[ACK] ,
         \south_out_b[ACK] , \west_out_b[ACK] , \resource_out_b[ACK] ;
  output \north_in_b[ACK] , \east_in_b[ACK] , \south_in_b[ACK] ,
         \west_in_b[ACK] , \resource_in_b[ACK] , \north_out_f[REQ] ,
         \north_out_f[DATA][34] , \north_out_f[DATA][33] ,
         \north_out_f[DATA][32] , \north_out_f[DATA][31] ,
         \north_out_f[DATA][30] , \north_out_f[DATA][29] ,
         \north_out_f[DATA][28] , \north_out_f[DATA][27] ,
         \north_out_f[DATA][26] , \north_out_f[DATA][25] ,
         \north_out_f[DATA][24] , \north_out_f[DATA][23] ,
         \north_out_f[DATA][22] , \north_out_f[DATA][21] ,
         \north_out_f[DATA][20] , \north_out_f[DATA][19] ,
         \north_out_f[DATA][18] , \north_out_f[DATA][17] ,
         \north_out_f[DATA][16] , \north_out_f[DATA][15] ,
         \north_out_f[DATA][14] , \north_out_f[DATA][13] ,
         \north_out_f[DATA][12] , \north_out_f[DATA][11] ,
         \north_out_f[DATA][10] , \north_out_f[DATA][9] ,
         \north_out_f[DATA][8] , \north_out_f[DATA][7] ,
         \north_out_f[DATA][6] , \north_out_f[DATA][5] ,
         \north_out_f[DATA][4] , \north_out_f[DATA][3] ,
         \north_out_f[DATA][2] , \north_out_f[DATA][1] ,
         \north_out_f[DATA][0] , \east_out_f[REQ] , \east_out_f[DATA][34] ,
         \east_out_f[DATA][33] , \east_out_f[DATA][32] ,
         \east_out_f[DATA][31] , \east_out_f[DATA][30] ,
         \east_out_f[DATA][29] , \east_out_f[DATA][28] ,
         \east_out_f[DATA][27] , \east_out_f[DATA][26] ,
         \east_out_f[DATA][25] , \east_out_f[DATA][24] ,
         \east_out_f[DATA][23] , \east_out_f[DATA][22] ,
         \east_out_f[DATA][21] , \east_out_f[DATA][20] ,
         \east_out_f[DATA][19] , \east_out_f[DATA][18] ,
         \east_out_f[DATA][17] , \east_out_f[DATA][16] ,
         \east_out_f[DATA][15] , \east_out_f[DATA][14] ,
         \east_out_f[DATA][13] , \east_out_f[DATA][12] ,
         \east_out_f[DATA][11] , \east_out_f[DATA][10] , \east_out_f[DATA][9] ,
         \east_out_f[DATA][8] , \east_out_f[DATA][7] , \east_out_f[DATA][6] ,
         \east_out_f[DATA][5] , \east_out_f[DATA][4] , \east_out_f[DATA][3] ,
         \east_out_f[DATA][2] , \east_out_f[DATA][1] , \east_out_f[DATA][0] ,
         \south_out_f[REQ] , \south_out_f[DATA][34] , \south_out_f[DATA][33] ,
         \south_out_f[DATA][32] , \south_out_f[DATA][31] ,
         \south_out_f[DATA][30] , \south_out_f[DATA][29] ,
         \south_out_f[DATA][28] , \south_out_f[DATA][27] ,
         \south_out_f[DATA][26] , \south_out_f[DATA][25] ,
         \south_out_f[DATA][24] , \south_out_f[DATA][23] ,
         \south_out_f[DATA][22] , \south_out_f[DATA][21] ,
         \south_out_f[DATA][20] , \south_out_f[DATA][19] ,
         \south_out_f[DATA][18] , \south_out_f[DATA][17] ,
         \south_out_f[DATA][16] , \south_out_f[DATA][15] ,
         \south_out_f[DATA][14] , \south_out_f[DATA][13] ,
         \south_out_f[DATA][12] , \south_out_f[DATA][11] ,
         \south_out_f[DATA][10] , \south_out_f[DATA][9] ,
         \south_out_f[DATA][8] , \south_out_f[DATA][7] ,
         \south_out_f[DATA][6] , \south_out_f[DATA][5] ,
         \south_out_f[DATA][4] , \south_out_f[DATA][3] ,
         \south_out_f[DATA][2] , \south_out_f[DATA][1] ,
         \south_out_f[DATA][0] , \west_out_f[REQ] , \west_out_f[DATA][34] ,
         \west_out_f[DATA][33] , \west_out_f[DATA][32] ,
         \west_out_f[DATA][31] , \west_out_f[DATA][30] ,
         \west_out_f[DATA][29] , \west_out_f[DATA][28] ,
         \west_out_f[DATA][27] , \west_out_f[DATA][26] ,
         \west_out_f[DATA][25] , \west_out_f[DATA][24] ,
         \west_out_f[DATA][23] , \west_out_f[DATA][22] ,
         \west_out_f[DATA][21] , \west_out_f[DATA][20] ,
         \west_out_f[DATA][19] , \west_out_f[DATA][18] ,
         \west_out_f[DATA][17] , \west_out_f[DATA][16] ,
         \west_out_f[DATA][15] , \west_out_f[DATA][14] ,
         \west_out_f[DATA][13] , \west_out_f[DATA][12] ,
         \west_out_f[DATA][11] , \west_out_f[DATA][10] , \west_out_f[DATA][9] ,
         \west_out_f[DATA][8] , \west_out_f[DATA][7] , \west_out_f[DATA][6] ,
         \west_out_f[DATA][5] , \west_out_f[DATA][4] , \west_out_f[DATA][3] ,
         \west_out_f[DATA][2] , \west_out_f[DATA][1] , \west_out_f[DATA][0] ,
         \resource_out_f[REQ] , \resource_out_f[DATA][34] ,
         \resource_out_f[DATA][33] , \resource_out_f[DATA][32] ,
         \resource_out_f[DATA][31] , \resource_out_f[DATA][30] ,
         \resource_out_f[DATA][29] , \resource_out_f[DATA][28] ,
         \resource_out_f[DATA][27] , \resource_out_f[DATA][26] ,
         \resource_out_f[DATA][25] , \resource_out_f[DATA][24] ,
         \resource_out_f[DATA][23] , \resource_out_f[DATA][22] ,
         \resource_out_f[DATA][21] , \resource_out_f[DATA][20] ,
         \resource_out_f[DATA][19] , \resource_out_f[DATA][18] ,
         \resource_out_f[DATA][17] , \resource_out_f[DATA][16] ,
         \resource_out_f[DATA][15] , \resource_out_f[DATA][14] ,
         \resource_out_f[DATA][13] , \resource_out_f[DATA][12] ,
         \resource_out_f[DATA][11] , \resource_out_f[DATA][10] ,
         \resource_out_f[DATA][9] , \resource_out_f[DATA][8] ,
         \resource_out_f[DATA][7] , \resource_out_f[DATA][6] ,
         \resource_out_f[DATA][5] , \resource_out_f[DATA][4] ,
         \resource_out_f[DATA][3] , \resource_out_f[DATA][2] ,
         \resource_out_f[DATA][1] , \resource_out_f[DATA][0] ;
  wire   \north_hpu_f[REQ] , \north_hpu_f[DATA][34] , \north_hpu_f[DATA][33] ,
         \north_hpu_f[DATA][32] , \north_hpu_f[DATA][31] ,
         \north_hpu_f[DATA][30] , \north_hpu_f[DATA][29] ,
         \north_hpu_f[DATA][28] , \north_hpu_f[DATA][27] ,
         \north_hpu_f[DATA][26] , \north_hpu_f[DATA][25] ,
         \north_hpu_f[DATA][24] , \north_hpu_f[DATA][23] ,
         \north_hpu_f[DATA][22] , \north_hpu_f[DATA][21] ,
         \north_hpu_f[DATA][20] , \north_hpu_f[DATA][19] ,
         \north_hpu_f[DATA][18] , \north_hpu_f[DATA][17] ,
         \north_hpu_f[DATA][16] , \north_hpu_f[DATA][15] ,
         \north_hpu_f[DATA][14] , \north_hpu_f[DATA][13] ,
         \north_hpu_f[DATA][12] , \north_hpu_f[DATA][11] ,
         \north_hpu_f[DATA][10] , \north_hpu_f[DATA][9] ,
         \north_hpu_f[DATA][8] , \north_hpu_f[DATA][7] ,
         \north_hpu_f[DATA][6] , \north_hpu_f[DATA][5] ,
         \north_hpu_f[DATA][4] , \north_hpu_f[DATA][3] ,
         \north_hpu_f[DATA][2] , \north_hpu_f[DATA][1] ,
         \north_hpu_f[DATA][0] , \north_hpu_b[ACK] , \south_hpu_f[REQ] ,
         \south_hpu_f[DATA][34] , \south_hpu_f[DATA][33] ,
         \south_hpu_f[DATA][32] , \south_hpu_f[DATA][31] ,
         \south_hpu_f[DATA][30] , \south_hpu_f[DATA][29] ,
         \south_hpu_f[DATA][28] , \south_hpu_f[DATA][27] ,
         \south_hpu_f[DATA][26] , \south_hpu_f[DATA][25] ,
         \south_hpu_f[DATA][24] , \south_hpu_f[DATA][23] ,
         \south_hpu_f[DATA][22] , \south_hpu_f[DATA][21] ,
         \south_hpu_f[DATA][20] , \south_hpu_f[DATA][19] ,
         \south_hpu_f[DATA][18] , \south_hpu_f[DATA][17] ,
         \south_hpu_f[DATA][16] , \south_hpu_f[DATA][15] ,
         \south_hpu_f[DATA][14] , \south_hpu_f[DATA][13] ,
         \south_hpu_f[DATA][12] , \south_hpu_f[DATA][11] ,
         \south_hpu_f[DATA][10] , \south_hpu_f[DATA][9] ,
         \south_hpu_f[DATA][8] , \south_hpu_f[DATA][7] ,
         \south_hpu_f[DATA][6] , \south_hpu_f[DATA][5] ,
         \south_hpu_f[DATA][4] , \south_hpu_f[DATA][3] ,
         \south_hpu_f[DATA][2] , \south_hpu_f[DATA][1] ,
         \south_hpu_f[DATA][0] , \south_hpu_b[ACK] , \east_hpu_f[REQ] ,
         \east_hpu_f[DATA][34] , \east_hpu_f[DATA][33] ,
         \east_hpu_f[DATA][32] , \east_hpu_f[DATA][31] ,
         \east_hpu_f[DATA][30] , \east_hpu_f[DATA][29] ,
         \east_hpu_f[DATA][28] , \east_hpu_f[DATA][27] ,
         \east_hpu_f[DATA][26] , \east_hpu_f[DATA][25] ,
         \east_hpu_f[DATA][24] , \east_hpu_f[DATA][23] ,
         \east_hpu_f[DATA][22] , \east_hpu_f[DATA][21] ,
         \east_hpu_f[DATA][20] , \east_hpu_f[DATA][19] ,
         \east_hpu_f[DATA][18] , \east_hpu_f[DATA][17] ,
         \east_hpu_f[DATA][16] , \east_hpu_f[DATA][15] ,
         \east_hpu_f[DATA][14] , \east_hpu_f[DATA][13] ,
         \east_hpu_f[DATA][12] , \east_hpu_f[DATA][11] ,
         \east_hpu_f[DATA][10] , \east_hpu_f[DATA][9] , \east_hpu_f[DATA][8] ,
         \east_hpu_f[DATA][7] , \east_hpu_f[DATA][6] , \east_hpu_f[DATA][5] ,
         \east_hpu_f[DATA][4] , \east_hpu_f[DATA][3] , \east_hpu_f[DATA][2] ,
         \east_hpu_f[DATA][1] , \east_hpu_f[DATA][0] , \east_hpu_b[ACK] ,
         \west_hpu_f[REQ] , \west_hpu_f[DATA][34] , \west_hpu_f[DATA][33] ,
         \west_hpu_f[DATA][32] , \west_hpu_f[DATA][31] ,
         \west_hpu_f[DATA][30] , \west_hpu_f[DATA][29] ,
         \west_hpu_f[DATA][28] , \west_hpu_f[DATA][27] ,
         \west_hpu_f[DATA][26] , \west_hpu_f[DATA][25] ,
         \west_hpu_f[DATA][24] , \west_hpu_f[DATA][23] ,
         \west_hpu_f[DATA][22] , \west_hpu_f[DATA][21] ,
         \west_hpu_f[DATA][20] , \west_hpu_f[DATA][19] ,
         \west_hpu_f[DATA][18] , \west_hpu_f[DATA][17] ,
         \west_hpu_f[DATA][16] , \west_hpu_f[DATA][15] ,
         \west_hpu_f[DATA][14] , \west_hpu_f[DATA][13] ,
         \west_hpu_f[DATA][12] , \west_hpu_f[DATA][11] ,
         \west_hpu_f[DATA][10] , \west_hpu_f[DATA][9] , \west_hpu_f[DATA][8] ,
         \west_hpu_f[DATA][7] , \west_hpu_f[DATA][6] , \west_hpu_f[DATA][5] ,
         \west_hpu_f[DATA][4] , \west_hpu_f[DATA][3] , \west_hpu_f[DATA][2] ,
         \west_hpu_f[DATA][1] , \west_hpu_f[DATA][0] , \west_hpu_b[ACK] ,
         \resource_hpu_f[REQ] , \resource_hpu_f[DATA][34] ,
         \resource_hpu_f[DATA][33] , \resource_hpu_f[DATA][32] ,
         \resource_hpu_f[DATA][31] , \resource_hpu_f[DATA][30] ,
         \resource_hpu_f[DATA][29] , \resource_hpu_f[DATA][28] ,
         \resource_hpu_f[DATA][27] , \resource_hpu_f[DATA][26] ,
         \resource_hpu_f[DATA][25] , \resource_hpu_f[DATA][24] ,
         \resource_hpu_f[DATA][23] , \resource_hpu_f[DATA][22] ,
         \resource_hpu_f[DATA][21] , \resource_hpu_f[DATA][20] ,
         \resource_hpu_f[DATA][19] , \resource_hpu_f[DATA][18] ,
         \resource_hpu_f[DATA][17] , \resource_hpu_f[DATA][16] ,
         \resource_hpu_f[DATA][15] , \resource_hpu_f[DATA][14] ,
         \resource_hpu_f[DATA][13] , \resource_hpu_f[DATA][12] ,
         \resource_hpu_f[DATA][11] , \resource_hpu_f[DATA][10] ,
         \resource_hpu_f[DATA][9] , \resource_hpu_f[DATA][8] ,
         \resource_hpu_f[DATA][7] , \resource_hpu_f[DATA][6] ,
         \resource_hpu_f[DATA][5] , \resource_hpu_f[DATA][4] ,
         \resource_hpu_f[DATA][3] , \resource_hpu_f[DATA][2] ,
         \resource_hpu_f[DATA][1] , \resource_hpu_f[DATA][0] ,
         \resource_hpu_b[ACK] , \chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] ,
         \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] ,
         \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] ,
         \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] ,
         \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] ,
         \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] ,
         \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] ,
         \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] ,
         \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] ,
         \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] ,
         \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] ,
         \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] ,
         \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] ,
         \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] ,
         \chs_in_f[4][DATA][7] , \chs_in_f[4][DATA][6] ,
         \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] ,
         \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] ,
         \chs_in_f[4][DATA][1] , \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] ,
         \chs_in_f[3][DATA][34] , \chs_in_f[3][DATA][33] ,
         \chs_in_f[3][DATA][32] , \chs_in_f[3][DATA][31] ,
         \chs_in_f[3][DATA][30] , \chs_in_f[3][DATA][29] ,
         \chs_in_f[3][DATA][28] , \chs_in_f[3][DATA][27] ,
         \chs_in_f[3][DATA][26] , \chs_in_f[3][DATA][25] ,
         \chs_in_f[3][DATA][24] , \chs_in_f[3][DATA][23] ,
         \chs_in_f[3][DATA][22] , \chs_in_f[3][DATA][21] ,
         \chs_in_f[3][DATA][20] , \chs_in_f[3][DATA][19] ,
         \chs_in_f[3][DATA][18] , \chs_in_f[3][DATA][17] ,
         \chs_in_f[3][DATA][16] , \chs_in_f[3][DATA][15] ,
         \chs_in_f[3][DATA][14] , \chs_in_f[3][DATA][13] ,
         \chs_in_f[3][DATA][12] , \chs_in_f[3][DATA][11] ,
         \chs_in_f[3][DATA][10] , \chs_in_f[3][DATA][9] ,
         \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] ,
         \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] ,
         \chs_in_f[3][DATA][4] , \chs_in_f[3][DATA][3] ,
         \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] ,
         \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] ,
         \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] ,
         \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] ,
         \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] ,
         \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] ,
         \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] ,
         \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] ,
         \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] ,
         \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] ,
         \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] ,
         \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] ,
         \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] ,
         \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] ,
         \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] ,
         \chs_in_f[2][DATA][7] , \chs_in_f[2][DATA][6] ,
         \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] ,
         \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] ,
         \chs_in_f[2][DATA][1] , \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] ,
         \chs_in_f[1][DATA][34] , \chs_in_f[1][DATA][33] ,
         \chs_in_f[1][DATA][32] , \chs_in_f[1][DATA][31] ,
         \chs_in_f[1][DATA][30] , \chs_in_f[1][DATA][29] ,
         \chs_in_f[1][DATA][28] , \chs_in_f[1][DATA][27] ,
         \chs_in_f[1][DATA][26] , \chs_in_f[1][DATA][25] ,
         \chs_in_f[1][DATA][24] , \chs_in_f[1][DATA][23] ,
         \chs_in_f[1][DATA][22] , \chs_in_f[1][DATA][21] ,
         \chs_in_f[1][DATA][20] , \chs_in_f[1][DATA][19] ,
         \chs_in_f[1][DATA][18] , \chs_in_f[1][DATA][17] ,
         \chs_in_f[1][DATA][16] , \chs_in_f[1][DATA][15] ,
         \chs_in_f[1][DATA][14] , \chs_in_f[1][DATA][13] ,
         \chs_in_f[1][DATA][12] , \chs_in_f[1][DATA][11] ,
         \chs_in_f[1][DATA][10] , \chs_in_f[1][DATA][9] ,
         \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] ,
         \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] ,
         \chs_in_f[1][DATA][4] , \chs_in_f[1][DATA][3] ,
         \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] ,
         \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] ,
         \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] ,
         \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] ,
         \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] ,
         \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] ,
         \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] ,
         \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] ,
         \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] ,
         \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] ,
         \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] ,
         \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] ,
         \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] ,
         \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] ,
         \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] ,
         \chs_in_f[0][DATA][7] , \chs_in_f[0][DATA][6] ,
         \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] ,
         \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] ,
         \chs_in_f[0][DATA][1] , \chs_in_f[0][DATA][0] , \chs_in_b[4][ACK] ,
         \chs_in_b[3][ACK] , \chs_in_b[2][ACK] , \chs_in_b[1][ACK] ,
         \chs_in_b[0][ACK] , \switch_sel[4][4] , \switch_sel[4][3] ,
         \switch_sel[4][2] , \switch_sel[4][1] , \switch_sel[4][0] ,
         \switch_sel[3][4] , \switch_sel[3][3] , \switch_sel[3][2] ,
         \switch_sel[3][1] , \switch_sel[3][0] , \switch_sel[2][4] ,
         \switch_sel[2][3] , \switch_sel[2][2] , \switch_sel[2][1] ,
         \switch_sel[2][0] , \switch_sel[1][4] , \switch_sel[1][3] ,
         \switch_sel[1][2] , \switch_sel[1][1] , \switch_sel[1][0] ,
         \switch_sel[0][4] , \switch_sel[0][3] , \switch_sel[0][2] ,
         \switch_sel[0][1] , \switch_sel[0][0] , n2, n3;

  channel_latch_1_xxxxxxxxx_0 north_in_latch ( .preset(n3), .left_in({
        \north_in_f[REQ] , \north_in_f[DATA][34] , \north_in_f[DATA][33] , 
        \north_in_f[DATA][32] , \north_in_f[DATA][31] , \north_in_f[DATA][30] , 
        \north_in_f[DATA][29] , \north_in_f[DATA][28] , \north_in_f[DATA][27] , 
        \north_in_f[DATA][26] , \north_in_f[DATA][25] , \north_in_f[DATA][24] , 
        \north_in_f[DATA][23] , \north_in_f[DATA][22] , \north_in_f[DATA][21] , 
        \north_in_f[DATA][20] , \north_in_f[DATA][19] , \north_in_f[DATA][18] , 
        \north_in_f[DATA][17] , \north_in_f[DATA][16] , \north_in_f[DATA][15] , 
        \north_in_f[DATA][14] , \north_in_f[DATA][13] , \north_in_f[DATA][12] , 
        \north_in_f[DATA][11] , \north_in_f[DATA][10] , \north_in_f[DATA][9] , 
        \north_in_f[DATA][8] , \north_in_f[DATA][7] , \north_in_f[DATA][6] , 
        \north_in_f[DATA][5] , \north_in_f[DATA][4] , \north_in_f[DATA][3] , 
        \north_in_f[DATA][2] , \north_in_f[DATA][1] , \north_in_f[DATA][0] }), 
        .left_out(\north_in_b[ACK] ), .right_out({\north_hpu_f[REQ] , 
        \north_hpu_f[DATA][34] , \north_hpu_f[DATA][33] , 
        \north_hpu_f[DATA][32] , \north_hpu_f[DATA][31] , 
        \north_hpu_f[DATA][30] , \north_hpu_f[DATA][29] , 
        \north_hpu_f[DATA][28] , \north_hpu_f[DATA][27] , 
        \north_hpu_f[DATA][26] , \north_hpu_f[DATA][25] , 
        \north_hpu_f[DATA][24] , \north_hpu_f[DATA][23] , 
        \north_hpu_f[DATA][22] , \north_hpu_f[DATA][21] , 
        \north_hpu_f[DATA][20] , \north_hpu_f[DATA][19] , 
        \north_hpu_f[DATA][18] , \north_hpu_f[DATA][17] , 
        \north_hpu_f[DATA][16] , \north_hpu_f[DATA][15] , 
        \north_hpu_f[DATA][14] , \north_hpu_f[DATA][13] , 
        \north_hpu_f[DATA][12] , \north_hpu_f[DATA][11] , 
        \north_hpu_f[DATA][10] , \north_hpu_f[DATA][9] , 
        \north_hpu_f[DATA][8] , \north_hpu_f[DATA][7] , \north_hpu_f[DATA][6] , 
        \north_hpu_f[DATA][5] , \north_hpu_f[DATA][4] , \north_hpu_f[DATA][3] , 
        \north_hpu_f[DATA][2] , \north_hpu_f[DATA][1] , \north_hpu_f[DATA][0] }), .right_in(\north_hpu_b[ACK] ) );
  channel_latch_1_xxxxxxxxx_39 south_in_latch ( .preset(n3), .left_in({
        \south_in_f[REQ] , \south_in_f[DATA][34] , \south_in_f[DATA][33] , 
        \south_in_f[DATA][32] , \south_in_f[DATA][31] , \south_in_f[DATA][30] , 
        \south_in_f[DATA][29] , \south_in_f[DATA][28] , \south_in_f[DATA][27] , 
        \south_in_f[DATA][26] , \south_in_f[DATA][25] , \south_in_f[DATA][24] , 
        \south_in_f[DATA][23] , \south_in_f[DATA][22] , \south_in_f[DATA][21] , 
        \south_in_f[DATA][20] , \south_in_f[DATA][19] , \south_in_f[DATA][18] , 
        \south_in_f[DATA][17] , \south_in_f[DATA][16] , \south_in_f[DATA][15] , 
        \south_in_f[DATA][14] , \south_in_f[DATA][13] , \south_in_f[DATA][12] , 
        \south_in_f[DATA][11] , \south_in_f[DATA][10] , \south_in_f[DATA][9] , 
        \south_in_f[DATA][8] , \south_in_f[DATA][7] , \south_in_f[DATA][6] , 
        \south_in_f[DATA][5] , \south_in_f[DATA][4] , \south_in_f[DATA][3] , 
        \south_in_f[DATA][2] , \south_in_f[DATA][1] , \south_in_f[DATA][0] }), 
        .left_out(\south_in_b[ACK] ), .right_out({\south_hpu_f[REQ] , 
        \south_hpu_f[DATA][34] , \south_hpu_f[DATA][33] , 
        \south_hpu_f[DATA][32] , \south_hpu_f[DATA][31] , 
        \south_hpu_f[DATA][30] , \south_hpu_f[DATA][29] , 
        \south_hpu_f[DATA][28] , \south_hpu_f[DATA][27] , 
        \south_hpu_f[DATA][26] , \south_hpu_f[DATA][25] , 
        \south_hpu_f[DATA][24] , \south_hpu_f[DATA][23] , 
        \south_hpu_f[DATA][22] , \south_hpu_f[DATA][21] , 
        \south_hpu_f[DATA][20] , \south_hpu_f[DATA][19] , 
        \south_hpu_f[DATA][18] , \south_hpu_f[DATA][17] , 
        \south_hpu_f[DATA][16] , \south_hpu_f[DATA][15] , 
        \south_hpu_f[DATA][14] , \south_hpu_f[DATA][13] , 
        \south_hpu_f[DATA][12] , \south_hpu_f[DATA][11] , 
        \south_hpu_f[DATA][10] , \south_hpu_f[DATA][9] , 
        \south_hpu_f[DATA][8] , \south_hpu_f[DATA][7] , \south_hpu_f[DATA][6] , 
        \south_hpu_f[DATA][5] , \south_hpu_f[DATA][4] , \south_hpu_f[DATA][3] , 
        \south_hpu_f[DATA][2] , \south_hpu_f[DATA][1] , \south_hpu_f[DATA][0] }), .right_in(\south_hpu_b[ACK] ) );
  channel_latch_1_xxxxxxxxx_38 east_in_latch ( .preset(n3), .left_in({
        \east_in_f[REQ] , \east_in_f[DATA][34] , \east_in_f[DATA][33] , 
        \east_in_f[DATA][32] , \east_in_f[DATA][31] , \east_in_f[DATA][30] , 
        \east_in_f[DATA][29] , \east_in_f[DATA][28] , \east_in_f[DATA][27] , 
        \east_in_f[DATA][26] , \east_in_f[DATA][25] , \east_in_f[DATA][24] , 
        \east_in_f[DATA][23] , \east_in_f[DATA][22] , \east_in_f[DATA][21] , 
        \east_in_f[DATA][20] , \east_in_f[DATA][19] , \east_in_f[DATA][18] , 
        \east_in_f[DATA][17] , \east_in_f[DATA][16] , \east_in_f[DATA][15] , 
        \east_in_f[DATA][14] , \east_in_f[DATA][13] , \east_in_f[DATA][12] , 
        \east_in_f[DATA][11] , \east_in_f[DATA][10] , \east_in_f[DATA][9] , 
        \east_in_f[DATA][8] , \east_in_f[DATA][7] , \east_in_f[DATA][6] , 
        \east_in_f[DATA][5] , \east_in_f[DATA][4] , \east_in_f[DATA][3] , 
        \east_in_f[DATA][2] , \east_in_f[DATA][1] , \east_in_f[DATA][0] }), 
        .left_out(\east_in_b[ACK] ), .right_out({\east_hpu_f[REQ] , 
        \east_hpu_f[DATA][34] , \east_hpu_f[DATA][33] , \east_hpu_f[DATA][32] , 
        \east_hpu_f[DATA][31] , \east_hpu_f[DATA][30] , \east_hpu_f[DATA][29] , 
        \east_hpu_f[DATA][28] , \east_hpu_f[DATA][27] , \east_hpu_f[DATA][26] , 
        \east_hpu_f[DATA][25] , \east_hpu_f[DATA][24] , \east_hpu_f[DATA][23] , 
        \east_hpu_f[DATA][22] , \east_hpu_f[DATA][21] , \east_hpu_f[DATA][20] , 
        \east_hpu_f[DATA][19] , \east_hpu_f[DATA][18] , \east_hpu_f[DATA][17] , 
        \east_hpu_f[DATA][16] , \east_hpu_f[DATA][15] , \east_hpu_f[DATA][14] , 
        \east_hpu_f[DATA][13] , \east_hpu_f[DATA][12] , \east_hpu_f[DATA][11] , 
        \east_hpu_f[DATA][10] , \east_hpu_f[DATA][9] , \east_hpu_f[DATA][8] , 
        \east_hpu_f[DATA][7] , \east_hpu_f[DATA][6] , \east_hpu_f[DATA][5] , 
        \east_hpu_f[DATA][4] , \east_hpu_f[DATA][3] , \east_hpu_f[DATA][2] , 
        \east_hpu_f[DATA][1] , \east_hpu_f[DATA][0] }), .right_in(
        \east_hpu_b[ACK] ) );
  channel_latch_1_xxxxxxxxx_37 west_in_latch ( .preset(n3), .left_in({
        \west_in_f[REQ] , \west_in_f[DATA][34] , \west_in_f[DATA][33] , 
        \west_in_f[DATA][32] , \west_in_f[DATA][31] , \west_in_f[DATA][30] , 
        \west_in_f[DATA][29] , \west_in_f[DATA][28] , \west_in_f[DATA][27] , 
        \west_in_f[DATA][26] , \west_in_f[DATA][25] , \west_in_f[DATA][24] , 
        \west_in_f[DATA][23] , \west_in_f[DATA][22] , \west_in_f[DATA][21] , 
        \west_in_f[DATA][20] , \west_in_f[DATA][19] , \west_in_f[DATA][18] , 
        \west_in_f[DATA][17] , \west_in_f[DATA][16] , \west_in_f[DATA][15] , 
        \west_in_f[DATA][14] , \west_in_f[DATA][13] , \west_in_f[DATA][12] , 
        \west_in_f[DATA][11] , \west_in_f[DATA][10] , \west_in_f[DATA][9] , 
        \west_in_f[DATA][8] , \west_in_f[DATA][7] , \west_in_f[DATA][6] , 
        \west_in_f[DATA][5] , \west_in_f[DATA][4] , \west_in_f[DATA][3] , 
        \west_in_f[DATA][2] , \west_in_f[DATA][1] , \west_in_f[DATA][0] }), 
        .left_out(\west_in_b[ACK] ), .right_out({\west_hpu_f[REQ] , 
        \west_hpu_f[DATA][34] , \west_hpu_f[DATA][33] , \west_hpu_f[DATA][32] , 
        \west_hpu_f[DATA][31] , \west_hpu_f[DATA][30] , \west_hpu_f[DATA][29] , 
        \west_hpu_f[DATA][28] , \west_hpu_f[DATA][27] , \west_hpu_f[DATA][26] , 
        \west_hpu_f[DATA][25] , \west_hpu_f[DATA][24] , \west_hpu_f[DATA][23] , 
        \west_hpu_f[DATA][22] , \west_hpu_f[DATA][21] , \west_hpu_f[DATA][20] , 
        \west_hpu_f[DATA][19] , \west_hpu_f[DATA][18] , \west_hpu_f[DATA][17] , 
        \west_hpu_f[DATA][16] , \west_hpu_f[DATA][15] , \west_hpu_f[DATA][14] , 
        \west_hpu_f[DATA][13] , \west_hpu_f[DATA][12] , \west_hpu_f[DATA][11] , 
        \west_hpu_f[DATA][10] , \west_hpu_f[DATA][9] , \west_hpu_f[DATA][8] , 
        \west_hpu_f[DATA][7] , \west_hpu_f[DATA][6] , \west_hpu_f[DATA][5] , 
        \west_hpu_f[DATA][4] , \west_hpu_f[DATA][3] , \west_hpu_f[DATA][2] , 
        \west_hpu_f[DATA][1] , \west_hpu_f[DATA][0] }), .right_in(
        \west_hpu_b[ACK] ) );
  channel_latch_1_xxxxxxxxx_36 resource_in_latch ( .preset(n3), .left_in({
        \resource_in_f[REQ] , \resource_in_f[DATA][34] , 
        \resource_in_f[DATA][33] , \resource_in_f[DATA][32] , 
        \resource_in_f[DATA][31] , \resource_in_f[DATA][30] , 
        \resource_in_f[DATA][29] , \resource_in_f[DATA][28] , 
        \resource_in_f[DATA][27] , \resource_in_f[DATA][26] , 
        \resource_in_f[DATA][25] , \resource_in_f[DATA][24] , 
        \resource_in_f[DATA][23] , \resource_in_f[DATA][22] , 
        \resource_in_f[DATA][21] , \resource_in_f[DATA][20] , 
        \resource_in_f[DATA][19] , \resource_in_f[DATA][18] , 
        \resource_in_f[DATA][17] , \resource_in_f[DATA][16] , 
        \resource_in_f[DATA][15] , \resource_in_f[DATA][14] , 
        \resource_in_f[DATA][13] , \resource_in_f[DATA][12] , 
        \resource_in_f[DATA][11] , \resource_in_f[DATA][10] , 
        \resource_in_f[DATA][9] , \resource_in_f[DATA][8] , 
        \resource_in_f[DATA][7] , \resource_in_f[DATA][6] , 
        \resource_in_f[DATA][5] , \resource_in_f[DATA][4] , 
        \resource_in_f[DATA][3] , \resource_in_f[DATA][2] , 
        \resource_in_f[DATA][1] , \resource_in_f[DATA][0] }), .left_out(
        \resource_in_b[ACK] ), .right_out({\resource_hpu_f[REQ] , 
        \resource_hpu_f[DATA][34] , \resource_hpu_f[DATA][33] , 
        \resource_hpu_f[DATA][32] , \resource_hpu_f[DATA][31] , 
        \resource_hpu_f[DATA][30] , \resource_hpu_f[DATA][29] , 
        \resource_hpu_f[DATA][28] , \resource_hpu_f[DATA][27] , 
        \resource_hpu_f[DATA][26] , \resource_hpu_f[DATA][25] , 
        \resource_hpu_f[DATA][24] , \resource_hpu_f[DATA][23] , 
        \resource_hpu_f[DATA][22] , \resource_hpu_f[DATA][21] , 
        \resource_hpu_f[DATA][20] , \resource_hpu_f[DATA][19] , 
        \resource_hpu_f[DATA][18] , \resource_hpu_f[DATA][17] , 
        \resource_hpu_f[DATA][16] , \resource_hpu_f[DATA][15] , 
        \resource_hpu_f[DATA][14] , \resource_hpu_f[DATA][13] , 
        \resource_hpu_f[DATA][12] , \resource_hpu_f[DATA][11] , 
        \resource_hpu_f[DATA][10] , \resource_hpu_f[DATA][9] , 
        \resource_hpu_f[DATA][8] , \resource_hpu_f[DATA][7] , 
        \resource_hpu_f[DATA][6] , \resource_hpu_f[DATA][5] , 
        \resource_hpu_f[DATA][4] , \resource_hpu_f[DATA][3] , 
        \resource_hpu_f[DATA][2] , \resource_hpu_f[DATA][1] , 
        \resource_hpu_f[DATA][0] }), .right_in(\resource_hpu_b[ACK] ) );
  hpu_0_0_0 north_hpu ( .preset(n2), .chan_in_f({\north_hpu_f[REQ] , 
        \north_hpu_f[DATA][34] , \north_hpu_f[DATA][33] , 
        \north_hpu_f[DATA][32] , \north_hpu_f[DATA][31] , 
        \north_hpu_f[DATA][30] , \north_hpu_f[DATA][29] , 
        \north_hpu_f[DATA][28] , \north_hpu_f[DATA][27] , 
        \north_hpu_f[DATA][26] , \north_hpu_f[DATA][25] , 
        \north_hpu_f[DATA][24] , \north_hpu_f[DATA][23] , 
        \north_hpu_f[DATA][22] , \north_hpu_f[DATA][21] , 
        \north_hpu_f[DATA][20] , \north_hpu_f[DATA][19] , 
        \north_hpu_f[DATA][18] , \north_hpu_f[DATA][17] , 
        \north_hpu_f[DATA][16] , \north_hpu_f[DATA][15] , 
        \north_hpu_f[DATA][14] , \north_hpu_f[DATA][13] , 
        \north_hpu_f[DATA][12] , \north_hpu_f[DATA][11] , 
        \north_hpu_f[DATA][10] , \north_hpu_f[DATA][9] , 
        \north_hpu_f[DATA][8] , \north_hpu_f[DATA][7] , \north_hpu_f[DATA][6] , 
        \north_hpu_f[DATA][5] , \north_hpu_f[DATA][4] , \north_hpu_f[DATA][3] , 
        \north_hpu_f[DATA][2] , \north_hpu_f[DATA][1] , \north_hpu_f[DATA][0] }), .chan_in_b(\north_hpu_b[ACK] ), .chan_out_f({\chs_in_f[0][REQ] , 
        \chs_in_f[0][DATA][34] , \chs_in_f[0][DATA][33] , 
        \chs_in_f[0][DATA][32] , \chs_in_f[0][DATA][31] , 
        \chs_in_f[0][DATA][30] , \chs_in_f[0][DATA][29] , 
        \chs_in_f[0][DATA][28] , \chs_in_f[0][DATA][27] , 
        \chs_in_f[0][DATA][26] , \chs_in_f[0][DATA][25] , 
        \chs_in_f[0][DATA][24] , \chs_in_f[0][DATA][23] , 
        \chs_in_f[0][DATA][22] , \chs_in_f[0][DATA][21] , 
        \chs_in_f[0][DATA][20] , \chs_in_f[0][DATA][19] , 
        \chs_in_f[0][DATA][18] , \chs_in_f[0][DATA][17] , 
        \chs_in_f[0][DATA][16] , \chs_in_f[0][DATA][15] , 
        \chs_in_f[0][DATA][14] , \chs_in_f[0][DATA][13] , 
        \chs_in_f[0][DATA][12] , \chs_in_f[0][DATA][11] , 
        \chs_in_f[0][DATA][10] , \chs_in_f[0][DATA][9] , 
        \chs_in_f[0][DATA][8] , \chs_in_f[0][DATA][7] , \chs_in_f[0][DATA][6] , 
        \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] , \chs_in_f[0][DATA][3] , 
        \chs_in_f[0][DATA][2] , \chs_in_f[0][DATA][1] , \chs_in_f[0][DATA][0] }), .chan_out_b(\chs_in_b[0][ACK] ), .sel({\switch_sel[0][4] , 
        \switch_sel[0][3] , \switch_sel[0][2] , \switch_sel[0][1] , 
        \switch_sel[0][0] }) );
  hpu_0_2_0 south_hpu ( .preset(n2), .chan_in_f({\south_hpu_f[REQ] , 
        \south_hpu_f[DATA][34] , \south_hpu_f[DATA][33] , 
        \south_hpu_f[DATA][32] , \south_hpu_f[DATA][31] , 
        \south_hpu_f[DATA][30] , \south_hpu_f[DATA][29] , 
        \south_hpu_f[DATA][28] , \south_hpu_f[DATA][27] , 
        \south_hpu_f[DATA][26] , \south_hpu_f[DATA][25] , 
        \south_hpu_f[DATA][24] , \south_hpu_f[DATA][23] , 
        \south_hpu_f[DATA][22] , \south_hpu_f[DATA][21] , 
        \south_hpu_f[DATA][20] , \south_hpu_f[DATA][19] , 
        \south_hpu_f[DATA][18] , \south_hpu_f[DATA][17] , 
        \south_hpu_f[DATA][16] , \south_hpu_f[DATA][15] , 
        \south_hpu_f[DATA][14] , \south_hpu_f[DATA][13] , 
        \south_hpu_f[DATA][12] , \south_hpu_f[DATA][11] , 
        \south_hpu_f[DATA][10] , \south_hpu_f[DATA][9] , 
        \south_hpu_f[DATA][8] , \south_hpu_f[DATA][7] , \south_hpu_f[DATA][6] , 
        \south_hpu_f[DATA][5] , \south_hpu_f[DATA][4] , \south_hpu_f[DATA][3] , 
        \south_hpu_f[DATA][2] , \south_hpu_f[DATA][1] , \south_hpu_f[DATA][0] }), .chan_in_b(\south_hpu_b[ACK] ), .chan_out_f({\chs_in_f[2][REQ] , 
        \chs_in_f[2][DATA][34] , \chs_in_f[2][DATA][33] , 
        \chs_in_f[2][DATA][32] , \chs_in_f[2][DATA][31] , 
        \chs_in_f[2][DATA][30] , \chs_in_f[2][DATA][29] , 
        \chs_in_f[2][DATA][28] , \chs_in_f[2][DATA][27] , 
        \chs_in_f[2][DATA][26] , \chs_in_f[2][DATA][25] , 
        \chs_in_f[2][DATA][24] , \chs_in_f[2][DATA][23] , 
        \chs_in_f[2][DATA][22] , \chs_in_f[2][DATA][21] , 
        \chs_in_f[2][DATA][20] , \chs_in_f[2][DATA][19] , 
        \chs_in_f[2][DATA][18] , \chs_in_f[2][DATA][17] , 
        \chs_in_f[2][DATA][16] , \chs_in_f[2][DATA][15] , 
        \chs_in_f[2][DATA][14] , \chs_in_f[2][DATA][13] , 
        \chs_in_f[2][DATA][12] , \chs_in_f[2][DATA][11] , 
        \chs_in_f[2][DATA][10] , \chs_in_f[2][DATA][9] , 
        \chs_in_f[2][DATA][8] , \chs_in_f[2][DATA][7] , \chs_in_f[2][DATA][6] , 
        \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] , \chs_in_f[2][DATA][3] , 
        \chs_in_f[2][DATA][2] , \chs_in_f[2][DATA][1] , \chs_in_f[2][DATA][0] }), .chan_out_b(\chs_in_b[2][ACK] ), .sel({\switch_sel[2][4] , 
        \switch_sel[2][3] , \switch_sel[2][2] , \switch_sel[2][1] , 
        \switch_sel[2][0] }) );
  hpu_0_1_0 east_hpu ( .preset(n2), .chan_in_f({\east_hpu_f[REQ] , 
        \east_hpu_f[DATA][34] , \east_hpu_f[DATA][33] , \east_hpu_f[DATA][32] , 
        \east_hpu_f[DATA][31] , \east_hpu_f[DATA][30] , \east_hpu_f[DATA][29] , 
        \east_hpu_f[DATA][28] , \east_hpu_f[DATA][27] , \east_hpu_f[DATA][26] , 
        \east_hpu_f[DATA][25] , \east_hpu_f[DATA][24] , \east_hpu_f[DATA][23] , 
        \east_hpu_f[DATA][22] , \east_hpu_f[DATA][21] , \east_hpu_f[DATA][20] , 
        \east_hpu_f[DATA][19] , \east_hpu_f[DATA][18] , \east_hpu_f[DATA][17] , 
        \east_hpu_f[DATA][16] , \east_hpu_f[DATA][15] , \east_hpu_f[DATA][14] , 
        \east_hpu_f[DATA][13] , \east_hpu_f[DATA][12] , \east_hpu_f[DATA][11] , 
        \east_hpu_f[DATA][10] , \east_hpu_f[DATA][9] , \east_hpu_f[DATA][8] , 
        \east_hpu_f[DATA][7] , \east_hpu_f[DATA][6] , \east_hpu_f[DATA][5] , 
        \east_hpu_f[DATA][4] , \east_hpu_f[DATA][3] , \east_hpu_f[DATA][2] , 
        \east_hpu_f[DATA][1] , \east_hpu_f[DATA][0] }), .chan_in_b(
        \east_hpu_b[ACK] ), .chan_out_f({\chs_in_f[1][REQ] , 
        \chs_in_f[1][DATA][34] , \chs_in_f[1][DATA][33] , 
        \chs_in_f[1][DATA][32] , \chs_in_f[1][DATA][31] , 
        \chs_in_f[1][DATA][30] , \chs_in_f[1][DATA][29] , 
        \chs_in_f[1][DATA][28] , \chs_in_f[1][DATA][27] , 
        \chs_in_f[1][DATA][26] , \chs_in_f[1][DATA][25] , 
        \chs_in_f[1][DATA][24] , \chs_in_f[1][DATA][23] , 
        \chs_in_f[1][DATA][22] , \chs_in_f[1][DATA][21] , 
        \chs_in_f[1][DATA][20] , \chs_in_f[1][DATA][19] , 
        \chs_in_f[1][DATA][18] , \chs_in_f[1][DATA][17] , 
        \chs_in_f[1][DATA][16] , \chs_in_f[1][DATA][15] , 
        \chs_in_f[1][DATA][14] , \chs_in_f[1][DATA][13] , 
        \chs_in_f[1][DATA][12] , \chs_in_f[1][DATA][11] , 
        \chs_in_f[1][DATA][10] , \chs_in_f[1][DATA][9] , 
        \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] , \chs_in_f[1][DATA][6] , 
        \chs_in_f[1][DATA][5] , \chs_in_f[1][DATA][4] , \chs_in_f[1][DATA][3] , 
        \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] , \chs_in_f[1][DATA][0] }), .chan_out_b(\chs_in_b[1][ACK] ), .sel({\switch_sel[1][4] , 
        \switch_sel[1][3] , \switch_sel[1][2] , \switch_sel[1][1] , 
        \switch_sel[1][0] }) );
  hpu_0_3_0 west_hpu ( .preset(n2), .chan_in_f({\west_hpu_f[REQ] , 
        \west_hpu_f[DATA][34] , \west_hpu_f[DATA][33] , \west_hpu_f[DATA][32] , 
        \west_hpu_f[DATA][31] , \west_hpu_f[DATA][30] , \west_hpu_f[DATA][29] , 
        \west_hpu_f[DATA][28] , \west_hpu_f[DATA][27] , \west_hpu_f[DATA][26] , 
        \west_hpu_f[DATA][25] , \west_hpu_f[DATA][24] , \west_hpu_f[DATA][23] , 
        \west_hpu_f[DATA][22] , \west_hpu_f[DATA][21] , \west_hpu_f[DATA][20] , 
        \west_hpu_f[DATA][19] , \west_hpu_f[DATA][18] , \west_hpu_f[DATA][17] , 
        \west_hpu_f[DATA][16] , \west_hpu_f[DATA][15] , \west_hpu_f[DATA][14] , 
        \west_hpu_f[DATA][13] , \west_hpu_f[DATA][12] , \west_hpu_f[DATA][11] , 
        \west_hpu_f[DATA][10] , \west_hpu_f[DATA][9] , \west_hpu_f[DATA][8] , 
        \west_hpu_f[DATA][7] , \west_hpu_f[DATA][6] , \west_hpu_f[DATA][5] , 
        \west_hpu_f[DATA][4] , \west_hpu_f[DATA][3] , \west_hpu_f[DATA][2] , 
        \west_hpu_f[DATA][1] , \west_hpu_f[DATA][0] }), .chan_in_b(
        \west_hpu_b[ACK] ), .chan_out_f({\chs_in_f[3][REQ] , 
        \chs_in_f[3][DATA][34] , \chs_in_f[3][DATA][33] , 
        \chs_in_f[3][DATA][32] , \chs_in_f[3][DATA][31] , 
        \chs_in_f[3][DATA][30] , \chs_in_f[3][DATA][29] , 
        \chs_in_f[3][DATA][28] , \chs_in_f[3][DATA][27] , 
        \chs_in_f[3][DATA][26] , \chs_in_f[3][DATA][25] , 
        \chs_in_f[3][DATA][24] , \chs_in_f[3][DATA][23] , 
        \chs_in_f[3][DATA][22] , \chs_in_f[3][DATA][21] , 
        \chs_in_f[3][DATA][20] , \chs_in_f[3][DATA][19] , 
        \chs_in_f[3][DATA][18] , \chs_in_f[3][DATA][17] , 
        \chs_in_f[3][DATA][16] , \chs_in_f[3][DATA][15] , 
        \chs_in_f[3][DATA][14] , \chs_in_f[3][DATA][13] , 
        \chs_in_f[3][DATA][12] , \chs_in_f[3][DATA][11] , 
        \chs_in_f[3][DATA][10] , \chs_in_f[3][DATA][9] , 
        \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] , \chs_in_f[3][DATA][6] , 
        \chs_in_f[3][DATA][5] , \chs_in_f[3][DATA][4] , \chs_in_f[3][DATA][3] , 
        \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] , \chs_in_f[3][DATA][0] }), .chan_out_b(\chs_in_b[3][ACK] ), .sel({\switch_sel[3][4] , 
        \switch_sel[3][3] , \switch_sel[3][2] , \switch_sel[3][1] , 
        \switch_sel[3][0] }) );
  hpu_1_x_0 resource_hpu ( .preset(n2), .chan_in_f({\resource_hpu_f[REQ] , 
        \resource_hpu_f[DATA][34] , \resource_hpu_f[DATA][33] , 
        \resource_hpu_f[DATA][32] , \resource_hpu_f[DATA][31] , 
        \resource_hpu_f[DATA][30] , \resource_hpu_f[DATA][29] , 
        \resource_hpu_f[DATA][28] , \resource_hpu_f[DATA][27] , 
        \resource_hpu_f[DATA][26] , \resource_hpu_f[DATA][25] , 
        \resource_hpu_f[DATA][24] , \resource_hpu_f[DATA][23] , 
        \resource_hpu_f[DATA][22] , \resource_hpu_f[DATA][21] , 
        \resource_hpu_f[DATA][20] , \resource_hpu_f[DATA][19] , 
        \resource_hpu_f[DATA][18] , \resource_hpu_f[DATA][17] , 
        \resource_hpu_f[DATA][16] , \resource_hpu_f[DATA][15] , 
        \resource_hpu_f[DATA][14] , \resource_hpu_f[DATA][13] , 
        \resource_hpu_f[DATA][12] , \resource_hpu_f[DATA][11] , 
        \resource_hpu_f[DATA][10] , \resource_hpu_f[DATA][9] , 
        \resource_hpu_f[DATA][8] , \resource_hpu_f[DATA][7] , 
        \resource_hpu_f[DATA][6] , \resource_hpu_f[DATA][5] , 
        \resource_hpu_f[DATA][4] , \resource_hpu_f[DATA][3] , 
        \resource_hpu_f[DATA][2] , \resource_hpu_f[DATA][1] , 
        \resource_hpu_f[DATA][0] }), .chan_in_b(\resource_hpu_b[ACK] ), 
        .chan_out_f({\chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] , 
        \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] , 
        \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] , 
        \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] , 
        \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] , 
        \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] , 
        \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] , 
        \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] , 
        \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] , 
        \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] , 
        \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] , 
        \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] , 
        \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] , 
        \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] , \chs_in_f[4][DATA][7] , 
        \chs_in_f[4][DATA][6] , \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] , 
        \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] , \chs_in_f[4][DATA][1] , 
        \chs_in_f[4][DATA][0] }), .chan_out_b(\chs_in_b[4][ACK] ), .sel({
        \switch_sel[4][4] , \switch_sel[4][3] , \switch_sel[4][2] , 
        \switch_sel[4][1] , \switch_sel[4][0] }) );
  crossbar_stage_0 xbar_with_latches ( .preset(n3), .switch_sel({1'b0, 
        \switch_sel[4][3] , \switch_sel[4][2] , \switch_sel[4][1] , 
        \switch_sel[4][0] , \switch_sel[3][4] , 1'b0, \switch_sel[3][2] , 
        \switch_sel[3][1] , \switch_sel[3][0] , \switch_sel[2][4] , 
        \switch_sel[2][3] , 1'b0, \switch_sel[2][1] , \switch_sel[2][0] , 
        \switch_sel[1][4] , \switch_sel[1][3] , \switch_sel[1][2] , 1'b0, 
        \switch_sel[1][0] , \switch_sel[0][4] , \switch_sel[0][3] , 
        \switch_sel[0][2] , \switch_sel[0][1] , 1'b0}), .chs_in_f({
        \chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] , \chs_in_f[4][DATA][33] , 
        \chs_in_f[4][DATA][32] , \chs_in_f[4][DATA][31] , 
        \chs_in_f[4][DATA][30] , \chs_in_f[4][DATA][29] , 
        \chs_in_f[4][DATA][28] , \chs_in_f[4][DATA][27] , 
        \chs_in_f[4][DATA][26] , \chs_in_f[4][DATA][25] , 
        \chs_in_f[4][DATA][24] , \chs_in_f[4][DATA][23] , 
        \chs_in_f[4][DATA][22] , \chs_in_f[4][DATA][21] , 
        \chs_in_f[4][DATA][20] , \chs_in_f[4][DATA][19] , 
        \chs_in_f[4][DATA][18] , \chs_in_f[4][DATA][17] , 
        \chs_in_f[4][DATA][16] , \chs_in_f[4][DATA][15] , 
        \chs_in_f[4][DATA][14] , \chs_in_f[4][DATA][13] , 
        \chs_in_f[4][DATA][12] , \chs_in_f[4][DATA][11] , 
        \chs_in_f[4][DATA][10] , \chs_in_f[4][DATA][9] , 
        \chs_in_f[4][DATA][8] , \chs_in_f[4][DATA][7] , \chs_in_f[4][DATA][6] , 
        \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] , \chs_in_f[4][DATA][3] , 
        \chs_in_f[4][DATA][2] , \chs_in_f[4][DATA][1] , \chs_in_f[4][DATA][0] , 
        \chs_in_f[3][REQ] , \chs_in_f[3][DATA][34] , \chs_in_f[3][DATA][33] , 
        \chs_in_f[3][DATA][32] , \chs_in_f[3][DATA][31] , 
        \chs_in_f[3][DATA][30] , \chs_in_f[3][DATA][29] , 
        \chs_in_f[3][DATA][28] , \chs_in_f[3][DATA][27] , 
        \chs_in_f[3][DATA][26] , \chs_in_f[3][DATA][25] , 
        \chs_in_f[3][DATA][24] , \chs_in_f[3][DATA][23] , 
        \chs_in_f[3][DATA][22] , \chs_in_f[3][DATA][21] , 
        \chs_in_f[3][DATA][20] , \chs_in_f[3][DATA][19] , 
        \chs_in_f[3][DATA][18] , \chs_in_f[3][DATA][17] , 
        \chs_in_f[3][DATA][16] , \chs_in_f[3][DATA][15] , 
        \chs_in_f[3][DATA][14] , \chs_in_f[3][DATA][13] , 
        \chs_in_f[3][DATA][12] , \chs_in_f[3][DATA][11] , 
        \chs_in_f[3][DATA][10] , \chs_in_f[3][DATA][9] , 
        \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] , \chs_in_f[3][DATA][6] , 
        \chs_in_f[3][DATA][5] , \chs_in_f[3][DATA][4] , \chs_in_f[3][DATA][3] , 
        \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] , \chs_in_f[3][DATA][0] , 
        \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] , \chs_in_f[2][DATA][33] , 
        \chs_in_f[2][DATA][32] , \chs_in_f[2][DATA][31] , 
        \chs_in_f[2][DATA][30] , \chs_in_f[2][DATA][29] , 
        \chs_in_f[2][DATA][28] , \chs_in_f[2][DATA][27] , 
        \chs_in_f[2][DATA][26] , \chs_in_f[2][DATA][25] , 
        \chs_in_f[2][DATA][24] , \chs_in_f[2][DATA][23] , 
        \chs_in_f[2][DATA][22] , \chs_in_f[2][DATA][21] , 
        \chs_in_f[2][DATA][20] , \chs_in_f[2][DATA][19] , 
        \chs_in_f[2][DATA][18] , \chs_in_f[2][DATA][17] , 
        \chs_in_f[2][DATA][16] , \chs_in_f[2][DATA][15] , 
        \chs_in_f[2][DATA][14] , \chs_in_f[2][DATA][13] , 
        \chs_in_f[2][DATA][12] , \chs_in_f[2][DATA][11] , 
        \chs_in_f[2][DATA][10] , \chs_in_f[2][DATA][9] , 
        \chs_in_f[2][DATA][8] , \chs_in_f[2][DATA][7] , \chs_in_f[2][DATA][6] , 
        \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] , \chs_in_f[2][DATA][3] , 
        \chs_in_f[2][DATA][2] , \chs_in_f[2][DATA][1] , \chs_in_f[2][DATA][0] , 
        \chs_in_f[1][REQ] , \chs_in_f[1][DATA][34] , \chs_in_f[1][DATA][33] , 
        \chs_in_f[1][DATA][32] , \chs_in_f[1][DATA][31] , 
        \chs_in_f[1][DATA][30] , \chs_in_f[1][DATA][29] , 
        \chs_in_f[1][DATA][28] , \chs_in_f[1][DATA][27] , 
        \chs_in_f[1][DATA][26] , \chs_in_f[1][DATA][25] , 
        \chs_in_f[1][DATA][24] , \chs_in_f[1][DATA][23] , 
        \chs_in_f[1][DATA][22] , \chs_in_f[1][DATA][21] , 
        \chs_in_f[1][DATA][20] , \chs_in_f[1][DATA][19] , 
        \chs_in_f[1][DATA][18] , \chs_in_f[1][DATA][17] , 
        \chs_in_f[1][DATA][16] , \chs_in_f[1][DATA][15] , 
        \chs_in_f[1][DATA][14] , \chs_in_f[1][DATA][13] , 
        \chs_in_f[1][DATA][12] , \chs_in_f[1][DATA][11] , 
        \chs_in_f[1][DATA][10] , \chs_in_f[1][DATA][9] , 
        \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] , \chs_in_f[1][DATA][6] , 
        \chs_in_f[1][DATA][5] , \chs_in_f[1][DATA][4] , \chs_in_f[1][DATA][3] , 
        \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] , \chs_in_f[1][DATA][0] , 
        \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] , \chs_in_f[0][DATA][33] , 
        \chs_in_f[0][DATA][32] , \chs_in_f[0][DATA][31] , 
        \chs_in_f[0][DATA][30] , \chs_in_f[0][DATA][29] , 
        \chs_in_f[0][DATA][28] , \chs_in_f[0][DATA][27] , 
        \chs_in_f[0][DATA][26] , \chs_in_f[0][DATA][25] , 
        \chs_in_f[0][DATA][24] , \chs_in_f[0][DATA][23] , 
        \chs_in_f[0][DATA][22] , \chs_in_f[0][DATA][21] , 
        \chs_in_f[0][DATA][20] , \chs_in_f[0][DATA][19] , 
        \chs_in_f[0][DATA][18] , \chs_in_f[0][DATA][17] , 
        \chs_in_f[0][DATA][16] , \chs_in_f[0][DATA][15] , 
        \chs_in_f[0][DATA][14] , \chs_in_f[0][DATA][13] , 
        \chs_in_f[0][DATA][12] , \chs_in_f[0][DATA][11] , 
        \chs_in_f[0][DATA][10] , \chs_in_f[0][DATA][9] , 
        \chs_in_f[0][DATA][8] , \chs_in_f[0][DATA][7] , \chs_in_f[0][DATA][6] , 
        \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] , \chs_in_f[0][DATA][3] , 
        \chs_in_f[0][DATA][2] , \chs_in_f[0][DATA][1] , \chs_in_f[0][DATA][0] }), .chs_in_b({\chs_in_b[4][ACK] , \chs_in_b[3][ACK] , \chs_in_b[2][ACK] , 
        \chs_in_b[1][ACK] , \chs_in_b[0][ACK] }), .latches_out_f({
        \resource_out_f[REQ] , \resource_out_f[DATA][34] , 
        \resource_out_f[DATA][33] , \resource_out_f[DATA][32] , 
        \resource_out_f[DATA][31] , \resource_out_f[DATA][30] , 
        \resource_out_f[DATA][29] , \resource_out_f[DATA][28] , 
        \resource_out_f[DATA][27] , \resource_out_f[DATA][26] , 
        \resource_out_f[DATA][25] , \resource_out_f[DATA][24] , 
        \resource_out_f[DATA][23] , \resource_out_f[DATA][22] , 
        \resource_out_f[DATA][21] , \resource_out_f[DATA][20] , 
        \resource_out_f[DATA][19] , \resource_out_f[DATA][18] , 
        \resource_out_f[DATA][17] , \resource_out_f[DATA][16] , 
        \resource_out_f[DATA][15] , \resource_out_f[DATA][14] , 
        \resource_out_f[DATA][13] , \resource_out_f[DATA][12] , 
        \resource_out_f[DATA][11] , \resource_out_f[DATA][10] , 
        \resource_out_f[DATA][9] , \resource_out_f[DATA][8] , 
        \resource_out_f[DATA][7] , \resource_out_f[DATA][6] , 
        \resource_out_f[DATA][5] , \resource_out_f[DATA][4] , 
        \resource_out_f[DATA][3] , \resource_out_f[DATA][2] , 
        \resource_out_f[DATA][1] , \resource_out_f[DATA][0] , 
        \west_out_f[REQ] , \west_out_f[DATA][34] , \west_out_f[DATA][33] , 
        \west_out_f[DATA][32] , \west_out_f[DATA][31] , \west_out_f[DATA][30] , 
        \west_out_f[DATA][29] , \west_out_f[DATA][28] , \west_out_f[DATA][27] , 
        \west_out_f[DATA][26] , \west_out_f[DATA][25] , \west_out_f[DATA][24] , 
        \west_out_f[DATA][23] , \west_out_f[DATA][22] , \west_out_f[DATA][21] , 
        \west_out_f[DATA][20] , \west_out_f[DATA][19] , \west_out_f[DATA][18] , 
        \west_out_f[DATA][17] , \west_out_f[DATA][16] , \west_out_f[DATA][15] , 
        \west_out_f[DATA][14] , \west_out_f[DATA][13] , \west_out_f[DATA][12] , 
        \west_out_f[DATA][11] , \west_out_f[DATA][10] , \west_out_f[DATA][9] , 
        \west_out_f[DATA][8] , \west_out_f[DATA][7] , \west_out_f[DATA][6] , 
        \west_out_f[DATA][5] , \west_out_f[DATA][4] , \west_out_f[DATA][3] , 
        \west_out_f[DATA][2] , \west_out_f[DATA][1] , \west_out_f[DATA][0] , 
        \south_out_f[REQ] , \south_out_f[DATA][34] , \south_out_f[DATA][33] , 
        \south_out_f[DATA][32] , \south_out_f[DATA][31] , 
        \south_out_f[DATA][30] , \south_out_f[DATA][29] , 
        \south_out_f[DATA][28] , \south_out_f[DATA][27] , 
        \south_out_f[DATA][26] , \south_out_f[DATA][25] , 
        \south_out_f[DATA][24] , \south_out_f[DATA][23] , 
        \south_out_f[DATA][22] , \south_out_f[DATA][21] , 
        \south_out_f[DATA][20] , \south_out_f[DATA][19] , 
        \south_out_f[DATA][18] , \south_out_f[DATA][17] , 
        \south_out_f[DATA][16] , \south_out_f[DATA][15] , 
        \south_out_f[DATA][14] , \south_out_f[DATA][13] , 
        \south_out_f[DATA][12] , \south_out_f[DATA][11] , 
        \south_out_f[DATA][10] , \south_out_f[DATA][9] , 
        \south_out_f[DATA][8] , \south_out_f[DATA][7] , \south_out_f[DATA][6] , 
        \south_out_f[DATA][5] , \south_out_f[DATA][4] , \south_out_f[DATA][3] , 
        \south_out_f[DATA][2] , \south_out_f[DATA][1] , \south_out_f[DATA][0] , 
        \east_out_f[REQ] , \east_out_f[DATA][34] , \east_out_f[DATA][33] , 
        \east_out_f[DATA][32] , \east_out_f[DATA][31] , \east_out_f[DATA][30] , 
        \east_out_f[DATA][29] , \east_out_f[DATA][28] , \east_out_f[DATA][27] , 
        \east_out_f[DATA][26] , \east_out_f[DATA][25] , \east_out_f[DATA][24] , 
        \east_out_f[DATA][23] , \east_out_f[DATA][22] , \east_out_f[DATA][21] , 
        \east_out_f[DATA][20] , \east_out_f[DATA][19] , \east_out_f[DATA][18] , 
        \east_out_f[DATA][17] , \east_out_f[DATA][16] , \east_out_f[DATA][15] , 
        \east_out_f[DATA][14] , \east_out_f[DATA][13] , \east_out_f[DATA][12] , 
        \east_out_f[DATA][11] , \east_out_f[DATA][10] , \east_out_f[DATA][9] , 
        \east_out_f[DATA][8] , \east_out_f[DATA][7] , \east_out_f[DATA][6] , 
        \east_out_f[DATA][5] , \east_out_f[DATA][4] , \east_out_f[DATA][3] , 
        \east_out_f[DATA][2] , \east_out_f[DATA][1] , \east_out_f[DATA][0] , 
        \north_out_f[REQ] , \north_out_f[DATA][34] , \north_out_f[DATA][33] , 
        \north_out_f[DATA][32] , \north_out_f[DATA][31] , 
        \north_out_f[DATA][30] , \north_out_f[DATA][29] , 
        \north_out_f[DATA][28] , \north_out_f[DATA][27] , 
        \north_out_f[DATA][26] , \north_out_f[DATA][25] , 
        \north_out_f[DATA][24] , \north_out_f[DATA][23] , 
        \north_out_f[DATA][22] , \north_out_f[DATA][21] , 
        \north_out_f[DATA][20] , \north_out_f[DATA][19] , 
        \north_out_f[DATA][18] , \north_out_f[DATA][17] , 
        \north_out_f[DATA][16] , \north_out_f[DATA][15] , 
        \north_out_f[DATA][14] , \north_out_f[DATA][13] , 
        \north_out_f[DATA][12] , \north_out_f[DATA][11] , 
        \north_out_f[DATA][10] , \north_out_f[DATA][9] , 
        \north_out_f[DATA][8] , \north_out_f[DATA][7] , \north_out_f[DATA][6] , 
        \north_out_f[DATA][5] , \north_out_f[DATA][4] , \north_out_f[DATA][3] , 
        \north_out_f[DATA][2] , \north_out_f[DATA][1] , \north_out_f[DATA][0] }), .latches_out_b({\resource_out_b[ACK] , \west_out_b[ACK] , 
        \south_out_b[ACK] , \east_out_b[ACK] , \north_out_b[ACK] }) );
  HS65_LS_BFX9 U1 ( .A(preset), .Z(n3) );
  HS65_LS_BFX9 U2 ( .A(preset), .Z(n2) );
endmodule


module noc_node_0 ( p_clk, n_clk, reset, .proc_in({\proc_in[MCMD][1] , 
        \proc_in[MCMD][0] , \proc_in[MADDR][31] , \proc_in[MADDR][30] , 
        \proc_in[MADDR][29] , \proc_in[MADDR][28] , \proc_in[MADDR][27] , 
        \proc_in[MADDR][26] , \proc_in[MADDR][25] , \proc_in[MADDR][24] , 
        \proc_in[MADDR][23] , \proc_in[MADDR][22] , \proc_in[MADDR][21] , 
        \proc_in[MADDR][20] , \proc_in[MADDR][19] , \proc_in[MADDR][18] , 
        \proc_in[MADDR][17] , \proc_in[MADDR][16] , \proc_in[MADDR][15] , 
        \proc_in[MADDR][14] , \proc_in[MADDR][13] , \proc_in[MADDR][12] , 
        \proc_in[MADDR][11] , \proc_in[MADDR][10] , \proc_in[MADDR][9] , 
        \proc_in[MADDR][8] , \proc_in[MADDR][7] , \proc_in[MADDR][6] , 
        \proc_in[MADDR][5] , \proc_in[MADDR][4] , \proc_in[MADDR][3] , 
        \proc_in[MADDR][2] , \proc_in[MADDR][1] , \proc_in[MADDR][0] , 
        \proc_in[MDATA][31] , \proc_in[MDATA][30] , \proc_in[MDATA][29] , 
        \proc_in[MDATA][28] , \proc_in[MDATA][27] , \proc_in[MDATA][26] , 
        \proc_in[MDATA][25] , \proc_in[MDATA][24] , \proc_in[MDATA][23] , 
        \proc_in[MDATA][22] , \proc_in[MDATA][21] , \proc_in[MDATA][20] , 
        \proc_in[MDATA][19] , \proc_in[MDATA][18] , \proc_in[MDATA][17] , 
        \proc_in[MDATA][16] , \proc_in[MDATA][15] , \proc_in[MDATA][14] , 
        \proc_in[MDATA][13] , \proc_in[MDATA][12] , \proc_in[MDATA][11] , 
        \proc_in[MDATA][10] , \proc_in[MDATA][9] , \proc_in[MDATA][8] , 
        \proc_in[MDATA][7] , \proc_in[MDATA][6] , \proc_in[MDATA][5] , 
        \proc_in[MDATA][4] , \proc_in[MDATA][3] , \proc_in[MDATA][2] , 
        \proc_in[MDATA][1] , \proc_in[MDATA][0] }), .proc_out({
        \proc_out[SCMDACCEPT] , \proc_out[SRESP] , \proc_out[SDATA][31] , 
        \proc_out[SDATA][30] , \proc_out[SDATA][29] , \proc_out[SDATA][28] , 
        \proc_out[SDATA][27] , \proc_out[SDATA][26] , \proc_out[SDATA][25] , 
        \proc_out[SDATA][24] , \proc_out[SDATA][23] , \proc_out[SDATA][22] , 
        \proc_out[SDATA][21] , \proc_out[SDATA][20] , \proc_out[SDATA][19] , 
        \proc_out[SDATA][18] , \proc_out[SDATA][17] , \proc_out[SDATA][16] , 
        \proc_out[SDATA][15] , \proc_out[SDATA][14] , \proc_out[SDATA][13] , 
        \proc_out[SDATA][12] , \proc_out[SDATA][11] , \proc_out[SDATA][10] , 
        \proc_out[SDATA][9] , \proc_out[SDATA][8] , \proc_out[SDATA][7] , 
        \proc_out[SDATA][6] , \proc_out[SDATA][5] , \proc_out[SDATA][4] , 
        \proc_out[SDATA][3] , \proc_out[SDATA][2] , \proc_out[SDATA][1] , 
        \proc_out[SDATA][0] }), .spm_in({\spm_in[SCMDACCEPT] , \spm_in[SRESP] , 
        \spm_in[SDATA][63] , \spm_in[SDATA][62] , \spm_in[SDATA][61] , 
        \spm_in[SDATA][60] , \spm_in[SDATA][59] , \spm_in[SDATA][58] , 
        \spm_in[SDATA][57] , \spm_in[SDATA][56] , \spm_in[SDATA][55] , 
        \spm_in[SDATA][54] , \spm_in[SDATA][53] , \spm_in[SDATA][52] , 
        \spm_in[SDATA][51] , \spm_in[SDATA][50] , \spm_in[SDATA][49] , 
        \spm_in[SDATA][48] , \spm_in[SDATA][47] , \spm_in[SDATA][46] , 
        \spm_in[SDATA][45] , \spm_in[SDATA][44] , \spm_in[SDATA][43] , 
        \spm_in[SDATA][42] , \spm_in[SDATA][41] , \spm_in[SDATA][40] , 
        \spm_in[SDATA][39] , \spm_in[SDATA][38] , \spm_in[SDATA][37] , 
        \spm_in[SDATA][36] , \spm_in[SDATA][35] , \spm_in[SDATA][34] , 
        \spm_in[SDATA][33] , \spm_in[SDATA][32] , \spm_in[SDATA][31] , 
        \spm_in[SDATA][30] , \spm_in[SDATA][29] , \spm_in[SDATA][28] , 
        \spm_in[SDATA][27] , \spm_in[SDATA][26] , \spm_in[SDATA][25] , 
        \spm_in[SDATA][24] , \spm_in[SDATA][23] , \spm_in[SDATA][22] , 
        \spm_in[SDATA][21] , \spm_in[SDATA][20] , \spm_in[SDATA][19] , 
        \spm_in[SDATA][18] , \spm_in[SDATA][17] , \spm_in[SDATA][16] , 
        \spm_in[SDATA][15] , \spm_in[SDATA][14] , \spm_in[SDATA][13] , 
        \spm_in[SDATA][12] , \spm_in[SDATA][11] , \spm_in[SDATA][10] , 
        \spm_in[SDATA][9] , \spm_in[SDATA][8] , \spm_in[SDATA][7] , 
        \spm_in[SDATA][6] , \spm_in[SDATA][5] , \spm_in[SDATA][4] , 
        \spm_in[SDATA][3] , \spm_in[SDATA][2] , \spm_in[SDATA][1] , 
        \spm_in[SDATA][0] }), .spm_out({\spm_out[MCMD][1] , \spm_out[MCMD][0] , 
        \spm_out[MADDR][31] , \spm_out[MADDR][30] , \spm_out[MADDR][29] , 
        \spm_out[MADDR][28] , \spm_out[MADDR][27] , \spm_out[MADDR][26] , 
        \spm_out[MADDR][25] , \spm_out[MADDR][24] , \spm_out[MADDR][23] , 
        \spm_out[MADDR][22] , \spm_out[MADDR][21] , \spm_out[MADDR][20] , 
        \spm_out[MADDR][19] , \spm_out[MADDR][18] , \spm_out[MADDR][17] , 
        \spm_out[MADDR][16] , \spm_out[MADDR][15] , \spm_out[MADDR][14] , 
        \spm_out[MADDR][13] , \spm_out[MADDR][12] , \spm_out[MADDR][11] , 
        \spm_out[MADDR][10] , \spm_out[MADDR][9] , \spm_out[MADDR][8] , 
        \spm_out[MADDR][7] , \spm_out[MADDR][6] , \spm_out[MADDR][5] , 
        \spm_out[MADDR][4] , \spm_out[MADDR][3] , \spm_out[MADDR][2] , 
        \spm_out[MADDR][1] , \spm_out[MADDR][0] , \spm_out[MDATA][63] , 
        \spm_out[MDATA][62] , \spm_out[MDATA][61] , \spm_out[MDATA][60] , 
        \spm_out[MDATA][59] , \spm_out[MDATA][58] , \spm_out[MDATA][57] , 
        \spm_out[MDATA][56] , \spm_out[MDATA][55] , \spm_out[MDATA][54] , 
        \spm_out[MDATA][53] , \spm_out[MDATA][52] , \spm_out[MDATA][51] , 
        \spm_out[MDATA][50] , \spm_out[MDATA][49] , \spm_out[MDATA][48] , 
        \spm_out[MDATA][47] , \spm_out[MDATA][46] , \spm_out[MDATA][45] , 
        \spm_out[MDATA][44] , \spm_out[MDATA][43] , \spm_out[MDATA][42] , 
        \spm_out[MDATA][41] , \spm_out[MDATA][40] , \spm_out[MDATA][39] , 
        \spm_out[MDATA][38] , \spm_out[MDATA][37] , \spm_out[MDATA][36] , 
        \spm_out[MDATA][35] , \spm_out[MDATA][34] , \spm_out[MDATA][33] , 
        \spm_out[MDATA][32] , \spm_out[MDATA][31] , \spm_out[MDATA][30] , 
        \spm_out[MDATA][29] , \spm_out[MDATA][28] , \spm_out[MDATA][27] , 
        \spm_out[MDATA][26] , \spm_out[MDATA][25] , \spm_out[MDATA][24] , 
        \spm_out[MDATA][23] , \spm_out[MDATA][22] , \spm_out[MDATA][21] , 
        \spm_out[MDATA][20] , \spm_out[MDATA][19] , \spm_out[MDATA][18] , 
        \spm_out[MDATA][17] , \spm_out[MDATA][16] , \spm_out[MDATA][15] , 
        \spm_out[MDATA][14] , \spm_out[MDATA][13] , \spm_out[MDATA][12] , 
        \spm_out[MDATA][11] , \spm_out[MDATA][10] , \spm_out[MDATA][9] , 
        \spm_out[MDATA][8] , \spm_out[MDATA][7] , \spm_out[MDATA][6] , 
        \spm_out[MDATA][5] , \spm_out[MDATA][4] , \spm_out[MDATA][3] , 
        \spm_out[MDATA][2] , \spm_out[MDATA][1] , \spm_out[MDATA][0] }), 
    .north_in_f({\north_in_f[REQ] , \north_in_f[DATA][34] , 
        \north_in_f[DATA][33] , \north_in_f[DATA][32] , \north_in_f[DATA][31] , 
        \north_in_f[DATA][30] , \north_in_f[DATA][29] , \north_in_f[DATA][28] , 
        \north_in_f[DATA][27] , \north_in_f[DATA][26] , \north_in_f[DATA][25] , 
        \north_in_f[DATA][24] , \north_in_f[DATA][23] , \north_in_f[DATA][22] , 
        \north_in_f[DATA][21] , \north_in_f[DATA][20] , \north_in_f[DATA][19] , 
        \north_in_f[DATA][18] , \north_in_f[DATA][17] , \north_in_f[DATA][16] , 
        \north_in_f[DATA][15] , \north_in_f[DATA][14] , \north_in_f[DATA][13] , 
        \north_in_f[DATA][12] , \north_in_f[DATA][11] , \north_in_f[DATA][10] , 
        \north_in_f[DATA][9] , \north_in_f[DATA][8] , \north_in_f[DATA][7] , 
        \north_in_f[DATA][6] , \north_in_f[DATA][5] , \north_in_f[DATA][4] , 
        \north_in_f[DATA][3] , \north_in_f[DATA][2] , \north_in_f[DATA][1] , 
        \north_in_f[DATA][0] }), .north_in_b(\north_in_b[ACK] ), .east_in_f({
        \east_in_f[REQ] , \east_in_f[DATA][34] , \east_in_f[DATA][33] , 
        \east_in_f[DATA][32] , \east_in_f[DATA][31] , \east_in_f[DATA][30] , 
        \east_in_f[DATA][29] , \east_in_f[DATA][28] , \east_in_f[DATA][27] , 
        \east_in_f[DATA][26] , \east_in_f[DATA][25] , \east_in_f[DATA][24] , 
        \east_in_f[DATA][23] , \east_in_f[DATA][22] , \east_in_f[DATA][21] , 
        \east_in_f[DATA][20] , \east_in_f[DATA][19] , \east_in_f[DATA][18] , 
        \east_in_f[DATA][17] , \east_in_f[DATA][16] , \east_in_f[DATA][15] , 
        \east_in_f[DATA][14] , \east_in_f[DATA][13] , \east_in_f[DATA][12] , 
        \east_in_f[DATA][11] , \east_in_f[DATA][10] , \east_in_f[DATA][9] , 
        \east_in_f[DATA][8] , \east_in_f[DATA][7] , \east_in_f[DATA][6] , 
        \east_in_f[DATA][5] , \east_in_f[DATA][4] , \east_in_f[DATA][3] , 
        \east_in_f[DATA][2] , \east_in_f[DATA][1] , \east_in_f[DATA][0] }), 
    .east_in_b(\east_in_b[ACK] ), .south_in_f({\south_in_f[REQ] , 
        \south_in_f[DATA][34] , \south_in_f[DATA][33] , \south_in_f[DATA][32] , 
        \south_in_f[DATA][31] , \south_in_f[DATA][30] , \south_in_f[DATA][29] , 
        \south_in_f[DATA][28] , \south_in_f[DATA][27] , \south_in_f[DATA][26] , 
        \south_in_f[DATA][25] , \south_in_f[DATA][24] , \south_in_f[DATA][23] , 
        \south_in_f[DATA][22] , \south_in_f[DATA][21] , \south_in_f[DATA][20] , 
        \south_in_f[DATA][19] , \south_in_f[DATA][18] , \south_in_f[DATA][17] , 
        \south_in_f[DATA][16] , \south_in_f[DATA][15] , \south_in_f[DATA][14] , 
        \south_in_f[DATA][13] , \south_in_f[DATA][12] , \south_in_f[DATA][11] , 
        \south_in_f[DATA][10] , \south_in_f[DATA][9] , \south_in_f[DATA][8] , 
        \south_in_f[DATA][7] , \south_in_f[DATA][6] , \south_in_f[DATA][5] , 
        \south_in_f[DATA][4] , \south_in_f[DATA][3] , \south_in_f[DATA][2] , 
        \south_in_f[DATA][1] , \south_in_f[DATA][0] }), .south_in_b(
        \south_in_b[ACK] ), .west_in_f({\west_in_f[REQ] , 
        \west_in_f[DATA][34] , \west_in_f[DATA][33] , \west_in_f[DATA][32] , 
        \west_in_f[DATA][31] , \west_in_f[DATA][30] , \west_in_f[DATA][29] , 
        \west_in_f[DATA][28] , \west_in_f[DATA][27] , \west_in_f[DATA][26] , 
        \west_in_f[DATA][25] , \west_in_f[DATA][24] , \west_in_f[DATA][23] , 
        \west_in_f[DATA][22] , \west_in_f[DATA][21] , \west_in_f[DATA][20] , 
        \west_in_f[DATA][19] , \west_in_f[DATA][18] , \west_in_f[DATA][17] , 
        \west_in_f[DATA][16] , \west_in_f[DATA][15] , \west_in_f[DATA][14] , 
        \west_in_f[DATA][13] , \west_in_f[DATA][12] , \west_in_f[DATA][11] , 
        \west_in_f[DATA][10] , \west_in_f[DATA][9] , \west_in_f[DATA][8] , 
        \west_in_f[DATA][7] , \west_in_f[DATA][6] , \west_in_f[DATA][5] , 
        \west_in_f[DATA][4] , \west_in_f[DATA][3] , \west_in_f[DATA][2] , 
        \west_in_f[DATA][1] , \west_in_f[DATA][0] }), .west_in_b(
        \west_in_b[ACK] ), .north_out_f({\north_out_f[REQ] , 
        \north_out_f[DATA][34] , \north_out_f[DATA][33] , 
        \north_out_f[DATA][32] , \north_out_f[DATA][31] , 
        \north_out_f[DATA][30] , \north_out_f[DATA][29] , 
        \north_out_f[DATA][28] , \north_out_f[DATA][27] , 
        \north_out_f[DATA][26] , \north_out_f[DATA][25] , 
        \north_out_f[DATA][24] , \north_out_f[DATA][23] , 
        \north_out_f[DATA][22] , \north_out_f[DATA][21] , 
        \north_out_f[DATA][20] , \north_out_f[DATA][19] , 
        \north_out_f[DATA][18] , \north_out_f[DATA][17] , 
        \north_out_f[DATA][16] , \north_out_f[DATA][15] , 
        \north_out_f[DATA][14] , \north_out_f[DATA][13] , 
        \north_out_f[DATA][12] , \north_out_f[DATA][11] , 
        \north_out_f[DATA][10] , \north_out_f[DATA][9] , 
        \north_out_f[DATA][8] , \north_out_f[DATA][7] , \north_out_f[DATA][6] , 
        \north_out_f[DATA][5] , \north_out_f[DATA][4] , \north_out_f[DATA][3] , 
        \north_out_f[DATA][2] , \north_out_f[DATA][1] , \north_out_f[DATA][0] 
        }), .north_out_b(\north_out_b[ACK] ), .east_out_f({\east_out_f[REQ] , 
        \east_out_f[DATA][34] , \east_out_f[DATA][33] , \east_out_f[DATA][32] , 
        \east_out_f[DATA][31] , \east_out_f[DATA][30] , \east_out_f[DATA][29] , 
        \east_out_f[DATA][28] , \east_out_f[DATA][27] , \east_out_f[DATA][26] , 
        \east_out_f[DATA][25] , \east_out_f[DATA][24] , \east_out_f[DATA][23] , 
        \east_out_f[DATA][22] , \east_out_f[DATA][21] , \east_out_f[DATA][20] , 
        \east_out_f[DATA][19] , \east_out_f[DATA][18] , \east_out_f[DATA][17] , 
        \east_out_f[DATA][16] , \east_out_f[DATA][15] , \east_out_f[DATA][14] , 
        \east_out_f[DATA][13] , \east_out_f[DATA][12] , \east_out_f[DATA][11] , 
        \east_out_f[DATA][10] , \east_out_f[DATA][9] , \east_out_f[DATA][8] , 
        \east_out_f[DATA][7] , \east_out_f[DATA][6] , \east_out_f[DATA][5] , 
        \east_out_f[DATA][4] , \east_out_f[DATA][3] , \east_out_f[DATA][2] , 
        \east_out_f[DATA][1] , \east_out_f[DATA][0] }), .east_out_b(
        \east_out_b[ACK] ), .south_out_f({\south_out_f[REQ] , 
        \south_out_f[DATA][34] , \south_out_f[DATA][33] , 
        \south_out_f[DATA][32] , \south_out_f[DATA][31] , 
        \south_out_f[DATA][30] , \south_out_f[DATA][29] , 
        \south_out_f[DATA][28] , \south_out_f[DATA][27] , 
        \south_out_f[DATA][26] , \south_out_f[DATA][25] , 
        \south_out_f[DATA][24] , \south_out_f[DATA][23] , 
        \south_out_f[DATA][22] , \south_out_f[DATA][21] , 
        \south_out_f[DATA][20] , \south_out_f[DATA][19] , 
        \south_out_f[DATA][18] , \south_out_f[DATA][17] , 
        \south_out_f[DATA][16] , \south_out_f[DATA][15] , 
        \south_out_f[DATA][14] , \south_out_f[DATA][13] , 
        \south_out_f[DATA][12] , \south_out_f[DATA][11] , 
        \south_out_f[DATA][10] , \south_out_f[DATA][9] , 
        \south_out_f[DATA][8] , \south_out_f[DATA][7] , \south_out_f[DATA][6] , 
        \south_out_f[DATA][5] , \south_out_f[DATA][4] , \south_out_f[DATA][3] , 
        \south_out_f[DATA][2] , \south_out_f[DATA][1] , \south_out_f[DATA][0] 
        }), .south_out_b(\south_out_b[ACK] ), .west_out_f({\west_out_f[REQ] , 
        \west_out_f[DATA][34] , \west_out_f[DATA][33] , \west_out_f[DATA][32] , 
        \west_out_f[DATA][31] , \west_out_f[DATA][30] , \west_out_f[DATA][29] , 
        \west_out_f[DATA][28] , \west_out_f[DATA][27] , \west_out_f[DATA][26] , 
        \west_out_f[DATA][25] , \west_out_f[DATA][24] , \west_out_f[DATA][23] , 
        \west_out_f[DATA][22] , \west_out_f[DATA][21] , \west_out_f[DATA][20] , 
        \west_out_f[DATA][19] , \west_out_f[DATA][18] , \west_out_f[DATA][17] , 
        \west_out_f[DATA][16] , \west_out_f[DATA][15] , \west_out_f[DATA][14] , 
        \west_out_f[DATA][13] , \west_out_f[DATA][12] , \west_out_f[DATA][11] , 
        \west_out_f[DATA][10] , \west_out_f[DATA][9] , \west_out_f[DATA][8] , 
        \west_out_f[DATA][7] , \west_out_f[DATA][6] , \west_out_f[DATA][5] , 
        \west_out_f[DATA][4] , \west_out_f[DATA][3] , \west_out_f[DATA][2] , 
        \west_out_f[DATA][1] , \west_out_f[DATA][0] }), .west_out_b(
        \west_out_b[ACK] ) );
  input p_clk, n_clk, reset, \proc_in[MCMD][1] , \proc_in[MCMD][0] ,
         \proc_in[MADDR][31] , \proc_in[MADDR][30] , \proc_in[MADDR][29] ,
         \proc_in[MADDR][28] , \proc_in[MADDR][27] , \proc_in[MADDR][26] ,
         \proc_in[MADDR][25] , \proc_in[MADDR][24] , \proc_in[MADDR][23] ,
         \proc_in[MADDR][22] , \proc_in[MADDR][21] , \proc_in[MADDR][20] ,
         \proc_in[MADDR][19] , \proc_in[MADDR][18] , \proc_in[MADDR][17] ,
         \proc_in[MADDR][16] , \proc_in[MADDR][15] , \proc_in[MADDR][14] ,
         \proc_in[MADDR][13] , \proc_in[MADDR][12] , \proc_in[MADDR][11] ,
         \proc_in[MADDR][10] , \proc_in[MADDR][9] , \proc_in[MADDR][8] ,
         \proc_in[MADDR][7] , \proc_in[MADDR][6] , \proc_in[MADDR][5] ,
         \proc_in[MADDR][4] , \proc_in[MADDR][3] , \proc_in[MADDR][2] ,
         \proc_in[MADDR][1] , \proc_in[MADDR][0] , \proc_in[MDATA][31] ,
         \proc_in[MDATA][30] , \proc_in[MDATA][29] , \proc_in[MDATA][28] ,
         \proc_in[MDATA][27] , \proc_in[MDATA][26] , \proc_in[MDATA][25] ,
         \proc_in[MDATA][24] , \proc_in[MDATA][23] , \proc_in[MDATA][22] ,
         \proc_in[MDATA][21] , \proc_in[MDATA][20] , \proc_in[MDATA][19] ,
         \proc_in[MDATA][18] , \proc_in[MDATA][17] , \proc_in[MDATA][16] ,
         \proc_in[MDATA][15] , \proc_in[MDATA][14] , \proc_in[MDATA][13] ,
         \proc_in[MDATA][12] , \proc_in[MDATA][11] , \proc_in[MDATA][10] ,
         \proc_in[MDATA][9] , \proc_in[MDATA][8] , \proc_in[MDATA][7] ,
         \proc_in[MDATA][6] , \proc_in[MDATA][5] , \proc_in[MDATA][4] ,
         \proc_in[MDATA][3] , \proc_in[MDATA][2] , \proc_in[MDATA][1] ,
         \proc_in[MDATA][0] , \spm_in[SCMDACCEPT] , \spm_in[SRESP] ,
         \spm_in[SDATA][63] , \spm_in[SDATA][62] , \spm_in[SDATA][61] ,
         \spm_in[SDATA][60] , \spm_in[SDATA][59] , \spm_in[SDATA][58] ,
         \spm_in[SDATA][57] , \spm_in[SDATA][56] , \spm_in[SDATA][55] ,
         \spm_in[SDATA][54] , \spm_in[SDATA][53] , \spm_in[SDATA][52] ,
         \spm_in[SDATA][51] , \spm_in[SDATA][50] , \spm_in[SDATA][49] ,
         \spm_in[SDATA][48] , \spm_in[SDATA][47] , \spm_in[SDATA][46] ,
         \spm_in[SDATA][45] , \spm_in[SDATA][44] , \spm_in[SDATA][43] ,
         \spm_in[SDATA][42] , \spm_in[SDATA][41] , \spm_in[SDATA][40] ,
         \spm_in[SDATA][39] , \spm_in[SDATA][38] , \spm_in[SDATA][37] ,
         \spm_in[SDATA][36] , \spm_in[SDATA][35] , \spm_in[SDATA][34] ,
         \spm_in[SDATA][33] , \spm_in[SDATA][32] , \spm_in[SDATA][31] ,
         \spm_in[SDATA][30] , \spm_in[SDATA][29] , \spm_in[SDATA][28] ,
         \spm_in[SDATA][27] , \spm_in[SDATA][26] , \spm_in[SDATA][25] ,
         \spm_in[SDATA][24] , \spm_in[SDATA][23] , \spm_in[SDATA][22] ,
         \spm_in[SDATA][21] , \spm_in[SDATA][20] , \spm_in[SDATA][19] ,
         \spm_in[SDATA][18] , \spm_in[SDATA][17] , \spm_in[SDATA][16] ,
         \spm_in[SDATA][15] , \spm_in[SDATA][14] , \spm_in[SDATA][13] ,
         \spm_in[SDATA][12] , \spm_in[SDATA][11] , \spm_in[SDATA][10] ,
         \spm_in[SDATA][9] , \spm_in[SDATA][8] , \spm_in[SDATA][7] ,
         \spm_in[SDATA][6] , \spm_in[SDATA][5] , \spm_in[SDATA][4] ,
         \spm_in[SDATA][3] , \spm_in[SDATA][2] , \spm_in[SDATA][1] ,
         \spm_in[SDATA][0] , \north_in_f[REQ] , \north_in_f[DATA][34] ,
         \north_in_f[DATA][33] , \north_in_f[DATA][32] ,
         \north_in_f[DATA][31] , \north_in_f[DATA][30] ,
         \north_in_f[DATA][29] , \north_in_f[DATA][28] ,
         \north_in_f[DATA][27] , \north_in_f[DATA][26] ,
         \north_in_f[DATA][25] , \north_in_f[DATA][24] ,
         \north_in_f[DATA][23] , \north_in_f[DATA][22] ,
         \north_in_f[DATA][21] , \north_in_f[DATA][20] ,
         \north_in_f[DATA][19] , \north_in_f[DATA][18] ,
         \north_in_f[DATA][17] , \north_in_f[DATA][16] ,
         \north_in_f[DATA][15] , \north_in_f[DATA][14] ,
         \north_in_f[DATA][13] , \north_in_f[DATA][12] ,
         \north_in_f[DATA][11] , \north_in_f[DATA][10] , \north_in_f[DATA][9] ,
         \north_in_f[DATA][8] , \north_in_f[DATA][7] , \north_in_f[DATA][6] ,
         \north_in_f[DATA][5] , \north_in_f[DATA][4] , \north_in_f[DATA][3] ,
         \north_in_f[DATA][2] , \north_in_f[DATA][1] , \north_in_f[DATA][0] ,
         \east_in_f[REQ] , \east_in_f[DATA][34] , \east_in_f[DATA][33] ,
         \east_in_f[DATA][32] , \east_in_f[DATA][31] , \east_in_f[DATA][30] ,
         \east_in_f[DATA][29] , \east_in_f[DATA][28] , \east_in_f[DATA][27] ,
         \east_in_f[DATA][26] , \east_in_f[DATA][25] , \east_in_f[DATA][24] ,
         \east_in_f[DATA][23] , \east_in_f[DATA][22] , \east_in_f[DATA][21] ,
         \east_in_f[DATA][20] , \east_in_f[DATA][19] , \east_in_f[DATA][18] ,
         \east_in_f[DATA][17] , \east_in_f[DATA][16] , \east_in_f[DATA][15] ,
         \east_in_f[DATA][14] , \east_in_f[DATA][13] , \east_in_f[DATA][12] ,
         \east_in_f[DATA][11] , \east_in_f[DATA][10] , \east_in_f[DATA][9] ,
         \east_in_f[DATA][8] , \east_in_f[DATA][7] , \east_in_f[DATA][6] ,
         \east_in_f[DATA][5] , \east_in_f[DATA][4] , \east_in_f[DATA][3] ,
         \east_in_f[DATA][2] , \east_in_f[DATA][1] , \east_in_f[DATA][0] ,
         \south_in_f[REQ] , \south_in_f[DATA][34] , \south_in_f[DATA][33] ,
         \south_in_f[DATA][32] , \south_in_f[DATA][31] ,
         \south_in_f[DATA][30] , \south_in_f[DATA][29] ,
         \south_in_f[DATA][28] , \south_in_f[DATA][27] ,
         \south_in_f[DATA][26] , \south_in_f[DATA][25] ,
         \south_in_f[DATA][24] , \south_in_f[DATA][23] ,
         \south_in_f[DATA][22] , \south_in_f[DATA][21] ,
         \south_in_f[DATA][20] , \south_in_f[DATA][19] ,
         \south_in_f[DATA][18] , \south_in_f[DATA][17] ,
         \south_in_f[DATA][16] , \south_in_f[DATA][15] ,
         \south_in_f[DATA][14] , \south_in_f[DATA][13] ,
         \south_in_f[DATA][12] , \south_in_f[DATA][11] ,
         \south_in_f[DATA][10] , \south_in_f[DATA][9] , \south_in_f[DATA][8] ,
         \south_in_f[DATA][7] , \south_in_f[DATA][6] , \south_in_f[DATA][5] ,
         \south_in_f[DATA][4] , \south_in_f[DATA][3] , \south_in_f[DATA][2] ,
         \south_in_f[DATA][1] , \south_in_f[DATA][0] , \west_in_f[REQ] ,
         \west_in_f[DATA][34] , \west_in_f[DATA][33] , \west_in_f[DATA][32] ,
         \west_in_f[DATA][31] , \west_in_f[DATA][30] , \west_in_f[DATA][29] ,
         \west_in_f[DATA][28] , \west_in_f[DATA][27] , \west_in_f[DATA][26] ,
         \west_in_f[DATA][25] , \west_in_f[DATA][24] , \west_in_f[DATA][23] ,
         \west_in_f[DATA][22] , \west_in_f[DATA][21] , \west_in_f[DATA][20] ,
         \west_in_f[DATA][19] , \west_in_f[DATA][18] , \west_in_f[DATA][17] ,
         \west_in_f[DATA][16] , \west_in_f[DATA][15] , \west_in_f[DATA][14] ,
         \west_in_f[DATA][13] , \west_in_f[DATA][12] , \west_in_f[DATA][11] ,
         \west_in_f[DATA][10] , \west_in_f[DATA][9] , \west_in_f[DATA][8] ,
         \west_in_f[DATA][7] , \west_in_f[DATA][6] , \west_in_f[DATA][5] ,
         \west_in_f[DATA][4] , \west_in_f[DATA][3] , \west_in_f[DATA][2] ,
         \west_in_f[DATA][1] , \west_in_f[DATA][0] , \north_out_b[ACK] ,
         \east_out_b[ACK] , \south_out_b[ACK] , \west_out_b[ACK] ;
  output \proc_out[SCMDACCEPT] , \proc_out[SRESP] , \proc_out[SDATA][31] ,
         \proc_out[SDATA][30] , \proc_out[SDATA][29] , \proc_out[SDATA][28] ,
         \proc_out[SDATA][27] , \proc_out[SDATA][26] , \proc_out[SDATA][25] ,
         \proc_out[SDATA][24] , \proc_out[SDATA][23] , \proc_out[SDATA][22] ,
         \proc_out[SDATA][21] , \proc_out[SDATA][20] , \proc_out[SDATA][19] ,
         \proc_out[SDATA][18] , \proc_out[SDATA][17] , \proc_out[SDATA][16] ,
         \proc_out[SDATA][15] , \proc_out[SDATA][14] , \proc_out[SDATA][13] ,
         \proc_out[SDATA][12] , \proc_out[SDATA][11] , \proc_out[SDATA][10] ,
         \proc_out[SDATA][9] , \proc_out[SDATA][8] , \proc_out[SDATA][7] ,
         \proc_out[SDATA][6] , \proc_out[SDATA][5] , \proc_out[SDATA][4] ,
         \proc_out[SDATA][3] , \proc_out[SDATA][2] , \proc_out[SDATA][1] ,
         \proc_out[SDATA][0] , \spm_out[MCMD][1] , \spm_out[MCMD][0] ,
         \spm_out[MADDR][31] , \spm_out[MADDR][30] , \spm_out[MADDR][29] ,
         \spm_out[MADDR][28] , \spm_out[MADDR][27] , \spm_out[MADDR][26] ,
         \spm_out[MADDR][25] , \spm_out[MADDR][24] , \spm_out[MADDR][23] ,
         \spm_out[MADDR][22] , \spm_out[MADDR][21] , \spm_out[MADDR][20] ,
         \spm_out[MADDR][19] , \spm_out[MADDR][18] , \spm_out[MADDR][17] ,
         \spm_out[MADDR][16] , \spm_out[MADDR][15] , \spm_out[MADDR][14] ,
         \spm_out[MADDR][13] , \spm_out[MADDR][12] , \spm_out[MADDR][11] ,
         \spm_out[MADDR][10] , \spm_out[MADDR][9] , \spm_out[MADDR][8] ,
         \spm_out[MADDR][7] , \spm_out[MADDR][6] , \spm_out[MADDR][5] ,
         \spm_out[MADDR][4] , \spm_out[MADDR][3] , \spm_out[MADDR][2] ,
         \spm_out[MADDR][1] , \spm_out[MADDR][0] , \spm_out[MDATA][63] ,
         \spm_out[MDATA][62] , \spm_out[MDATA][61] , \spm_out[MDATA][60] ,
         \spm_out[MDATA][59] , \spm_out[MDATA][58] , \spm_out[MDATA][57] ,
         \spm_out[MDATA][56] , \spm_out[MDATA][55] , \spm_out[MDATA][54] ,
         \spm_out[MDATA][53] , \spm_out[MDATA][52] , \spm_out[MDATA][51] ,
         \spm_out[MDATA][50] , \spm_out[MDATA][49] , \spm_out[MDATA][48] ,
         \spm_out[MDATA][47] , \spm_out[MDATA][46] , \spm_out[MDATA][45] ,
         \spm_out[MDATA][44] , \spm_out[MDATA][43] , \spm_out[MDATA][42] ,
         \spm_out[MDATA][41] , \spm_out[MDATA][40] , \spm_out[MDATA][39] ,
         \spm_out[MDATA][38] , \spm_out[MDATA][37] , \spm_out[MDATA][36] ,
         \spm_out[MDATA][35] , \spm_out[MDATA][34] , \spm_out[MDATA][33] ,
         \spm_out[MDATA][32] , \spm_out[MDATA][31] , \spm_out[MDATA][30] ,
         \spm_out[MDATA][29] , \spm_out[MDATA][28] , \spm_out[MDATA][27] ,
         \spm_out[MDATA][26] , \spm_out[MDATA][25] , \spm_out[MDATA][24] ,
         \spm_out[MDATA][23] , \spm_out[MDATA][22] , \spm_out[MDATA][21] ,
         \spm_out[MDATA][20] , \spm_out[MDATA][19] , \spm_out[MDATA][18] ,
         \spm_out[MDATA][17] , \spm_out[MDATA][16] , \spm_out[MDATA][15] ,
         \spm_out[MDATA][14] , \spm_out[MDATA][13] , \spm_out[MDATA][12] ,
         \spm_out[MDATA][11] , \spm_out[MDATA][10] , \spm_out[MDATA][9] ,
         \spm_out[MDATA][8] , \spm_out[MDATA][7] , \spm_out[MDATA][6] ,
         \spm_out[MDATA][5] , \spm_out[MDATA][4] , \spm_out[MDATA][3] ,
         \spm_out[MDATA][2] , \spm_out[MDATA][1] , \spm_out[MDATA][0] ,
         \north_in_b[ACK] , \east_in_b[ACK] , \south_in_b[ACK] ,
         \west_in_b[ACK] , \north_out_f[REQ] , \north_out_f[DATA][34] ,
         \north_out_f[DATA][33] , \north_out_f[DATA][32] ,
         \north_out_f[DATA][31] , \north_out_f[DATA][30] ,
         \north_out_f[DATA][29] , \north_out_f[DATA][28] ,
         \north_out_f[DATA][27] , \north_out_f[DATA][26] ,
         \north_out_f[DATA][25] , \north_out_f[DATA][24] ,
         \north_out_f[DATA][23] , \north_out_f[DATA][22] ,
         \north_out_f[DATA][21] , \north_out_f[DATA][20] ,
         \north_out_f[DATA][19] , \north_out_f[DATA][18] ,
         \north_out_f[DATA][17] , \north_out_f[DATA][16] ,
         \north_out_f[DATA][15] , \north_out_f[DATA][14] ,
         \north_out_f[DATA][13] , \north_out_f[DATA][12] ,
         \north_out_f[DATA][11] , \north_out_f[DATA][10] ,
         \north_out_f[DATA][9] , \north_out_f[DATA][8] ,
         \north_out_f[DATA][7] , \north_out_f[DATA][6] ,
         \north_out_f[DATA][5] , \north_out_f[DATA][4] ,
         \north_out_f[DATA][3] , \north_out_f[DATA][2] ,
         \north_out_f[DATA][1] , \north_out_f[DATA][0] , \east_out_f[REQ] ,
         \east_out_f[DATA][34] , \east_out_f[DATA][33] ,
         \east_out_f[DATA][32] , \east_out_f[DATA][31] ,
         \east_out_f[DATA][30] , \east_out_f[DATA][29] ,
         \east_out_f[DATA][28] , \east_out_f[DATA][27] ,
         \east_out_f[DATA][26] , \east_out_f[DATA][25] ,
         \east_out_f[DATA][24] , \east_out_f[DATA][23] ,
         \east_out_f[DATA][22] , \east_out_f[DATA][21] ,
         \east_out_f[DATA][20] , \east_out_f[DATA][19] ,
         \east_out_f[DATA][18] , \east_out_f[DATA][17] ,
         \east_out_f[DATA][16] , \east_out_f[DATA][15] ,
         \east_out_f[DATA][14] , \east_out_f[DATA][13] ,
         \east_out_f[DATA][12] , \east_out_f[DATA][11] ,
         \east_out_f[DATA][10] , \east_out_f[DATA][9] , \east_out_f[DATA][8] ,
         \east_out_f[DATA][7] , \east_out_f[DATA][6] , \east_out_f[DATA][5] ,
         \east_out_f[DATA][4] , \east_out_f[DATA][3] , \east_out_f[DATA][2] ,
         \east_out_f[DATA][1] , \east_out_f[DATA][0] , \south_out_f[REQ] ,
         \south_out_f[DATA][34] , \south_out_f[DATA][33] ,
         \south_out_f[DATA][32] , \south_out_f[DATA][31] ,
         \south_out_f[DATA][30] , \south_out_f[DATA][29] ,
         \south_out_f[DATA][28] , \south_out_f[DATA][27] ,
         \south_out_f[DATA][26] , \south_out_f[DATA][25] ,
         \south_out_f[DATA][24] , \south_out_f[DATA][23] ,
         \south_out_f[DATA][22] , \south_out_f[DATA][21] ,
         \south_out_f[DATA][20] , \south_out_f[DATA][19] ,
         \south_out_f[DATA][18] , \south_out_f[DATA][17] ,
         \south_out_f[DATA][16] , \south_out_f[DATA][15] ,
         \south_out_f[DATA][14] , \south_out_f[DATA][13] ,
         \south_out_f[DATA][12] , \south_out_f[DATA][11] ,
         \south_out_f[DATA][10] , \south_out_f[DATA][9] ,
         \south_out_f[DATA][8] , \south_out_f[DATA][7] ,
         \south_out_f[DATA][6] , \south_out_f[DATA][5] ,
         \south_out_f[DATA][4] , \south_out_f[DATA][3] ,
         \south_out_f[DATA][2] , \south_out_f[DATA][1] ,
         \south_out_f[DATA][0] , \west_out_f[REQ] , \west_out_f[DATA][34] ,
         \west_out_f[DATA][33] , \west_out_f[DATA][32] ,
         \west_out_f[DATA][31] , \west_out_f[DATA][30] ,
         \west_out_f[DATA][29] , \west_out_f[DATA][28] ,
         \west_out_f[DATA][27] , \west_out_f[DATA][26] ,
         \west_out_f[DATA][25] , \west_out_f[DATA][24] ,
         \west_out_f[DATA][23] , \west_out_f[DATA][22] ,
         \west_out_f[DATA][21] , \west_out_f[DATA][20] ,
         \west_out_f[DATA][19] , \west_out_f[DATA][18] ,
         \west_out_f[DATA][17] , \west_out_f[DATA][16] ,
         \west_out_f[DATA][15] , \west_out_f[DATA][14] ,
         \west_out_f[DATA][13] , \west_out_f[DATA][12] ,
         \west_out_f[DATA][11] , \west_out_f[DATA][10] , \west_out_f[DATA][9] ,
         \west_out_f[DATA][8] , \west_out_f[DATA][7] , \west_out_f[DATA][6] ,
         \west_out_f[DATA][5] , \west_out_f[DATA][4] , \west_out_f[DATA][3] ,
         \west_out_f[DATA][2] , \west_out_f[DATA][1] , \west_out_f[DATA][0] ;
  wire   del_half_clk0, \ip_to_net_f[REQ] , n2, n1, n3, n4, n5, n6, n7, n8, n9,
         n10;
  wire   [34:0] net_to_ip;
  wire   [34:0] ip_to_net;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17;
  assign \spm_out[MADDR][31]  = 1'b0;
  assign \spm_out[MADDR][30]  = 1'b0;
  assign \spm_out[MADDR][29]  = 1'b0;
  assign \spm_out[MADDR][28]  = 1'b0;
  assign \spm_out[MADDR][27]  = 1'b0;
  assign \spm_out[MADDR][26]  = 1'b0;
  assign \spm_out[MADDR][25]  = 1'b0;
  assign \spm_out[MADDR][24]  = 1'b0;
  assign \spm_out[MADDR][23]  = 1'b0;
  assign \spm_out[MADDR][22]  = 1'b0;
  assign \spm_out[MADDR][21]  = 1'b0;
  assign \spm_out[MADDR][20]  = 1'b0;
  assign \spm_out[MADDR][19]  = 1'b0;
  assign \spm_out[MADDR][18]  = 1'b0;
  assign \spm_out[MADDR][17]  = 1'b0;
  assign \spm_out[MADDR][16]  = 1'b0;
  assign \spm_out[MADDR][15]  = 1'b0;

  nAdapter_0 na ( .na_clk(n_clk), .na_reset(reset), .proc_in({
        \proc_in[MCMD][1] , \proc_in[MCMD][0] , \proc_in[MADDR][31] , 
        \proc_in[MADDR][30] , \proc_in[MADDR][29] , \proc_in[MADDR][28] , 
        \proc_in[MADDR][27] , \proc_in[MADDR][26] , \proc_in[MADDR][25] , 
        \proc_in[MADDR][24] , \proc_in[MADDR][23] , \proc_in[MADDR][22] , 
        \proc_in[MADDR][21] , \proc_in[MADDR][20] , \proc_in[MADDR][19] , 
        \proc_in[MADDR][18] , \proc_in[MADDR][17] , \proc_in[MADDR][16] , 
        \proc_in[MADDR][15] , \proc_in[MADDR][14] , \proc_in[MADDR][13] , 
        \proc_in[MADDR][12] , \proc_in[MADDR][11] , \proc_in[MADDR][10] , 
        \proc_in[MADDR][9] , \proc_in[MADDR][8] , \proc_in[MADDR][7] , 
        \proc_in[MADDR][6] , \proc_in[MADDR][5] , \proc_in[MADDR][4] , 
        \proc_in[MADDR][3] , \proc_in[MADDR][2] , \proc_in[MADDR][1] , 
        \proc_in[MADDR][0] , \proc_in[MDATA][31] , \proc_in[MDATA][30] , 
        \proc_in[MDATA][29] , \proc_in[MDATA][28] , \proc_in[MDATA][27] , 
        \proc_in[MDATA][26] , \proc_in[MDATA][25] , \proc_in[MDATA][24] , 
        \proc_in[MDATA][23] , \proc_in[MDATA][22] , \proc_in[MDATA][21] , 
        \proc_in[MDATA][20] , \proc_in[MDATA][19] , \proc_in[MDATA][18] , 
        \proc_in[MDATA][17] , \proc_in[MDATA][16] , \proc_in[MDATA][15] , 
        \proc_in[MDATA][14] , \proc_in[MDATA][13] , \proc_in[MDATA][12] , 
        \proc_in[MDATA][11] , \proc_in[MDATA][10] , \proc_in[MDATA][9] , 
        \proc_in[MDATA][8] , \proc_in[MDATA][7] , \proc_in[MDATA][6] , 
        \proc_in[MDATA][5] , \proc_in[MDATA][4] , \proc_in[MDATA][3] , 
        \proc_in[MDATA][2] , \proc_in[MDATA][1] , \proc_in[MDATA][0] }), 
        .proc_out({\proc_out[SCMDACCEPT] , \proc_out[SRESP] , 
        \proc_out[SDATA][31] , \proc_out[SDATA][30] , \proc_out[SDATA][29] , 
        \proc_out[SDATA][28] , \proc_out[SDATA][27] , \proc_out[SDATA][26] , 
        \proc_out[SDATA][25] , \proc_out[SDATA][24] , \proc_out[SDATA][23] , 
        \proc_out[SDATA][22] , \proc_out[SDATA][21] , \proc_out[SDATA][20] , 
        \proc_out[SDATA][19] , \proc_out[SDATA][18] , \proc_out[SDATA][17] , 
        \proc_out[SDATA][16] , \proc_out[SDATA][15] , \proc_out[SDATA][14] , 
        \proc_out[SDATA][13] , \proc_out[SDATA][12] , \proc_out[SDATA][11] , 
        \proc_out[SDATA][10] , \proc_out[SDATA][9] , \proc_out[SDATA][8] , 
        \proc_out[SDATA][7] , \proc_out[SDATA][6] , \proc_out[SDATA][5] , 
        \proc_out[SDATA][4] , \proc_out[SDATA][3] , \proc_out[SDATA][2] , 
        \proc_out[SDATA][1] , \proc_out[SDATA][0] }), .spm_in({
        \spm_in[SCMDACCEPT] , \spm_in[SRESP] , \spm_in[SDATA][63] , 
        \spm_in[SDATA][62] , \spm_in[SDATA][61] , \spm_in[SDATA][60] , 
        \spm_in[SDATA][59] , \spm_in[SDATA][58] , \spm_in[SDATA][57] , 
        \spm_in[SDATA][56] , \spm_in[SDATA][55] , \spm_in[SDATA][54] , 
        \spm_in[SDATA][53] , \spm_in[SDATA][52] , \spm_in[SDATA][51] , 
        \spm_in[SDATA][50] , \spm_in[SDATA][49] , \spm_in[SDATA][48] , 
        \spm_in[SDATA][47] , \spm_in[SDATA][46] , \spm_in[SDATA][45] , 
        \spm_in[SDATA][44] , \spm_in[SDATA][43] , \spm_in[SDATA][42] , 
        \spm_in[SDATA][41] , \spm_in[SDATA][40] , \spm_in[SDATA][39] , 
        \spm_in[SDATA][38] , \spm_in[SDATA][37] , \spm_in[SDATA][36] , 
        \spm_in[SDATA][35] , \spm_in[SDATA][34] , \spm_in[SDATA][33] , 
        \spm_in[SDATA][32] , \spm_in[SDATA][31] , \spm_in[SDATA][30] , 
        \spm_in[SDATA][29] , \spm_in[SDATA][28] , \spm_in[SDATA][27] , 
        \spm_in[SDATA][26] , \spm_in[SDATA][25] , \spm_in[SDATA][24] , 
        \spm_in[SDATA][23] , \spm_in[SDATA][22] , \spm_in[SDATA][21] , 
        \spm_in[SDATA][20] , \spm_in[SDATA][19] , \spm_in[SDATA][18] , 
        \spm_in[SDATA][17] , \spm_in[SDATA][16] , \spm_in[SDATA][15] , 
        \spm_in[SDATA][14] , \spm_in[SDATA][13] , \spm_in[SDATA][12] , 
        \spm_in[SDATA][11] , \spm_in[SDATA][10] , \spm_in[SDATA][9] , 
        \spm_in[SDATA][8] , \spm_in[SDATA][7] , \spm_in[SDATA][6] , 
        \spm_in[SDATA][5] , \spm_in[SDATA][4] , \spm_in[SDATA][3] , 
        \spm_in[SDATA][2] , \spm_in[SDATA][1] , \spm_in[SDATA][0] }), 
        .spm_out({\spm_out[MCMD][1] , \spm_out[MCMD][0] , 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, \spm_out[MADDR][14] , \spm_out[MADDR][13] , 
        \spm_out[MADDR][12] , \spm_out[MADDR][11] , \spm_out[MADDR][10] , 
        \spm_out[MADDR][9] , \spm_out[MADDR][8] , \spm_out[MADDR][7] , 
        \spm_out[MADDR][6] , \spm_out[MADDR][5] , \spm_out[MADDR][4] , 
        \spm_out[MADDR][3] , \spm_out[MADDR][2] , \spm_out[MADDR][1] , 
        \spm_out[MADDR][0] , \spm_out[MDATA][63] , \spm_out[MDATA][62] , 
        \spm_out[MDATA][61] , \spm_out[MDATA][60] , \spm_out[MDATA][59] , 
        \spm_out[MDATA][58] , \spm_out[MDATA][57] , \spm_out[MDATA][56] , 
        \spm_out[MDATA][55] , \spm_out[MDATA][54] , \spm_out[MDATA][53] , 
        \spm_out[MDATA][52] , \spm_out[MDATA][51] , \spm_out[MDATA][50] , 
        \spm_out[MDATA][49] , \spm_out[MDATA][48] , \spm_out[MDATA][47] , 
        \spm_out[MDATA][46] , \spm_out[MDATA][45] , \spm_out[MDATA][44] , 
        \spm_out[MDATA][43] , \spm_out[MDATA][42] , \spm_out[MDATA][41] , 
        \spm_out[MDATA][40] , \spm_out[MDATA][39] , \spm_out[MDATA][38] , 
        \spm_out[MDATA][37] , \spm_out[MDATA][36] , \spm_out[MDATA][35] , 
        \spm_out[MDATA][34] , \spm_out[MDATA][33] , \spm_out[MDATA][32] , 
        \spm_out[MDATA][31] , \spm_out[MDATA][30] , \spm_out[MDATA][29] , 
        \spm_out[MDATA][28] , \spm_out[MDATA][27] , \spm_out[MDATA][26] , 
        \spm_out[MDATA][25] , \spm_out[MDATA][24] , \spm_out[MDATA][23] , 
        \spm_out[MDATA][22] , \spm_out[MDATA][21] , \spm_out[MDATA][20] , 
        \spm_out[MDATA][19] , \spm_out[MDATA][18] , \spm_out[MDATA][17] , 
        \spm_out[MDATA][16] , \spm_out[MDATA][15] , \spm_out[MDATA][14] , 
        \spm_out[MDATA][13] , \spm_out[MDATA][12] , \spm_out[MDATA][11] , 
        \spm_out[MDATA][10] , \spm_out[MDATA][9] , \spm_out[MDATA][8] , 
        \spm_out[MDATA][7] , \spm_out[MDATA][6] , \spm_out[MDATA][5] , 
        \spm_out[MDATA][4] , \spm_out[MDATA][3] , \spm_out[MDATA][2] , 
        \spm_out[MDATA][1] , \spm_out[MDATA][0] }), .pkt_in(net_to_ip), 
        .pkt_out(ip_to_net) );
  noc_switch_0 r ( .preset(reset), .north_in_f({\north_in_f[REQ] , 
        \north_in_f[DATA][34] , \north_in_f[DATA][33] , \north_in_f[DATA][32] , 
        \north_in_f[DATA][31] , \north_in_f[DATA][30] , \north_in_f[DATA][29] , 
        \north_in_f[DATA][28] , \north_in_f[DATA][27] , \north_in_f[DATA][26] , 
        \north_in_f[DATA][25] , \north_in_f[DATA][24] , \north_in_f[DATA][23] , 
        \north_in_f[DATA][22] , \north_in_f[DATA][21] , \north_in_f[DATA][20] , 
        \north_in_f[DATA][19] , \north_in_f[DATA][18] , \north_in_f[DATA][17] , 
        \north_in_f[DATA][16] , \north_in_f[DATA][15] , \north_in_f[DATA][14] , 
        \north_in_f[DATA][13] , \north_in_f[DATA][12] , \north_in_f[DATA][11] , 
        \north_in_f[DATA][10] , \north_in_f[DATA][9] , \north_in_f[DATA][8] , 
        \north_in_f[DATA][7] , \north_in_f[DATA][6] , \north_in_f[DATA][5] , 
        \north_in_f[DATA][4] , \north_in_f[DATA][3] , \north_in_f[DATA][2] , 
        \north_in_f[DATA][1] , \north_in_f[DATA][0] }), .north_in_b(
        \north_in_b[ACK] ), .east_in_f({\east_in_f[REQ] , 
        \east_in_f[DATA][34] , \east_in_f[DATA][33] , \east_in_f[DATA][32] , 
        \east_in_f[DATA][31] , \east_in_f[DATA][30] , \east_in_f[DATA][29] , 
        \east_in_f[DATA][28] , \east_in_f[DATA][27] , \east_in_f[DATA][26] , 
        \east_in_f[DATA][25] , \east_in_f[DATA][24] , \east_in_f[DATA][23] , 
        \east_in_f[DATA][22] , \east_in_f[DATA][21] , \east_in_f[DATA][20] , 
        \east_in_f[DATA][19] , \east_in_f[DATA][18] , \east_in_f[DATA][17] , 
        \east_in_f[DATA][16] , \east_in_f[DATA][15] , \east_in_f[DATA][14] , 
        \east_in_f[DATA][13] , \east_in_f[DATA][12] , \east_in_f[DATA][11] , 
        \east_in_f[DATA][10] , \east_in_f[DATA][9] , \east_in_f[DATA][8] , 
        \east_in_f[DATA][7] , \east_in_f[DATA][6] , \east_in_f[DATA][5] , 
        \east_in_f[DATA][4] , \east_in_f[DATA][3] , \east_in_f[DATA][2] , 
        \east_in_f[DATA][1] , \east_in_f[DATA][0] }), .east_in_b(
        \east_in_b[ACK] ), .south_in_f({\south_in_f[REQ] , 
        \south_in_f[DATA][34] , \south_in_f[DATA][33] , \south_in_f[DATA][32] , 
        \south_in_f[DATA][31] , \south_in_f[DATA][30] , \south_in_f[DATA][29] , 
        \south_in_f[DATA][28] , \south_in_f[DATA][27] , \south_in_f[DATA][26] , 
        \south_in_f[DATA][25] , \south_in_f[DATA][24] , \south_in_f[DATA][23] , 
        \south_in_f[DATA][22] , \south_in_f[DATA][21] , \south_in_f[DATA][20] , 
        \south_in_f[DATA][19] , \south_in_f[DATA][18] , \south_in_f[DATA][17] , 
        \south_in_f[DATA][16] , \south_in_f[DATA][15] , \south_in_f[DATA][14] , 
        \south_in_f[DATA][13] , \south_in_f[DATA][12] , \south_in_f[DATA][11] , 
        \south_in_f[DATA][10] , \south_in_f[DATA][9] , \south_in_f[DATA][8] , 
        \south_in_f[DATA][7] , \south_in_f[DATA][6] , \south_in_f[DATA][5] , 
        \south_in_f[DATA][4] , \south_in_f[DATA][3] , \south_in_f[DATA][2] , 
        \south_in_f[DATA][1] , \south_in_f[DATA][0] }), .south_in_b(
        \south_in_b[ACK] ), .west_in_f({\west_in_f[REQ] , 
        \west_in_f[DATA][34] , \west_in_f[DATA][33] , \west_in_f[DATA][32] , 
        \west_in_f[DATA][31] , \west_in_f[DATA][30] , \west_in_f[DATA][29] , 
        \west_in_f[DATA][28] , \west_in_f[DATA][27] , \west_in_f[DATA][26] , 
        \west_in_f[DATA][25] , \west_in_f[DATA][24] , \west_in_f[DATA][23] , 
        \west_in_f[DATA][22] , \west_in_f[DATA][21] , \west_in_f[DATA][20] , 
        \west_in_f[DATA][19] , \west_in_f[DATA][18] , \west_in_f[DATA][17] , 
        \west_in_f[DATA][16] , \west_in_f[DATA][15] , \west_in_f[DATA][14] , 
        \west_in_f[DATA][13] , \west_in_f[DATA][12] , \west_in_f[DATA][11] , 
        \west_in_f[DATA][10] , \west_in_f[DATA][9] , \west_in_f[DATA][8] , 
        \west_in_f[DATA][7] , \west_in_f[DATA][6] , \west_in_f[DATA][5] , 
        \west_in_f[DATA][4] , \west_in_f[DATA][3] , \west_in_f[DATA][2] , 
        \west_in_f[DATA][1] , \west_in_f[DATA][0] }), .west_in_b(
        \west_in_b[ACK] ), .resource_in_f({\ip_to_net_f[REQ] , ip_to_net}), 
        .north_out_f({\north_out_f[REQ] , \north_out_f[DATA][34] , 
        \north_out_f[DATA][33] , \north_out_f[DATA][32] , 
        \north_out_f[DATA][31] , \north_out_f[DATA][30] , 
        \north_out_f[DATA][29] , \north_out_f[DATA][28] , 
        \north_out_f[DATA][27] , \north_out_f[DATA][26] , 
        \north_out_f[DATA][25] , \north_out_f[DATA][24] , 
        \north_out_f[DATA][23] , \north_out_f[DATA][22] , 
        \north_out_f[DATA][21] , \north_out_f[DATA][20] , 
        \north_out_f[DATA][19] , \north_out_f[DATA][18] , 
        \north_out_f[DATA][17] , \north_out_f[DATA][16] , 
        \north_out_f[DATA][15] , \north_out_f[DATA][14] , 
        \north_out_f[DATA][13] , \north_out_f[DATA][12] , 
        \north_out_f[DATA][11] , \north_out_f[DATA][10] , 
        \north_out_f[DATA][9] , \north_out_f[DATA][8] , \north_out_f[DATA][7] , 
        \north_out_f[DATA][6] , \north_out_f[DATA][5] , \north_out_f[DATA][4] , 
        \north_out_f[DATA][3] , \north_out_f[DATA][2] , \north_out_f[DATA][1] , 
        \north_out_f[DATA][0] }), .north_out_b(\north_out_b[ACK] ), 
        .east_out_f({\east_out_f[REQ] , \east_out_f[DATA][34] , 
        \east_out_f[DATA][33] , \east_out_f[DATA][32] , \east_out_f[DATA][31] , 
        \east_out_f[DATA][30] , \east_out_f[DATA][29] , \east_out_f[DATA][28] , 
        \east_out_f[DATA][27] , \east_out_f[DATA][26] , \east_out_f[DATA][25] , 
        \east_out_f[DATA][24] , \east_out_f[DATA][23] , \east_out_f[DATA][22] , 
        \east_out_f[DATA][21] , \east_out_f[DATA][20] , \east_out_f[DATA][19] , 
        \east_out_f[DATA][18] , \east_out_f[DATA][17] , \east_out_f[DATA][16] , 
        \east_out_f[DATA][15] , \east_out_f[DATA][14] , \east_out_f[DATA][13] , 
        \east_out_f[DATA][12] , \east_out_f[DATA][11] , \east_out_f[DATA][10] , 
        \east_out_f[DATA][9] , \east_out_f[DATA][8] , \east_out_f[DATA][7] , 
        \east_out_f[DATA][6] , \east_out_f[DATA][5] , \east_out_f[DATA][4] , 
        \east_out_f[DATA][3] , \east_out_f[DATA][2] , \east_out_f[DATA][1] , 
        \east_out_f[DATA][0] }), .east_out_b(\east_out_b[ACK] ), .south_out_f(
        {\south_out_f[REQ] , \south_out_f[DATA][34] , \south_out_f[DATA][33] , 
        \south_out_f[DATA][32] , \south_out_f[DATA][31] , 
        \south_out_f[DATA][30] , \south_out_f[DATA][29] , 
        \south_out_f[DATA][28] , \south_out_f[DATA][27] , 
        \south_out_f[DATA][26] , \south_out_f[DATA][25] , 
        \south_out_f[DATA][24] , \south_out_f[DATA][23] , 
        \south_out_f[DATA][22] , \south_out_f[DATA][21] , 
        \south_out_f[DATA][20] , \south_out_f[DATA][19] , 
        \south_out_f[DATA][18] , \south_out_f[DATA][17] , 
        \south_out_f[DATA][16] , \south_out_f[DATA][15] , 
        \south_out_f[DATA][14] , \south_out_f[DATA][13] , 
        \south_out_f[DATA][12] , \south_out_f[DATA][11] , 
        \south_out_f[DATA][10] , \south_out_f[DATA][9] , 
        \south_out_f[DATA][8] , \south_out_f[DATA][7] , \south_out_f[DATA][6] , 
        \south_out_f[DATA][5] , \south_out_f[DATA][4] , \south_out_f[DATA][3] , 
        \south_out_f[DATA][2] , \south_out_f[DATA][1] , \south_out_f[DATA][0] }), .south_out_b(\south_out_b[ACK] ), .west_out_f({\west_out_f[REQ] , 
        \west_out_f[DATA][34] , \west_out_f[DATA][33] , \west_out_f[DATA][32] , 
        \west_out_f[DATA][31] , \west_out_f[DATA][30] , \west_out_f[DATA][29] , 
        \west_out_f[DATA][28] , \west_out_f[DATA][27] , \west_out_f[DATA][26] , 
        \west_out_f[DATA][25] , \west_out_f[DATA][24] , \west_out_f[DATA][23] , 
        \west_out_f[DATA][22] , \west_out_f[DATA][21] , \west_out_f[DATA][20] , 
        \west_out_f[DATA][19] , \west_out_f[DATA][18] , \west_out_f[DATA][17] , 
        \west_out_f[DATA][16] , \west_out_f[DATA][15] , \west_out_f[DATA][14] , 
        \west_out_f[DATA][13] , \west_out_f[DATA][12] , \west_out_f[DATA][11] , 
        \west_out_f[DATA][10] , \west_out_f[DATA][9] , \west_out_f[DATA][8] , 
        \west_out_f[DATA][7] , \west_out_f[DATA][6] , \west_out_f[DATA][5] , 
        \west_out_f[DATA][4] , \west_out_f[DATA][3] , \west_out_f[DATA][2] , 
        \west_out_f[DATA][1] , \west_out_f[DATA][0] }), .west_out_b(
        \west_out_b[ACK] ), .resource_out_f({SYNOPSYS_UNCONNECTED__17, 
        net_to_ip}), .resource_out_b(n9) );
  HS65_LS_DFPRQNX9 half_clk_reg ( .D(n2), .CP(n_clk), .RN(n8), .QN(n2) );
  HS65_LS_IVX9 I_2 ( .A(n4), .Z(\ip_to_net_f[REQ] ) );
  HS65_LH_IVX2 I_1 ( .A(n10), .Z(del_half_clk0) );
  HS65_LS_IVX9 U3 ( .A(n2), .Z(n10) );
  HS65_LH_IVX2 U4 ( .A(n1), .Z(n3) );
  HS65_LS_IVX106 U5 ( .A(del_half_clk0), .Z(n1) );
  HS65_LS_BFX9 U6 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U7 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U8 ( .A(n7), .Z(n6) );
  HS65_LS_BFX9 U9 ( .A(n3), .Z(n7) );
  HS65_LS_IVX9 U10 ( .A(reset), .Z(n8) );
  HS65_LS_IVX9 U11 ( .A(del_half_clk0), .Z(n9) );
endmodule


module counter_WIDTH3_3 ( clk, reset, enable, cnt );
  output [2:0] cnt;
  input clk, reset, enable;
  wire   n1, n2, n3, n4, n5, n8, n9, n10, n11;

  HS65_LS_DFPRQX9 \reg_reg[0]  ( .D(n5), .CP(clk), .RN(n1), .Q(cnt[0]) );
  HS65_LS_DFPRQX9 \reg_reg[2]  ( .D(n8), .CP(clk), .RN(n1), .Q(cnt[2]) );
  HS65_LS_DFPRQX9 \reg_reg[1]  ( .D(n9), .CP(clk), .RN(n1), .Q(cnt[1]) );
  HS65_LS_IVX9 U3 ( .A(reset), .Z(n1) );
  HS65_LS_OAI32X5 U4 ( .A(n4), .B(n11), .C(n2), .D(enable), .E(n3), .Z(n8) );
  HS65_LS_NAND2X7 U5 ( .A(enable), .B(n3), .Z(n11) );
  HS65_LS_OAI32X5 U6 ( .A(n2), .B(cnt[1]), .C(n11), .D(n10), .E(n4), .Z(n9) );
  HS65_LS_OA12X9 U7 ( .A(cnt[0]), .B(cnt[2]), .C(enable), .Z(n10) );
  HS65_LS_OAI22X6 U8 ( .A(enable), .B(n2), .C(cnt[0]), .D(n11), .Z(n5) );
  HS65_LS_IVX9 U9 ( .A(cnt[0]), .Z(n2) );
  HS65_LS_IVX9 U10 ( .A(cnt[1]), .Z(n4) );
  HS65_LS_IVX9 U11 ( .A(cnt[2]), .Z(n3) );
endmodule


module bram_DATA16_ADDR2_6 ( clk, reset, rd_addr, wr_addr, wr_data, wr_ena, 
        rd_data );
  input [1:0] rd_addr;
  input [1:0] wr_addr;
  input [15:0] wr_data;
  output [15:0] rd_data;
  input clk, reset, wr_ena;
  wire   \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] ,
         \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][15] , \mem[1][14] , \mem[1][13] ,
         \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] , \mem[1][8] ,
         \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] ,
         \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][15] , \mem[0][14] ,
         \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] ,
         \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] ,
         \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, n1,
         n2, n3, n4, n5, n6, n7, n8, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162;

  HS65_LS_DFPRQX9 \mem_reg[3][15]  ( .D(n91), .CP(clk), .RN(n1), .Q(
        \mem[3][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][14]  ( .D(n92), .CP(clk), .RN(n1), .Q(
        \mem[3][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][13]  ( .D(n93), .CP(clk), .RN(n1), .Q(
        \mem[3][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][12]  ( .D(n94), .CP(clk), .RN(n1), .Q(
        \mem[3][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][11]  ( .D(n95), .CP(clk), .RN(n1), .Q(
        \mem[3][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][10]  ( .D(n96), .CP(clk), .RN(n1), .Q(
        \mem[3][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][9]  ( .D(n97), .CP(clk), .RN(n1), .Q(\mem[3][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][8]  ( .D(n98), .CP(clk), .RN(n1), .Q(\mem[3][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][7]  ( .D(n99), .CP(clk), .RN(n1), .Q(\mem[3][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][6]  ( .D(n100), .CP(clk), .RN(n1), .Q(
        \mem[3][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][5]  ( .D(n101), .CP(clk), .RN(n1), .Q(
        \mem[3][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][4]  ( .D(n102), .CP(clk), .RN(n1), .Q(
        \mem[3][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][3]  ( .D(n103), .CP(clk), .RN(n1), .Q(
        \mem[3][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][2]  ( .D(n104), .CP(clk), .RN(n2), .Q(
        \mem[3][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][1]  ( .D(n105), .CP(clk), .RN(n2), .Q(
        \mem[3][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][0]  ( .D(n106), .CP(clk), .RN(n2), .Q(
        \mem[3][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][15]  ( .D(n107), .CP(clk), .RN(n2), .Q(
        \mem[2][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][14]  ( .D(n108), .CP(clk), .RN(n2), .Q(
        \mem[2][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][13]  ( .D(n109), .CP(clk), .RN(n2), .Q(
        \mem[2][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][12]  ( .D(n110), .CP(clk), .RN(n2), .Q(
        \mem[2][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][11]  ( .D(n111), .CP(clk), .RN(n2), .Q(
        \mem[2][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][10]  ( .D(n112), .CP(clk), .RN(n2), .Q(
        \mem[2][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][9]  ( .D(n113), .CP(clk), .RN(n2), .Q(
        \mem[2][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][8]  ( .D(n114), .CP(clk), .RN(n2), .Q(
        \mem[2][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][7]  ( .D(n115), .CP(clk), .RN(n2), .Q(
        \mem[2][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][6]  ( .D(n116), .CP(clk), .RN(n2), .Q(
        \mem[2][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][5]  ( .D(n117), .CP(clk), .RN(n3), .Q(
        \mem[2][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][4]  ( .D(n118), .CP(clk), .RN(n3), .Q(
        \mem[2][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][3]  ( .D(n119), .CP(clk), .RN(n3), .Q(
        \mem[2][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][2]  ( .D(n120), .CP(clk), .RN(n3), .Q(
        \mem[2][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][1]  ( .D(n121), .CP(clk), .RN(n3), .Q(
        \mem[2][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][0]  ( .D(n122), .CP(clk), .RN(n3), .Q(
        \mem[2][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][15]  ( .D(n123), .CP(clk), .RN(n3), .Q(
        \mem[1][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][14]  ( .D(n124), .CP(clk), .RN(n3), .Q(
        \mem[1][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][13]  ( .D(n125), .CP(clk), .RN(n3), .Q(
        \mem[1][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][12]  ( .D(n126), .CP(clk), .RN(n3), .Q(
        \mem[1][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][11]  ( .D(n127), .CP(clk), .RN(n3), .Q(
        \mem[1][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][10]  ( .D(n128), .CP(clk), .RN(n3), .Q(
        \mem[1][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][9]  ( .D(n129), .CP(clk), .RN(n3), .Q(
        \mem[1][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][8]  ( .D(n130), .CP(clk), .RN(n4), .Q(
        \mem[1][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][7]  ( .D(n131), .CP(clk), .RN(n4), .Q(
        \mem[1][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][6]  ( .D(n132), .CP(clk), .RN(n4), .Q(
        \mem[1][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][5]  ( .D(n133), .CP(clk), .RN(n4), .Q(
        \mem[1][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][4]  ( .D(n134), .CP(clk), .RN(n4), .Q(
        \mem[1][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][3]  ( .D(n135), .CP(clk), .RN(n4), .Q(
        \mem[1][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][2]  ( .D(n136), .CP(clk), .RN(n4), .Q(
        \mem[1][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][1]  ( .D(n137), .CP(clk), .RN(n4), .Q(
        \mem[1][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][0]  ( .D(n138), .CP(clk), .RN(n4), .Q(
        \mem[1][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][15]  ( .D(n139), .CP(clk), .RN(n4), .Q(
        \mem[0][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][14]  ( .D(n140), .CP(clk), .RN(n4), .Q(
        \mem[0][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][13]  ( .D(n141), .CP(clk), .RN(n4), .Q(
        \mem[0][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][12]  ( .D(n142), .CP(clk), .RN(n4), .Q(
        \mem[0][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][11]  ( .D(n143), .CP(clk), .RN(n5), .Q(
        \mem[0][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][10]  ( .D(n144), .CP(clk), .RN(n5), .Q(
        \mem[0][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][9]  ( .D(n145), .CP(clk), .RN(n5), .Q(
        \mem[0][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][8]  ( .D(n146), .CP(clk), .RN(n5), .Q(
        \mem[0][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][7]  ( .D(n147), .CP(clk), .RN(n5), .Q(
        \mem[0][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][6]  ( .D(n148), .CP(clk), .RN(n5), .Q(
        \mem[0][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][5]  ( .D(n149), .CP(clk), .RN(n5), .Q(
        \mem[0][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][4]  ( .D(n150), .CP(clk), .RN(n5), .Q(
        \mem[0][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][3]  ( .D(n151), .CP(clk), .RN(n5), .Q(
        \mem[0][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][2]  ( .D(n152), .CP(clk), .RN(n5), .Q(
        \mem[0][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][1]  ( .D(n153), .CP(clk), .RN(n5), .Q(
        \mem[0][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][0]  ( .D(n154), .CP(clk), .RN(n5), .Q(
        \mem[0][0] ) );
  HS65_LS_DFPRQX9 \rd_data_reg[15]  ( .D(N17), .CP(clk), .RN(n5), .Q(
        rd_data[15]) );
  HS65_LS_DFPRQX9 \rd_data_reg[14]  ( .D(N18), .CP(clk), .RN(n6), .Q(
        rd_data[14]) );
  HS65_LS_DFPRQX9 \rd_data_reg[13]  ( .D(N19), .CP(clk), .RN(n6), .Q(
        rd_data[13]) );
  HS65_LS_DFPRQX9 \rd_data_reg[12]  ( .D(N20), .CP(clk), .RN(n6), .Q(
        rd_data[12]) );
  HS65_LS_DFPRQX9 \rd_data_reg[11]  ( .D(N21), .CP(clk), .RN(n6), .Q(
        rd_data[11]) );
  HS65_LS_DFPRQX9 \rd_data_reg[10]  ( .D(N22), .CP(clk), .RN(n6), .Q(
        rd_data[10]) );
  HS65_LS_DFPRQX9 \rd_data_reg[9]  ( .D(N23), .CP(clk), .RN(n6), .Q(rd_data[9]) );
  HS65_LS_DFPRQX9 \rd_data_reg[8]  ( .D(N24), .CP(clk), .RN(n6), .Q(rd_data[8]) );
  HS65_LS_DFPRQX9 \rd_data_reg[7]  ( .D(N25), .CP(clk), .RN(n6), .Q(rd_data[7]) );
  HS65_LS_DFPRQX9 \rd_data_reg[6]  ( .D(N26), .CP(clk), .RN(n6), .Q(rd_data[6]) );
  HS65_LS_DFPRQX9 \rd_data_reg[5]  ( .D(N27), .CP(clk), .RN(n6), .Q(rd_data[5]) );
  HS65_LS_DFPRQX9 \rd_data_reg[4]  ( .D(N28), .CP(clk), .RN(n6), .Q(rd_data[4]) );
  HS65_LS_DFPRQX9 \rd_data_reg[3]  ( .D(N29), .CP(clk), .RN(n6), .Q(rd_data[3]) );
  HS65_LS_DFPRQX9 \rd_data_reg[2]  ( .D(N30), .CP(clk), .RN(n6), .Q(rd_data[2]) );
  HS65_LS_DFPRQX9 \rd_data_reg[1]  ( .D(N31), .CP(clk), .RN(n7), .Q(rd_data[1]) );
  HS65_LS_DFPRQX9 \rd_data_reg[0]  ( .D(N32), .CP(clk), .RN(n7), .Q(rd_data[0]) );
  HS65_LS_BFX9 U3 ( .A(n81), .Z(n4) );
  HS65_LS_BFX9 U4 ( .A(n81), .Z(n3) );
  HS65_LS_BFX9 U5 ( .A(n81), .Z(n2) );
  HS65_LS_BFX9 U6 ( .A(n83), .Z(n81) );
  HS65_LS_BFX9 U7 ( .A(n8), .Z(n6) );
  HS65_LS_BFX9 U8 ( .A(n8), .Z(n5) );
  HS65_LS_BFX9 U9 ( .A(n82), .Z(n1) );
  HS65_LS_BFX9 U10 ( .A(n83), .Z(n82) );
  HS65_LS_BFX9 U11 ( .A(n8), .Z(n7) );
  HS65_LS_BFX9 U12 ( .A(n83), .Z(n8) );
  HS65_LS_IVX9 U13 ( .A(reset), .Z(n83) );
  HS65_LS_IVX9 U14 ( .A(n161), .Z(n86) );
  HS65_LS_IVX9 U15 ( .A(n162), .Z(n87) );
  HS65_LS_NAND3X5 U16 ( .A(wr_ena), .B(n88), .C(wr_addr[0]), .Z(n161) );
  HS65_LS_IVX9 U17 ( .A(wr_addr[0]), .Z(n89) );
  HS65_LS_NAND3X5 U18 ( .A(n89), .B(n88), .C(wr_ena), .Z(n162) );
  HS65_LS_IVX9 U19 ( .A(n160), .Z(n85) );
  HS65_LS_IVX9 U20 ( .A(n159), .Z(n84) );
  HS65_LS_NAND3X5 U21 ( .A(wr_ena), .B(n89), .C(wr_addr[1]), .Z(n160) );
  HS65_LS_NOR2X6 U22 ( .A(n90), .B(rd_addr[1]), .Z(n157) );
  HS65_LS_NOR2X6 U23 ( .A(rd_addr[0]), .B(rd_addr[1]), .Z(n158) );
  HS65_LS_IVX9 U24 ( .A(wr_addr[1]), .Z(n88) );
  HS65_LS_NAND3X5 U25 ( .A(wr_addr[0]), .B(wr_ena), .C(wr_addr[1]), .Z(n159)
         );
  HS65_LS_AND2X4 U26 ( .A(rd_addr[1]), .B(n90), .Z(n156) );
  HS65_LS_AND2X4 U27 ( .A(rd_addr[1]), .B(rd_addr[0]), .Z(n155) );
  HS65_LS_IVX9 U28 ( .A(rd_addr[0]), .Z(n90) );
  HS65_LS_MX41X7 U29 ( .D0(n158), .S0(\mem[0][0] ), .D1(n157), .S1(\mem[1][0] ), .D2(n156), .S2(\mem[2][0] ), .D3(n155), .S3(\mem[3][0] ), .Z(N32) );
  HS65_LS_MX41X7 U30 ( .D0(n158), .S0(\mem[0][1] ), .D1(n157), .S1(\mem[1][1] ), .D2(n156), .S2(\mem[2][1] ), .D3(n155), .S3(\mem[3][1] ), .Z(N31) );
  HS65_LS_MX41X7 U31 ( .D0(n158), .S0(\mem[0][2] ), .D1(n157), .S1(\mem[1][2] ), .D2(n156), .S2(\mem[2][2] ), .D3(n155), .S3(\mem[3][2] ), .Z(N30) );
  HS65_LS_MX41X7 U32 ( .D0(n158), .S0(\mem[0][3] ), .D1(n157), .S1(\mem[1][3] ), .D2(n156), .S2(\mem[2][3] ), .D3(n155), .S3(\mem[3][3] ), .Z(N29) );
  HS65_LS_MX41X7 U33 ( .D0(n158), .S0(\mem[0][4] ), .D1(n157), .S1(\mem[1][4] ), .D2(n156), .S2(\mem[2][4] ), .D3(n155), .S3(\mem[3][4] ), .Z(N28) );
  HS65_LS_MX41X7 U34 ( .D0(n158), .S0(\mem[0][5] ), .D1(n157), .S1(\mem[1][5] ), .D2(n156), .S2(\mem[2][5] ), .D3(n155), .S3(\mem[3][5] ), .Z(N27) );
  HS65_LS_MX41X7 U35 ( .D0(n158), .S0(\mem[0][6] ), .D1(n157), .S1(\mem[1][6] ), .D2(n156), .S2(\mem[2][6] ), .D3(n155), .S3(\mem[3][6] ), .Z(N26) );
  HS65_LS_MX41X7 U36 ( .D0(n158), .S0(\mem[0][7] ), .D1(n157), .S1(\mem[1][7] ), .D2(n156), .S2(\mem[2][7] ), .D3(n155), .S3(\mem[3][7] ), .Z(N25) );
  HS65_LS_MX41X7 U37 ( .D0(n158), .S0(\mem[0][8] ), .D1(n157), .S1(\mem[1][8] ), .D2(n156), .S2(\mem[2][8] ), .D3(n155), .S3(\mem[3][8] ), .Z(N24) );
  HS65_LS_MX41X7 U38 ( .D0(n158), .S0(\mem[0][9] ), .D1(n157), .S1(\mem[1][9] ), .D2(n156), .S2(\mem[2][9] ), .D3(n155), .S3(\mem[3][9] ), .Z(N23) );
  HS65_LS_MX41X7 U39 ( .D0(n158), .S0(\mem[0][10] ), .D1(n157), .S1(
        \mem[1][10] ), .D2(n156), .S2(\mem[2][10] ), .D3(n155), .S3(
        \mem[3][10] ), .Z(N22) );
  HS65_LS_MX41X7 U40 ( .D0(n158), .S0(\mem[0][11] ), .D1(n157), .S1(
        \mem[1][11] ), .D2(n156), .S2(\mem[2][11] ), .D3(n155), .S3(
        \mem[3][11] ), .Z(N21) );
  HS65_LS_MX41X7 U41 ( .D0(n158), .S0(\mem[0][12] ), .D1(n157), .S1(
        \mem[1][12] ), .D2(n156), .S2(\mem[2][12] ), .D3(n155), .S3(
        \mem[3][12] ), .Z(N20) );
  HS65_LS_MX41X7 U42 ( .D0(n158), .S0(\mem[0][13] ), .D1(n157), .S1(
        \mem[1][13] ), .D2(n156), .S2(\mem[2][13] ), .D3(n155), .S3(
        \mem[3][13] ), .Z(N19) );
  HS65_LS_MX41X7 U43 ( .D0(n158), .S0(\mem[0][14] ), .D1(n157), .S1(
        \mem[1][14] ), .D2(n156), .S2(\mem[2][14] ), .D3(n155), .S3(
        \mem[3][14] ), .Z(N18) );
  HS65_LS_MX41X7 U44 ( .D0(n158), .S0(\mem[0][15] ), .D1(n157), .S1(
        \mem[1][15] ), .D2(n156), .S2(\mem[2][15] ), .D3(n155), .S3(
        \mem[3][15] ), .Z(N17) );
  HS65_LS_AO22X9 U45 ( .A(wr_data[0]), .B(n86), .C(n161), .D(\mem[1][0] ), .Z(
        n138) );
  HS65_LS_AO22X9 U46 ( .A(wr_data[1]), .B(n86), .C(n161), .D(\mem[1][1] ), .Z(
        n137) );
  HS65_LS_AO22X9 U47 ( .A(wr_data[2]), .B(n86), .C(n161), .D(\mem[1][2] ), .Z(
        n136) );
  HS65_LS_AO22X9 U48 ( .A(wr_data[3]), .B(n86), .C(n161), .D(\mem[1][3] ), .Z(
        n135) );
  HS65_LS_AO22X9 U49 ( .A(wr_data[4]), .B(n86), .C(n161), .D(\mem[1][4] ), .Z(
        n134) );
  HS65_LS_AO22X9 U50 ( .A(wr_data[5]), .B(n86), .C(n161), .D(\mem[1][5] ), .Z(
        n133) );
  HS65_LS_AO22X9 U51 ( .A(wr_data[6]), .B(n86), .C(n161), .D(\mem[1][6] ), .Z(
        n132) );
  HS65_LS_AO22X9 U52 ( .A(wr_data[7]), .B(n86), .C(n161), .D(\mem[1][7] ), .Z(
        n131) );
  HS65_LS_AO22X9 U53 ( .A(wr_data[8]), .B(n86), .C(n161), .D(\mem[1][8] ), .Z(
        n130) );
  HS65_LS_AO22X9 U54 ( .A(wr_data[9]), .B(n86), .C(n161), .D(\mem[1][9] ), .Z(
        n129) );
  HS65_LS_AO22X9 U55 ( .A(wr_data[10]), .B(n86), .C(n161), .D(\mem[1][10] ), 
        .Z(n128) );
  HS65_LS_AO22X9 U56 ( .A(wr_data[11]), .B(n86), .C(n161), .D(\mem[1][11] ), 
        .Z(n127) );
  HS65_LS_AO22X9 U57 ( .A(wr_data[12]), .B(n86), .C(n161), .D(\mem[1][12] ), 
        .Z(n126) );
  HS65_LS_AO22X9 U58 ( .A(wr_data[13]), .B(n86), .C(n161), .D(\mem[1][13] ), 
        .Z(n125) );
  HS65_LS_AO22X9 U59 ( .A(wr_data[14]), .B(n86), .C(n161), .D(\mem[1][14] ), 
        .Z(n124) );
  HS65_LS_AO22X9 U60 ( .A(wr_data[15]), .B(n86), .C(n161), .D(\mem[1][15] ), 
        .Z(n123) );
  HS65_LS_AO22X9 U61 ( .A(wr_data[0]), .B(n85), .C(n160), .D(\mem[2][0] ), .Z(
        n122) );
  HS65_LS_AO22X9 U62 ( .A(wr_data[1]), .B(n85), .C(n160), .D(\mem[2][1] ), .Z(
        n121) );
  HS65_LS_AO22X9 U63 ( .A(wr_data[2]), .B(n85), .C(n160), .D(\mem[2][2] ), .Z(
        n120) );
  HS65_LS_AO22X9 U64 ( .A(wr_data[3]), .B(n85), .C(n160), .D(\mem[2][3] ), .Z(
        n119) );
  HS65_LS_AO22X9 U65 ( .A(wr_data[4]), .B(n85), .C(n160), .D(\mem[2][4] ), .Z(
        n118) );
  HS65_LS_AO22X9 U66 ( .A(wr_data[5]), .B(n85), .C(n160), .D(\mem[2][5] ), .Z(
        n117) );
  HS65_LS_AO22X9 U67 ( .A(wr_data[6]), .B(n85), .C(n160), .D(\mem[2][6] ), .Z(
        n116) );
  HS65_LS_AO22X9 U68 ( .A(wr_data[7]), .B(n85), .C(n160), .D(\mem[2][7] ), .Z(
        n115) );
  HS65_LS_AO22X9 U69 ( .A(wr_data[8]), .B(n85), .C(n160), .D(\mem[2][8] ), .Z(
        n114) );
  HS65_LS_AO22X9 U70 ( .A(wr_data[9]), .B(n85), .C(n160), .D(\mem[2][9] ), .Z(
        n113) );
  HS65_LS_AO22X9 U71 ( .A(wr_data[10]), .B(n85), .C(n160), .D(\mem[2][10] ), 
        .Z(n112) );
  HS65_LS_AO22X9 U72 ( .A(wr_data[11]), .B(n85), .C(n160), .D(\mem[2][11] ), 
        .Z(n111) );
  HS65_LS_AO22X9 U73 ( .A(wr_data[12]), .B(n85), .C(n160), .D(\mem[2][12] ), 
        .Z(n110) );
  HS65_LS_AO22X9 U74 ( .A(wr_data[13]), .B(n85), .C(n160), .D(\mem[2][13] ), 
        .Z(n109) );
  HS65_LS_AO22X9 U75 ( .A(wr_data[14]), .B(n85), .C(n160), .D(\mem[2][14] ), 
        .Z(n108) );
  HS65_LS_AO22X9 U76 ( .A(wr_data[15]), .B(n85), .C(n160), .D(\mem[2][15] ), 
        .Z(n107) );
  HS65_LS_AO22X9 U77 ( .A(n87), .B(wr_data[0]), .C(n162), .D(\mem[0][0] ), .Z(
        n154) );
  HS65_LS_AO22X9 U78 ( .A(n87), .B(wr_data[1]), .C(n162), .D(\mem[0][1] ), .Z(
        n153) );
  HS65_LS_AO22X9 U79 ( .A(n87), .B(wr_data[2]), .C(n162), .D(\mem[0][2] ), .Z(
        n152) );
  HS65_LS_AO22X9 U80 ( .A(n87), .B(wr_data[3]), .C(n162), .D(\mem[0][3] ), .Z(
        n151) );
  HS65_LS_AO22X9 U81 ( .A(n87), .B(wr_data[4]), .C(n162), .D(\mem[0][4] ), .Z(
        n150) );
  HS65_LS_AO22X9 U82 ( .A(n87), .B(wr_data[5]), .C(n162), .D(\mem[0][5] ), .Z(
        n149) );
  HS65_LS_AO22X9 U83 ( .A(n87), .B(wr_data[6]), .C(n162), .D(\mem[0][6] ), .Z(
        n148) );
  HS65_LS_AO22X9 U84 ( .A(n87), .B(wr_data[7]), .C(n162), .D(\mem[0][7] ), .Z(
        n147) );
  HS65_LS_AO22X9 U85 ( .A(n87), .B(wr_data[8]), .C(n162), .D(\mem[0][8] ), .Z(
        n146) );
  HS65_LS_AO22X9 U86 ( .A(n87), .B(wr_data[9]), .C(n162), .D(\mem[0][9] ), .Z(
        n145) );
  HS65_LS_AO22X9 U87 ( .A(n87), .B(wr_data[10]), .C(n162), .D(\mem[0][10] ), 
        .Z(n144) );
  HS65_LS_AO22X9 U88 ( .A(n87), .B(wr_data[11]), .C(n162), .D(\mem[0][11] ), 
        .Z(n143) );
  HS65_LS_AO22X9 U89 ( .A(n87), .B(wr_data[12]), .C(n162), .D(\mem[0][12] ), 
        .Z(n142) );
  HS65_LS_AO22X9 U90 ( .A(n87), .B(wr_data[13]), .C(n162), .D(\mem[0][13] ), 
        .Z(n141) );
  HS65_LS_AO22X9 U91 ( .A(n87), .B(wr_data[14]), .C(n162), .D(\mem[0][14] ), 
        .Z(n140) );
  HS65_LS_AO22X9 U92 ( .A(n87), .B(wr_data[15]), .C(n162), .D(\mem[0][15] ), 
        .Z(n139) );
  HS65_LS_AO22X9 U93 ( .A(wr_data[0]), .B(n84), .C(n159), .D(\mem[3][0] ), .Z(
        n106) );
  HS65_LS_AO22X9 U94 ( .A(wr_data[1]), .B(n84), .C(n159), .D(\mem[3][1] ), .Z(
        n105) );
  HS65_LS_AO22X9 U95 ( .A(wr_data[2]), .B(n84), .C(n159), .D(\mem[3][2] ), .Z(
        n104) );
  HS65_LS_AO22X9 U96 ( .A(wr_data[3]), .B(n84), .C(n159), .D(\mem[3][3] ), .Z(
        n103) );
  HS65_LS_AO22X9 U97 ( .A(wr_data[4]), .B(n84), .C(n159), .D(\mem[3][4] ), .Z(
        n102) );
  HS65_LS_AO22X9 U98 ( .A(wr_data[5]), .B(n84), .C(n159), .D(\mem[3][5] ), .Z(
        n101) );
  HS65_LS_AO22X9 U99 ( .A(wr_data[6]), .B(n84), .C(n159), .D(\mem[3][6] ), .Z(
        n100) );
  HS65_LS_AO22X9 U100 ( .A(wr_data[7]), .B(n84), .C(n159), .D(\mem[3][7] ), 
        .Z(n99) );
  HS65_LS_AO22X9 U101 ( .A(wr_data[8]), .B(n84), .C(n159), .D(\mem[3][8] ), 
        .Z(n98) );
  HS65_LS_AO22X9 U102 ( .A(wr_data[9]), .B(n84), .C(n159), .D(\mem[3][9] ), 
        .Z(n97) );
  HS65_LS_AO22X9 U103 ( .A(wr_data[10]), .B(n84), .C(n159), .D(\mem[3][10] ), 
        .Z(n96) );
  HS65_LS_AO22X9 U104 ( .A(wr_data[11]), .B(n84), .C(n159), .D(\mem[3][11] ), 
        .Z(n95) );
  HS65_LS_AO22X9 U105 ( .A(wr_data[12]), .B(n84), .C(n159), .D(\mem[3][12] ), 
        .Z(n94) );
  HS65_LS_AO22X9 U106 ( .A(wr_data[13]), .B(n84), .C(n159), .D(\mem[3][13] ), 
        .Z(n93) );
  HS65_LS_AO22X9 U107 ( .A(wr_data[14]), .B(n84), .C(n159), .D(\mem[3][14] ), 
        .Z(n92) );
  HS65_LS_AO22X9 U108 ( .A(wr_data[15]), .B(n84), .C(n159), .D(\mem[3][15] ), 
        .Z(n91) );
endmodule


module bram_DATA32_ADDR2_3 ( clk, reset, rd_addr, wr_addr, wr_data, wr_ena, 
        rd_data );
  input [1:0] rd_addr;
  input [1:0] wr_addr;
  input [31:0] wr_data;
  output [31:0] rd_data;
  input clk, reset, wr_ena;
  wire   \mem[3][31] , \mem[3][30] , \mem[3][29] , \mem[3][28] , \mem[3][27] ,
         \mem[3][26] , \mem[3][25] , \mem[3][24] , \mem[3][23] , \mem[3][22] ,
         \mem[3][21] , \mem[3][20] , \mem[3][19] , \mem[3][18] , \mem[3][17] ,
         \mem[3][16] , \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] ,
         \mem[3][11] , \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] ,
         \mem[3][6] , \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] ,
         \mem[3][1] , \mem[3][0] , \mem[2][31] , \mem[2][30] , \mem[2][29] ,
         \mem[2][28] , \mem[2][27] , \mem[2][26] , \mem[2][25] , \mem[2][24] ,
         \mem[2][23] , \mem[2][22] , \mem[2][21] , \mem[2][20] , \mem[2][19] ,
         \mem[2][18] , \mem[2][17] , \mem[2][16] , \mem[2][15] , \mem[2][14] ,
         \mem[2][13] , \mem[2][12] , \mem[2][11] , \mem[2][10] , \mem[2][9] ,
         \mem[2][8] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][31] ,
         \mem[1][30] , \mem[1][29] , \mem[1][28] , \mem[1][27] , \mem[1][26] ,
         \mem[1][25] , \mem[1][24] , \mem[1][23] , \mem[1][22] , \mem[1][21] ,
         \mem[1][20] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][31] , \mem[0][30] , \mem[0][29] , \mem[0][28] ,
         \mem[0][27] , \mem[0][26] , \mem[0][25] , \mem[0][24] , \mem[0][23] ,
         \mem[0][22] , \mem[0][21] , \mem[0][20] , \mem[0][19] , \mem[0][18] ,
         \mem[0][17] , \mem[0][16] , \mem[0][15] , \mem[0][14] , \mem[0][13] ,
         \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] , \mem[0][8] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N17, N18, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36,
         N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327;

  HS65_LS_DFPRQX9 \mem_reg[3][31]  ( .D(n193), .CP(clk), .RN(n171), .Q(
        \mem[3][31] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][30]  ( .D(n194), .CP(clk), .RN(n171), .Q(
        \mem[3][30] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][29]  ( .D(n195), .CP(clk), .RN(n171), .Q(
        \mem[3][29] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][28]  ( .D(n196), .CP(clk), .RN(n171), .Q(
        \mem[3][28] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][27]  ( .D(n197), .CP(clk), .RN(n171), .Q(
        \mem[3][27] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][26]  ( .D(n198), .CP(clk), .RN(n171), .Q(
        \mem[3][26] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][25]  ( .D(n199), .CP(clk), .RN(n171), .Q(
        \mem[3][25] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][24]  ( .D(n200), .CP(clk), .RN(n171), .Q(
        \mem[3][24] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][23]  ( .D(n201), .CP(clk), .RN(n171), .Q(
        \mem[3][23] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][22]  ( .D(n202), .CP(clk), .RN(n171), .Q(
        \mem[3][22] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][21]  ( .D(n203), .CP(clk), .RN(n171), .Q(
        \mem[3][21] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][20]  ( .D(n204), .CP(clk), .RN(n171), .Q(
        \mem[3][20] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][19]  ( .D(n205), .CP(clk), .RN(n171), .Q(
        \mem[3][19] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][18]  ( .D(n206), .CP(clk), .RN(n172), .Q(
        \mem[3][18] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][17]  ( .D(n207), .CP(clk), .RN(n172), .Q(
        \mem[3][17] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][16]  ( .D(n208), .CP(clk), .RN(n172), .Q(
        \mem[3][16] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][15]  ( .D(n209), .CP(clk), .RN(n172), .Q(
        \mem[3][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][14]  ( .D(n210), .CP(clk), .RN(n172), .Q(
        \mem[3][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][13]  ( .D(n211), .CP(clk), .RN(n172), .Q(
        \mem[3][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][12]  ( .D(n212), .CP(clk), .RN(n172), .Q(
        \mem[3][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][11]  ( .D(n213), .CP(clk), .RN(n172), .Q(
        \mem[3][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][10]  ( .D(n214), .CP(clk), .RN(n172), .Q(
        \mem[3][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][9]  ( .D(n215), .CP(clk), .RN(n172), .Q(
        \mem[3][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][8]  ( .D(n216), .CP(clk), .RN(n172), .Q(
        \mem[3][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][7]  ( .D(n217), .CP(clk), .RN(n172), .Q(
        \mem[3][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][6]  ( .D(n218), .CP(clk), .RN(n172), .Q(
        \mem[3][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][5]  ( .D(n219), .CP(clk), .RN(n173), .Q(
        \mem[3][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][4]  ( .D(n220), .CP(clk), .RN(n173), .Q(
        \mem[3][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][3]  ( .D(n221), .CP(clk), .RN(n173), .Q(
        \mem[3][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][2]  ( .D(n222), .CP(clk), .RN(n173), .Q(
        \mem[3][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][1]  ( .D(n223), .CP(clk), .RN(n173), .Q(
        \mem[3][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][0]  ( .D(n224), .CP(clk), .RN(n173), .Q(
        \mem[3][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][31]  ( .D(n225), .CP(clk), .RN(n173), .Q(
        \mem[2][31] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][30]  ( .D(n226), .CP(clk), .RN(n173), .Q(
        \mem[2][30] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][29]  ( .D(n227), .CP(clk), .RN(n173), .Q(
        \mem[2][29] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][28]  ( .D(n228), .CP(clk), .RN(n173), .Q(
        \mem[2][28] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][27]  ( .D(n229), .CP(clk), .RN(n173), .Q(
        \mem[2][27] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][26]  ( .D(n230), .CP(clk), .RN(n173), .Q(
        \mem[2][26] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][25]  ( .D(n231), .CP(clk), .RN(n173), .Q(
        \mem[2][25] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][24]  ( .D(n232), .CP(clk), .RN(n174), .Q(
        \mem[2][24] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][23]  ( .D(n233), .CP(clk), .RN(n174), .Q(
        \mem[2][23] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][22]  ( .D(n234), .CP(clk), .RN(n174), .Q(
        \mem[2][22] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][21]  ( .D(n235), .CP(clk), .RN(n174), .Q(
        \mem[2][21] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][20]  ( .D(n236), .CP(clk), .RN(n174), .Q(
        \mem[2][20] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][19]  ( .D(n237), .CP(clk), .RN(n174), .Q(
        \mem[2][19] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][18]  ( .D(n238), .CP(clk), .RN(n174), .Q(
        \mem[2][18] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][17]  ( .D(n239), .CP(clk), .RN(n174), .Q(
        \mem[2][17] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][16]  ( .D(n240), .CP(clk), .RN(n174), .Q(
        \mem[2][16] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][15]  ( .D(n241), .CP(clk), .RN(n174), .Q(
        \mem[2][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][14]  ( .D(n242), .CP(clk), .RN(n174), .Q(
        \mem[2][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][13]  ( .D(n243), .CP(clk), .RN(n174), .Q(
        \mem[2][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][12]  ( .D(n244), .CP(clk), .RN(n174), .Q(
        \mem[2][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][11]  ( .D(n245), .CP(clk), .RN(n175), .Q(
        \mem[2][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][10]  ( .D(n246), .CP(clk), .RN(n175), .Q(
        \mem[2][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][9]  ( .D(n247), .CP(clk), .RN(n175), .Q(
        \mem[2][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][8]  ( .D(n248), .CP(clk), .RN(n175), .Q(
        \mem[2][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][7]  ( .D(n249), .CP(clk), .RN(n175), .Q(
        \mem[2][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][6]  ( .D(n250), .CP(clk), .RN(n175), .Q(
        \mem[2][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][5]  ( .D(n251), .CP(clk), .RN(n175), .Q(
        \mem[2][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][4]  ( .D(n252), .CP(clk), .RN(n175), .Q(
        \mem[2][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][3]  ( .D(n253), .CP(clk), .RN(n175), .Q(
        \mem[2][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][2]  ( .D(n254), .CP(clk), .RN(n175), .Q(
        \mem[2][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][1]  ( .D(n255), .CP(clk), .RN(n175), .Q(
        \mem[2][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][0]  ( .D(n256), .CP(clk), .RN(n175), .Q(
        \mem[2][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][31]  ( .D(n257), .CP(clk), .RN(n175), .Q(
        \mem[1][31] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][30]  ( .D(n258), .CP(clk), .RN(n176), .Q(
        \mem[1][30] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][29]  ( .D(n259), .CP(clk), .RN(n176), .Q(
        \mem[1][29] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][28]  ( .D(n260), .CP(clk), .RN(n176), .Q(
        \mem[1][28] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][27]  ( .D(n261), .CP(clk), .RN(n176), .Q(
        \mem[1][27] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][26]  ( .D(n262), .CP(clk), .RN(n176), .Q(
        \mem[1][26] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][25]  ( .D(n263), .CP(clk), .RN(n176), .Q(
        \mem[1][25] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][24]  ( .D(n264), .CP(clk), .RN(n176), .Q(
        \mem[1][24] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][23]  ( .D(n265), .CP(clk), .RN(n176), .Q(
        \mem[1][23] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][22]  ( .D(n266), .CP(clk), .RN(n176), .Q(
        \mem[1][22] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][21]  ( .D(n267), .CP(clk), .RN(n176), .Q(
        \mem[1][21] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][20]  ( .D(n268), .CP(clk), .RN(n176), .Q(
        \mem[1][20] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][19]  ( .D(n269), .CP(clk), .RN(n176), .Q(
        \mem[1][19] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][18]  ( .D(n270), .CP(clk), .RN(n176), .Q(
        \mem[1][18] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][17]  ( .D(n271), .CP(clk), .RN(n177), .Q(
        \mem[1][17] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][16]  ( .D(n272), .CP(clk), .RN(n177), .Q(
        \mem[1][16] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][15]  ( .D(n273), .CP(clk), .RN(n177), .Q(
        \mem[1][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][14]  ( .D(n274), .CP(clk), .RN(n177), .Q(
        \mem[1][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][13]  ( .D(n275), .CP(clk), .RN(n177), .Q(
        \mem[1][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][12]  ( .D(n276), .CP(clk), .RN(n177), .Q(
        \mem[1][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][11]  ( .D(n277), .CP(clk), .RN(n177), .Q(
        \mem[1][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][10]  ( .D(n278), .CP(clk), .RN(n177), .Q(
        \mem[1][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][9]  ( .D(n279), .CP(clk), .RN(n177), .Q(
        \mem[1][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][8]  ( .D(n280), .CP(clk), .RN(n177), .Q(
        \mem[1][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][7]  ( .D(n281), .CP(clk), .RN(n177), .Q(
        \mem[1][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][6]  ( .D(n282), .CP(clk), .RN(n177), .Q(
        \mem[1][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][5]  ( .D(n283), .CP(clk), .RN(n177), .Q(
        \mem[1][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][4]  ( .D(n284), .CP(clk), .RN(n178), .Q(
        \mem[1][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][3]  ( .D(n285), .CP(clk), .RN(n178), .Q(
        \mem[1][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][2]  ( .D(n286), .CP(clk), .RN(n178), .Q(
        \mem[1][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][1]  ( .D(n287), .CP(clk), .RN(n178), .Q(
        \mem[1][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][0]  ( .D(n288), .CP(clk), .RN(n178), .Q(
        \mem[1][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][31]  ( .D(n289), .CP(clk), .RN(n178), .Q(
        \mem[0][31] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][30]  ( .D(n290), .CP(clk), .RN(n178), .Q(
        \mem[0][30] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][29]  ( .D(n291), .CP(clk), .RN(n178), .Q(
        \mem[0][29] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][28]  ( .D(n292), .CP(clk), .RN(n178), .Q(
        \mem[0][28] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][27]  ( .D(n293), .CP(clk), .RN(n178), .Q(
        \mem[0][27] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][26]  ( .D(n294), .CP(clk), .RN(n178), .Q(
        \mem[0][26] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][25]  ( .D(n295), .CP(clk), .RN(n178), .Q(
        \mem[0][25] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][24]  ( .D(n296), .CP(clk), .RN(n178), .Q(
        \mem[0][24] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][23]  ( .D(n297), .CP(clk), .RN(n179), .Q(
        \mem[0][23] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][22]  ( .D(n298), .CP(clk), .RN(n179), .Q(
        \mem[0][22] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][21]  ( .D(n299), .CP(clk), .RN(n179), .Q(
        \mem[0][21] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][20]  ( .D(n300), .CP(clk), .RN(n179), .Q(
        \mem[0][20] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][19]  ( .D(n301), .CP(clk), .RN(n179), .Q(
        \mem[0][19] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][18]  ( .D(n302), .CP(clk), .RN(n179), .Q(
        \mem[0][18] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][17]  ( .D(n303), .CP(clk), .RN(n179), .Q(
        \mem[0][17] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][16]  ( .D(n304), .CP(clk), .RN(n179), .Q(
        \mem[0][16] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][15]  ( .D(n305), .CP(clk), .RN(n179), .Q(
        \mem[0][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][14]  ( .D(n306), .CP(clk), .RN(n179), .Q(
        \mem[0][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][13]  ( .D(n307), .CP(clk), .RN(n179), .Q(
        \mem[0][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][12]  ( .D(n308), .CP(clk), .RN(n179), .Q(
        \mem[0][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][11]  ( .D(n309), .CP(clk), .RN(n179), .Q(
        \mem[0][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][10]  ( .D(n310), .CP(clk), .RN(n180), .Q(
        \mem[0][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][9]  ( .D(n311), .CP(clk), .RN(n180), .Q(
        \mem[0][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][8]  ( .D(n312), .CP(clk), .RN(n180), .Q(
        \mem[0][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][7]  ( .D(n313), .CP(clk), .RN(n180), .Q(
        \mem[0][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][6]  ( .D(n314), .CP(clk), .RN(n180), .Q(
        \mem[0][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][5]  ( .D(n315), .CP(clk), .RN(n180), .Q(
        \mem[0][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][4]  ( .D(n316), .CP(clk), .RN(n180), .Q(
        \mem[0][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][3]  ( .D(n317), .CP(clk), .RN(n180), .Q(
        \mem[0][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][2]  ( .D(n318), .CP(clk), .RN(n180), .Q(
        \mem[0][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][1]  ( .D(n319), .CP(clk), .RN(n180), .Q(
        \mem[0][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][0]  ( .D(n320), .CP(clk), .RN(n180), .Q(
        \mem[0][0] ) );
  HS65_LS_DFPRQX9 \rd_data_reg[31]  ( .D(N17), .CP(clk), .RN(n180), .Q(
        rd_data[31]) );
  HS65_LS_DFPRQX9 \rd_data_reg[30]  ( .D(N18), .CP(clk), .RN(n180), .Q(
        rd_data[30]) );
  HS65_LS_DFPRQX9 \rd_data_reg[29]  ( .D(N19), .CP(clk), .RN(n181), .Q(
        rd_data[29]) );
  HS65_LS_DFPRQX9 \rd_data_reg[28]  ( .D(N20), .CP(clk), .RN(n181), .Q(
        rd_data[28]) );
  HS65_LS_DFPRQX9 \rd_data_reg[27]  ( .D(N21), .CP(clk), .RN(n181), .Q(
        rd_data[27]) );
  HS65_LS_DFPRQX9 \rd_data_reg[26]  ( .D(N22), .CP(clk), .RN(n181), .Q(
        rd_data[26]) );
  HS65_LS_DFPRQX9 \rd_data_reg[25]  ( .D(N23), .CP(clk), .RN(n181), .Q(
        rd_data[25]) );
  HS65_LS_DFPRQX9 \rd_data_reg[24]  ( .D(N24), .CP(clk), .RN(n181), .Q(
        rd_data[24]) );
  HS65_LS_DFPRQX9 \rd_data_reg[23]  ( .D(N25), .CP(clk), .RN(n181), .Q(
        rd_data[23]) );
  HS65_LS_DFPRQX9 \rd_data_reg[22]  ( .D(N26), .CP(clk), .RN(n181), .Q(
        rd_data[22]) );
  HS65_LS_DFPRQX9 \rd_data_reg[21]  ( .D(N27), .CP(clk), .RN(n181), .Q(
        rd_data[21]) );
  HS65_LS_DFPRQX9 \rd_data_reg[20]  ( .D(N28), .CP(clk), .RN(n181), .Q(
        rd_data[20]) );
  HS65_LS_DFPRQX9 \rd_data_reg[19]  ( .D(N29), .CP(clk), .RN(n181), .Q(
        rd_data[19]) );
  HS65_LS_DFPRQX9 \rd_data_reg[18]  ( .D(N30), .CP(clk), .RN(n181), .Q(
        rd_data[18]) );
  HS65_LS_DFPRQX9 \rd_data_reg[17]  ( .D(N31), .CP(clk), .RN(n181), .Q(
        rd_data[17]) );
  HS65_LS_DFPRQX9 \rd_data_reg[16]  ( .D(N32), .CP(clk), .RN(n182), .Q(
        rd_data[16]) );
  HS65_LS_DFPRQX9 \rd_data_reg[15]  ( .D(N33), .CP(clk), .RN(n182), .Q(
        rd_data[15]) );
  HS65_LS_DFPRQX9 \rd_data_reg[14]  ( .D(N34), .CP(clk), .RN(n182), .Q(
        rd_data[14]) );
  HS65_LS_DFPRQX9 \rd_data_reg[13]  ( .D(N35), .CP(clk), .RN(n182), .Q(
        rd_data[13]) );
  HS65_LS_DFPRQX9 \rd_data_reg[12]  ( .D(N36), .CP(clk), .RN(n182), .Q(
        rd_data[12]) );
  HS65_LS_DFPRQX9 \rd_data_reg[11]  ( .D(N37), .CP(clk), .RN(n182), .Q(
        rd_data[11]) );
  HS65_LS_DFPRQX9 \rd_data_reg[10]  ( .D(N38), .CP(clk), .RN(n182), .Q(
        rd_data[10]) );
  HS65_LS_DFPRQX9 \rd_data_reg[9]  ( .D(N39), .CP(clk), .RN(n182), .Q(
        rd_data[9]) );
  HS65_LS_DFPRQX9 \rd_data_reg[8]  ( .D(N40), .CP(clk), .RN(n182), .Q(
        rd_data[8]) );
  HS65_LS_DFPRQX9 \rd_data_reg[7]  ( .D(N41), .CP(clk), .RN(n182), .Q(
        rd_data[7]) );
  HS65_LS_DFPRQX9 \rd_data_reg[6]  ( .D(N42), .CP(clk), .RN(n182), .Q(
        rd_data[6]) );
  HS65_LS_DFPRQX9 \rd_data_reg[5]  ( .D(N43), .CP(clk), .RN(n182), .Q(
        rd_data[5]) );
  HS65_LS_DFPRQX9 \rd_data_reg[4]  ( .D(N44), .CP(clk), .RN(n182), .Q(
        rd_data[4]) );
  HS65_LS_DFPRQX9 \rd_data_reg[3]  ( .D(N45), .CP(clk), .RN(n183), .Q(
        rd_data[3]) );
  HS65_LS_DFPRQX9 \rd_data_reg[2]  ( .D(N46), .CP(clk), .RN(n183), .Q(
        rd_data[2]) );
  HS65_LS_DFPRQX9 \rd_data_reg[1]  ( .D(N47), .CP(clk), .RN(n183), .Q(
        rd_data[1]) );
  HS65_LS_DFPRQX9 \rd_data_reg[0]  ( .D(N48), .CP(clk), .RN(n183), .Q(
        rd_data[0]) );
  HS65_LS_AND3X9 U3 ( .A(n191), .B(n190), .C(wr_ena), .Z(n1) );
  HS65_LS_BFX9 U4 ( .A(n165), .Z(n162) );
  HS65_LS_BFX9 U5 ( .A(n1), .Z(n168) );
  HS65_LS_BFX9 U6 ( .A(n160), .Z(n157) );
  HS65_LS_BFX9 U7 ( .A(n155), .Z(n152) );
  HS65_LS_AND2X4 U8 ( .A(rd_addr[1]), .B(rd_addr[0]), .Z(n321) );
  HS65_LS_AND2X4 U9 ( .A(rd_addr[1]), .B(n192), .Z(n322) );
  HS65_LS_BFX9 U10 ( .A(n185), .Z(n180) );
  HS65_LS_BFX9 U11 ( .A(n185), .Z(n179) );
  HS65_LS_BFX9 U12 ( .A(n185), .Z(n178) );
  HS65_LS_BFX9 U13 ( .A(n186), .Z(n177) );
  HS65_LS_BFX9 U14 ( .A(n186), .Z(n176) );
  HS65_LS_BFX9 U15 ( .A(n186), .Z(n175) );
  HS65_LS_BFX9 U16 ( .A(n187), .Z(n174) );
  HS65_LS_BFX9 U17 ( .A(n187), .Z(n173) );
  HS65_LS_BFX9 U18 ( .A(n187), .Z(n172) );
  HS65_LS_BFX9 U19 ( .A(n188), .Z(n185) );
  HS65_LS_BFX9 U20 ( .A(n188), .Z(n186) );
  HS65_LS_BFX9 U21 ( .A(n189), .Z(n187) );
  HS65_LS_BFX9 U22 ( .A(n184), .Z(n182) );
  HS65_LS_BFX9 U23 ( .A(n184), .Z(n181) );
  HS65_LS_BFX9 U24 ( .A(n188), .Z(n171) );
  HS65_LS_BFX9 U25 ( .A(n189), .Z(n188) );
  HS65_LS_BFX9 U26 ( .A(n184), .Z(n183) );
  HS65_LS_BFX9 U27 ( .A(n189), .Z(n184) );
  HS65_LS_IVX9 U28 ( .A(reset), .Z(n189) );
  HS65_LS_IVX9 U29 ( .A(n168), .Z(n167) );
  HS65_LS_IVX9 U30 ( .A(n168), .Z(n166) );
  HS65_LS_IVX9 U31 ( .A(n162), .Z(n161) );
  HS65_LS_BFX9 U32 ( .A(n1), .Z(n169) );
  HS65_LS_BFX9 U33 ( .A(n165), .Z(n163) );
  HS65_LS_BFX9 U34 ( .A(n1), .Z(n170) );
  HS65_LS_BFX9 U35 ( .A(n162), .Z(n164) );
  HS65_LS_IVX9 U36 ( .A(n157), .Z(n156) );
  HS65_LS_IVX9 U37 ( .A(n152), .Z(n151) );
  HS65_LS_BFX9 U38 ( .A(n160), .Z(n158) );
  HS65_LS_BFX9 U39 ( .A(n155), .Z(n153) );
  HS65_LS_BFX9 U40 ( .A(n157), .Z(n159) );
  HS65_LS_BFX9 U41 ( .A(n152), .Z(n154) );
  HS65_LS_IVX9 U42 ( .A(n327), .Z(n165) );
  HS65_LS_IVX9 U43 ( .A(wr_addr[0]), .Z(n191) );
  HS65_LS_NAND3X5 U44 ( .A(wr_ena), .B(n190), .C(wr_addr[0]), .Z(n327) );
  HS65_LS_BFX9 U45 ( .A(n322), .Z(n6) );
  HS65_LS_BFX9 U46 ( .A(n322), .Z(n5) );
  HS65_LS_BFX9 U47 ( .A(n321), .Z(n3) );
  HS65_LS_BFX9 U48 ( .A(n321), .Z(n2) );
  HS65_LS_BFX9 U49 ( .A(n8), .Z(n145) );
  HS65_LS_BFX9 U50 ( .A(n8), .Z(n9) );
  HS65_LS_BFX9 U51 ( .A(n147), .Z(n149) );
  HS65_LS_BFX9 U52 ( .A(n147), .Z(n148) );
  HS65_LS_BFX9 U53 ( .A(n321), .Z(n4) );
  HS65_LS_BFX9 U54 ( .A(n322), .Z(n7) );
  HS65_LS_BFX9 U55 ( .A(n8), .Z(n146) );
  HS65_LS_BFX9 U56 ( .A(n147), .Z(n150) );
  HS65_LS_IVX9 U57 ( .A(n326), .Z(n160) );
  HS65_LS_IVX9 U58 ( .A(n325), .Z(n155) );
  HS65_LS_IVX9 U59 ( .A(wr_addr[1]), .Z(n190) );
  HS65_LS_IVX9 U60 ( .A(rd_addr[0]), .Z(n192) );
  HS65_LS_NAND3X5 U61 ( .A(wr_addr[0]), .B(wr_ena), .C(wr_addr[1]), .Z(n325)
         );
  HS65_LS_NAND3X5 U62 ( .A(wr_ena), .B(n191), .C(wr_addr[1]), .Z(n326) );
  HS65_LS_BFX9 U63 ( .A(n324), .Z(n147) );
  HS65_LS_NOR2X6 U64 ( .A(rd_addr[0]), .B(rd_addr[1]), .Z(n324) );
  HS65_LS_BFX9 U65 ( .A(n323), .Z(n8) );
  HS65_LH_NOR2X2 U66 ( .A(n192), .B(rd_addr[1]), .Z(n323) );
  HS65_LS_MX41X7 U67 ( .D0(n150), .S0(\mem[0][0] ), .D1(n146), .S1(\mem[1][0] ), .D2(n7), .S2(\mem[2][0] ), .D3(n4), .S3(\mem[3][0] ), .Z(N48) );
  HS65_LS_MX41X7 U68 ( .D0(n150), .S0(\mem[0][1] ), .D1(n146), .S1(\mem[1][1] ), .D2(n7), .S2(\mem[2][1] ), .D3(n4), .S3(\mem[3][1] ), .Z(N47) );
  HS65_LS_MX41X7 U69 ( .D0(n150), .S0(\mem[0][2] ), .D1(n146), .S1(\mem[1][2] ), .D2(n7), .S2(\mem[2][2] ), .D3(n4), .S3(\mem[3][2] ), .Z(N46) );
  HS65_LS_MX41X7 U70 ( .D0(n150), .S0(\mem[0][3] ), .D1(n146), .S1(\mem[1][3] ), .D2(n7), .S2(\mem[2][3] ), .D3(n4), .S3(\mem[3][3] ), .Z(N45) );
  HS65_LS_MX41X7 U71 ( .D0(n150), .S0(\mem[0][4] ), .D1(n146), .S1(\mem[1][4] ), .D2(n7), .S2(\mem[2][4] ), .D3(n4), .S3(\mem[3][4] ), .Z(N44) );
  HS65_LS_MX41X7 U72 ( .D0(n150), .S0(\mem[0][5] ), .D1(n146), .S1(\mem[1][5] ), .D2(n7), .S2(\mem[2][5] ), .D3(n4), .S3(\mem[3][5] ), .Z(N43) );
  HS65_LS_MX41X7 U73 ( .D0(n150), .S0(\mem[0][6] ), .D1(n146), .S1(\mem[1][6] ), .D2(n6), .S2(\mem[2][6] ), .D3(n4), .S3(\mem[3][6] ), .Z(N42) );
  HS65_LS_MX41X7 U74 ( .D0(n150), .S0(\mem[0][7] ), .D1(n146), .S1(\mem[1][7] ), .D2(n6), .S2(\mem[2][7] ), .D3(n4), .S3(\mem[3][7] ), .Z(N41) );
  HS65_LS_MX41X7 U75 ( .D0(n149), .S0(\mem[0][8] ), .D1(n145), .S1(\mem[1][8] ), .D2(n6), .S2(\mem[2][8] ), .D3(n3), .S3(\mem[3][8] ), .Z(N40) );
  HS65_LS_MX41X7 U76 ( .D0(n149), .S0(\mem[0][9] ), .D1(n145), .S1(\mem[1][9] ), .D2(n6), .S2(\mem[2][9] ), .D3(n3), .S3(\mem[3][9] ), .Z(N39) );
  HS65_LS_MX41X7 U77 ( .D0(n149), .S0(\mem[0][10] ), .D1(n145), .S1(
        \mem[1][10] ), .D2(n6), .S2(\mem[2][10] ), .D3(n3), .S3(\mem[3][10] ), 
        .Z(N38) );
  HS65_LS_MX41X7 U78 ( .D0(n149), .S0(\mem[0][11] ), .D1(n145), .S1(
        \mem[1][11] ), .D2(n6), .S2(\mem[2][11] ), .D3(n3), .S3(\mem[3][11] ), 
        .Z(N37) );
  HS65_LS_MX41X7 U79 ( .D0(n149), .S0(\mem[0][12] ), .D1(n145), .S1(
        \mem[1][12] ), .D2(n6), .S2(\mem[2][12] ), .D3(n3), .S3(\mem[3][12] ), 
        .Z(N36) );
  HS65_LS_MX41X7 U80 ( .D0(n149), .S0(\mem[0][13] ), .D1(n145), .S1(
        \mem[1][13] ), .D2(n6), .S2(\mem[2][13] ), .D3(n3), .S3(\mem[3][13] ), 
        .Z(N35) );
  HS65_LS_MX41X7 U81 ( .D0(n149), .S0(\mem[0][14] ), .D1(n145), .S1(
        \mem[1][14] ), .D2(n6), .S2(\mem[2][14] ), .D3(n3), .S3(\mem[3][14] ), 
        .Z(N34) );
  HS65_LS_MX41X7 U82 ( .D0(n149), .S0(\mem[0][15] ), .D1(n145), .S1(
        \mem[1][15] ), .D2(n6), .S2(\mem[2][15] ), .D3(n3), .S3(\mem[3][15] ), 
        .Z(N33) );
  HS65_LS_MX41X7 U83 ( .D0(n149), .S0(\mem[0][16] ), .D1(n145), .S1(
        \mem[1][16] ), .D2(n6), .S2(\mem[2][16] ), .D3(n3), .S3(\mem[3][16] ), 
        .Z(N32) );
  HS65_LS_MX41X7 U84 ( .D0(n149), .S0(\mem[0][17] ), .D1(n145), .S1(
        \mem[1][17] ), .D2(n6), .S2(\mem[2][17] ), .D3(n3), .S3(\mem[3][17] ), 
        .Z(N31) );
  HS65_LS_MX41X7 U85 ( .D0(n149), .S0(\mem[0][18] ), .D1(n145), .S1(
        \mem[1][18] ), .D2(n6), .S2(\mem[2][18] ), .D3(n3), .S3(\mem[3][18] ), 
        .Z(N30) );
  HS65_LS_MX41X7 U86 ( .D0(n149), .S0(\mem[0][19] ), .D1(n145), .S1(
        \mem[1][19] ), .D2(n5), .S2(\mem[2][19] ), .D3(n3), .S3(\mem[3][19] ), 
        .Z(N29) );
  HS65_LS_MX41X7 U87 ( .D0(n148), .S0(\mem[0][20] ), .D1(n9), .S1(\mem[1][20] ), .D2(n5), .S2(\mem[2][20] ), .D3(n2), .S3(\mem[3][20] ), .Z(N28) );
  HS65_LS_MX41X7 U88 ( .D0(n148), .S0(\mem[0][21] ), .D1(n9), .S1(\mem[1][21] ), .D2(n5), .S2(\mem[2][21] ), .D3(n2), .S3(\mem[3][21] ), .Z(N27) );
  HS65_LS_MX41X7 U89 ( .D0(n148), .S0(\mem[0][22] ), .D1(n9), .S1(\mem[1][22] ), .D2(n5), .S2(\mem[2][22] ), .D3(n2), .S3(\mem[3][22] ), .Z(N26) );
  HS65_LS_MX41X7 U90 ( .D0(n148), .S0(\mem[0][23] ), .D1(n9), .S1(\mem[1][23] ), .D2(n5), .S2(\mem[2][23] ), .D3(n2), .S3(\mem[3][23] ), .Z(N25) );
  HS65_LS_MX41X7 U91 ( .D0(n148), .S0(\mem[0][24] ), .D1(n9), .S1(\mem[1][24] ), .D2(n5), .S2(\mem[2][24] ), .D3(n2), .S3(\mem[3][24] ), .Z(N24) );
  HS65_LS_MX41X7 U92 ( .D0(n148), .S0(\mem[0][25] ), .D1(n9), .S1(\mem[1][25] ), .D2(n5), .S2(\mem[2][25] ), .D3(n2), .S3(\mem[3][25] ), .Z(N23) );
  HS65_LS_MX41X7 U93 ( .D0(n148), .S0(\mem[0][26] ), .D1(n9), .S1(\mem[1][26] ), .D2(n5), .S2(\mem[2][26] ), .D3(n2), .S3(\mem[3][26] ), .Z(N22) );
  HS65_LS_MX41X7 U94 ( .D0(n148), .S0(\mem[0][27] ), .D1(n9), .S1(\mem[1][27] ), .D2(n5), .S2(\mem[2][27] ), .D3(n2), .S3(\mem[3][27] ), .Z(N21) );
  HS65_LS_MX41X7 U95 ( .D0(n148), .S0(\mem[0][28] ), .D1(n9), .S1(\mem[1][28] ), .D2(n5), .S2(\mem[2][28] ), .D3(n2), .S3(\mem[3][28] ), .Z(N20) );
  HS65_LS_MX41X7 U96 ( .D0(n148), .S0(\mem[0][29] ), .D1(n9), .S1(\mem[1][29] ), .D2(n5), .S2(\mem[2][29] ), .D3(n2), .S3(\mem[3][29] ), .Z(N19) );
  HS65_LS_MX41X7 U97 ( .D0(n148), .S0(\mem[0][30] ), .D1(n9), .S1(\mem[1][30] ), .D2(n5), .S2(\mem[2][30] ), .D3(n2), .S3(\mem[3][30] ), .Z(N18) );
  HS65_LS_MX41X7 U98 ( .D0(n148), .S0(\mem[0][31] ), .D1(n9), .S1(\mem[1][31] ), .D2(n5), .S2(\mem[2][31] ), .D3(n2), .S3(\mem[3][31] ), .Z(N17) );
  HS65_LS_AO22X9 U99 ( .A(wr_data[0]), .B(n154), .C(n151), .D(\mem[3][0] ), 
        .Z(n224) );
  HS65_LS_AO22X9 U100 ( .A(wr_data[1]), .B(n154), .C(n151), .D(\mem[3][1] ), 
        .Z(n223) );
  HS65_LS_AO22X9 U101 ( .A(wr_data[2]), .B(n154), .C(n151), .D(\mem[3][2] ), 
        .Z(n222) );
  HS65_LS_AO22X9 U102 ( .A(wr_data[3]), .B(n154), .C(n151), .D(\mem[3][3] ), 
        .Z(n221) );
  HS65_LS_AO22X9 U103 ( .A(wr_data[4]), .B(n154), .C(n151), .D(\mem[3][4] ), 
        .Z(n220) );
  HS65_LS_AO22X9 U104 ( .A(wr_data[5]), .B(n154), .C(n151), .D(\mem[3][5] ), 
        .Z(n219) );
  HS65_LS_AO22X9 U105 ( .A(wr_data[6]), .B(n154), .C(n151), .D(\mem[3][6] ), 
        .Z(n218) );
  HS65_LS_AO22X9 U106 ( .A(wr_data[7]), .B(n154), .C(n151), .D(\mem[3][7] ), 
        .Z(n217) );
  HS65_LS_AO22X9 U107 ( .A(wr_data[8]), .B(n154), .C(n151), .D(\mem[3][8] ), 
        .Z(n216) );
  HS65_LS_AO22X9 U108 ( .A(wr_data[9]), .B(n154), .C(n151), .D(\mem[3][9] ), 
        .Z(n215) );
  HS65_LS_AO22X9 U109 ( .A(wr_data[10]), .B(n154), .C(n151), .D(\mem[3][10] ), 
        .Z(n214) );
  HS65_LS_AO22X9 U110 ( .A(wr_data[11]), .B(n153), .C(n151), .D(\mem[3][11] ), 
        .Z(n213) );
  HS65_LS_AO22X9 U111 ( .A(wr_data[12]), .B(n153), .C(n151), .D(\mem[3][12] ), 
        .Z(n212) );
  HS65_LS_AO22X9 U112 ( .A(wr_data[13]), .B(n153), .C(n151), .D(\mem[3][13] ), 
        .Z(n211) );
  HS65_LS_AO22X9 U113 ( .A(wr_data[14]), .B(n153), .C(n151), .D(\mem[3][14] ), 
        .Z(n210) );
  HS65_LS_AO22X9 U114 ( .A(wr_data[15]), .B(n153), .C(n151), .D(\mem[3][15] ), 
        .Z(n209) );
  HS65_LS_AO22X9 U115 ( .A(wr_data[16]), .B(n153), .C(n151), .D(\mem[3][16] ), 
        .Z(n208) );
  HS65_LS_AO22X9 U116 ( .A(wr_data[17]), .B(n153), .C(n151), .D(\mem[3][17] ), 
        .Z(n207) );
  HS65_LS_AO22X9 U117 ( .A(wr_data[18]), .B(n153), .C(n151), .D(\mem[3][18] ), 
        .Z(n206) );
  HS65_LS_AO22X9 U118 ( .A(wr_data[19]), .B(n153), .C(n151), .D(\mem[3][19] ), 
        .Z(n205) );
  HS65_LS_AO22X9 U119 ( .A(wr_data[20]), .B(n153), .C(n325), .D(\mem[3][20] ), 
        .Z(n204) );
  HS65_LS_AO22X9 U120 ( .A(wr_data[21]), .B(n153), .C(n325), .D(\mem[3][21] ), 
        .Z(n203) );
  HS65_LS_AO22X9 U121 ( .A(wr_data[22]), .B(n153), .C(n325), .D(\mem[3][22] ), 
        .Z(n202) );
  HS65_LS_AO22X9 U122 ( .A(wr_data[23]), .B(n153), .C(n325), .D(\mem[3][23] ), 
        .Z(n201) );
  HS65_LS_AO22X9 U123 ( .A(wr_data[24]), .B(n153), .C(n325), .D(\mem[3][24] ), 
        .Z(n200) );
  HS65_LS_AO22X9 U124 ( .A(wr_data[25]), .B(n153), .C(n325), .D(\mem[3][25] ), 
        .Z(n199) );
  HS65_LS_AO22X9 U125 ( .A(wr_data[26]), .B(n153), .C(n325), .D(\mem[3][26] ), 
        .Z(n198) );
  HS65_LS_AO22X9 U126 ( .A(wr_data[27]), .B(n153), .C(n325), .D(\mem[3][27] ), 
        .Z(n197) );
  HS65_LS_AO22X9 U127 ( .A(wr_data[28]), .B(n153), .C(n325), .D(\mem[3][28] ), 
        .Z(n196) );
  HS65_LS_AO22X9 U128 ( .A(wr_data[29]), .B(n153), .C(n325), .D(\mem[3][29] ), 
        .Z(n195) );
  HS65_LS_AO22X9 U129 ( .A(wr_data[30]), .B(n153), .C(n325), .D(\mem[3][30] ), 
        .Z(n194) );
  HS65_LS_AO22X9 U130 ( .A(wr_data[31]), .B(n152), .C(n325), .D(\mem[3][31] ), 
        .Z(n193) );
  HS65_LS_AO22X9 U131 ( .A(wr_data[0]), .B(n164), .C(n161), .D(\mem[1][0] ), 
        .Z(n288) );
  HS65_LS_AO22X9 U132 ( .A(wr_data[1]), .B(n164), .C(n161), .D(\mem[1][1] ), 
        .Z(n287) );
  HS65_LS_AO22X9 U133 ( .A(wr_data[2]), .B(n164), .C(n161), .D(\mem[1][2] ), 
        .Z(n286) );
  HS65_LS_AO22X9 U134 ( .A(wr_data[3]), .B(n164), .C(n161), .D(\mem[1][3] ), 
        .Z(n285) );
  HS65_LS_AO22X9 U135 ( .A(wr_data[4]), .B(n164), .C(n161), .D(\mem[1][4] ), 
        .Z(n284) );
  HS65_LS_AO22X9 U136 ( .A(wr_data[5]), .B(n164), .C(n161), .D(\mem[1][5] ), 
        .Z(n283) );
  HS65_LS_AO22X9 U137 ( .A(wr_data[6]), .B(n164), .C(n161), .D(\mem[1][6] ), 
        .Z(n282) );
  HS65_LS_AO22X9 U138 ( .A(wr_data[7]), .B(n164), .C(n161), .D(\mem[1][7] ), 
        .Z(n281) );
  HS65_LS_AO22X9 U139 ( .A(wr_data[8]), .B(n164), .C(n161), .D(\mem[1][8] ), 
        .Z(n280) );
  HS65_LS_AO22X9 U140 ( .A(wr_data[9]), .B(n164), .C(n161), .D(\mem[1][9] ), 
        .Z(n279) );
  HS65_LS_AO22X9 U141 ( .A(wr_data[10]), .B(n164), .C(n161), .D(\mem[1][10] ), 
        .Z(n278) );
  HS65_LS_AO22X9 U142 ( .A(wr_data[11]), .B(n163), .C(n161), .D(\mem[1][11] ), 
        .Z(n277) );
  HS65_LS_AO22X9 U143 ( .A(wr_data[12]), .B(n163), .C(n161), .D(\mem[1][12] ), 
        .Z(n276) );
  HS65_LS_AO22X9 U144 ( .A(wr_data[13]), .B(n163), .C(n161), .D(\mem[1][13] ), 
        .Z(n275) );
  HS65_LS_AO22X9 U145 ( .A(wr_data[14]), .B(n163), .C(n161), .D(\mem[1][14] ), 
        .Z(n274) );
  HS65_LS_AO22X9 U146 ( .A(wr_data[15]), .B(n163), .C(n161), .D(\mem[1][15] ), 
        .Z(n273) );
  HS65_LS_AO22X9 U147 ( .A(wr_data[16]), .B(n163), .C(n161), .D(\mem[1][16] ), 
        .Z(n272) );
  HS65_LS_AO22X9 U148 ( .A(wr_data[17]), .B(n163), .C(n161), .D(\mem[1][17] ), 
        .Z(n271) );
  HS65_LS_AO22X9 U149 ( .A(wr_data[18]), .B(n163), .C(n161), .D(\mem[1][18] ), 
        .Z(n270) );
  HS65_LS_AO22X9 U150 ( .A(wr_data[19]), .B(n163), .C(n161), .D(\mem[1][19] ), 
        .Z(n269) );
  HS65_LS_AO22X9 U151 ( .A(wr_data[20]), .B(n163), .C(n327), .D(\mem[1][20] ), 
        .Z(n268) );
  HS65_LS_AO22X9 U152 ( .A(wr_data[21]), .B(n163), .C(n327), .D(\mem[1][21] ), 
        .Z(n267) );
  HS65_LS_AO22X9 U153 ( .A(wr_data[22]), .B(n163), .C(n327), .D(\mem[1][22] ), 
        .Z(n266) );
  HS65_LS_AO22X9 U154 ( .A(wr_data[23]), .B(n163), .C(n327), .D(\mem[1][23] ), 
        .Z(n265) );
  HS65_LS_AO22X9 U155 ( .A(wr_data[24]), .B(n163), .C(n327), .D(\mem[1][24] ), 
        .Z(n264) );
  HS65_LS_AO22X9 U156 ( .A(wr_data[25]), .B(n163), .C(n327), .D(\mem[1][25] ), 
        .Z(n263) );
  HS65_LS_AO22X9 U157 ( .A(wr_data[26]), .B(n163), .C(n327), .D(\mem[1][26] ), 
        .Z(n262) );
  HS65_LS_AO22X9 U158 ( .A(wr_data[27]), .B(n163), .C(n327), .D(\mem[1][27] ), 
        .Z(n261) );
  HS65_LS_AO22X9 U159 ( .A(wr_data[28]), .B(n163), .C(n327), .D(\mem[1][28] ), 
        .Z(n260) );
  HS65_LS_AO22X9 U160 ( .A(wr_data[29]), .B(n163), .C(n327), .D(\mem[1][29] ), 
        .Z(n259) );
  HS65_LS_AO22X9 U161 ( .A(wr_data[30]), .B(n163), .C(n327), .D(\mem[1][30] ), 
        .Z(n258) );
  HS65_LS_AO22X9 U162 ( .A(wr_data[31]), .B(n162), .C(n327), .D(\mem[1][31] ), 
        .Z(n257) );
  HS65_LS_AO22X9 U163 ( .A(n170), .B(wr_data[0]), .C(n167), .D(\mem[0][0] ), 
        .Z(n320) );
  HS65_LS_AO22X9 U164 ( .A(n170), .B(wr_data[1]), .C(n166), .D(\mem[0][1] ), 
        .Z(n319) );
  HS65_LS_AO22X9 U165 ( .A(n170), .B(wr_data[2]), .C(n167), .D(\mem[0][2] ), 
        .Z(n318) );
  HS65_LS_AO22X9 U166 ( .A(n170), .B(wr_data[3]), .C(n166), .D(\mem[0][3] ), 
        .Z(n317) );
  HS65_LS_AO22X9 U167 ( .A(n170), .B(wr_data[4]), .C(n167), .D(\mem[0][4] ), 
        .Z(n316) );
  HS65_LS_AO22X9 U168 ( .A(n170), .B(wr_data[5]), .C(n166), .D(\mem[0][5] ), 
        .Z(n315) );
  HS65_LS_AO22X9 U169 ( .A(n170), .B(wr_data[6]), .C(n167), .D(\mem[0][6] ), 
        .Z(n314) );
  HS65_LS_AO22X9 U170 ( .A(n170), .B(wr_data[7]), .C(n167), .D(\mem[0][7] ), 
        .Z(n313) );
  HS65_LS_AO22X9 U171 ( .A(n170), .B(wr_data[8]), .C(n167), .D(\mem[0][8] ), 
        .Z(n312) );
  HS65_LS_AO22X9 U172 ( .A(n170), .B(wr_data[9]), .C(n167), .D(\mem[0][9] ), 
        .Z(n311) );
  HS65_LS_AO22X9 U173 ( .A(n170), .B(wr_data[10]), .C(n167), .D(\mem[0][10] ), 
        .Z(n310) );
  HS65_LS_AO22X9 U174 ( .A(n169), .B(wr_data[11]), .C(n167), .D(\mem[0][11] ), 
        .Z(n309) );
  HS65_LS_AO22X9 U175 ( .A(n169), .B(wr_data[12]), .C(n167), .D(\mem[0][12] ), 
        .Z(n308) );
  HS65_LS_AO22X9 U176 ( .A(n169), .B(wr_data[13]), .C(n167), .D(\mem[0][13] ), 
        .Z(n307) );
  HS65_LS_AO22X9 U177 ( .A(n169), .B(wr_data[14]), .C(n167), .D(\mem[0][14] ), 
        .Z(n306) );
  HS65_LS_AO22X9 U178 ( .A(n169), .B(wr_data[15]), .C(n167), .D(\mem[0][15] ), 
        .Z(n305) );
  HS65_LS_AO22X9 U179 ( .A(n169), .B(wr_data[16]), .C(n167), .D(\mem[0][16] ), 
        .Z(n304) );
  HS65_LS_AO22X9 U180 ( .A(n169), .B(wr_data[17]), .C(n167), .D(\mem[0][17] ), 
        .Z(n303) );
  HS65_LS_AO22X9 U181 ( .A(n169), .B(wr_data[18]), .C(n167), .D(\mem[0][18] ), 
        .Z(n302) );
  HS65_LS_AO22X9 U182 ( .A(n169), .B(wr_data[19]), .C(n166), .D(\mem[0][19] ), 
        .Z(n301) );
  HS65_LS_AO22X9 U183 ( .A(n169), .B(wr_data[20]), .C(n166), .D(\mem[0][20] ), 
        .Z(n300) );
  HS65_LS_AO22X9 U184 ( .A(n169), .B(wr_data[21]), .C(n166), .D(\mem[0][21] ), 
        .Z(n299) );
  HS65_LS_AO22X9 U185 ( .A(n169), .B(wr_data[22]), .C(n166), .D(\mem[0][22] ), 
        .Z(n298) );
  HS65_LS_AO22X9 U186 ( .A(n169), .B(wr_data[23]), .C(n166), .D(\mem[0][23] ), 
        .Z(n297) );
  HS65_LS_AO22X9 U187 ( .A(n169), .B(wr_data[24]), .C(n166), .D(\mem[0][24] ), 
        .Z(n296) );
  HS65_LS_AO22X9 U188 ( .A(n169), .B(wr_data[25]), .C(n166), .D(\mem[0][25] ), 
        .Z(n295) );
  HS65_LS_AO22X9 U189 ( .A(n169), .B(wr_data[26]), .C(n166), .D(\mem[0][26] ), 
        .Z(n294) );
  HS65_LS_AO22X9 U190 ( .A(n169), .B(wr_data[27]), .C(n166), .D(\mem[0][27] ), 
        .Z(n293) );
  HS65_LS_AO22X9 U191 ( .A(n169), .B(wr_data[28]), .C(n166), .D(\mem[0][28] ), 
        .Z(n292) );
  HS65_LS_AO22X9 U192 ( .A(n169), .B(wr_data[29]), .C(n166), .D(\mem[0][29] ), 
        .Z(n291) );
  HS65_LS_AO22X9 U193 ( .A(n169), .B(wr_data[30]), .C(n166), .D(\mem[0][30] ), 
        .Z(n290) );
  HS65_LS_AO22X9 U194 ( .A(n168), .B(wr_data[31]), .C(n166), .D(\mem[0][31] ), 
        .Z(n289) );
  HS65_LS_AO22X9 U195 ( .A(wr_data[0]), .B(n159), .C(n156), .D(\mem[2][0] ), 
        .Z(n256) );
  HS65_LS_AO22X9 U196 ( .A(wr_data[1]), .B(n159), .C(n156), .D(\mem[2][1] ), 
        .Z(n255) );
  HS65_LS_AO22X9 U197 ( .A(wr_data[2]), .B(n159), .C(n156), .D(\mem[2][2] ), 
        .Z(n254) );
  HS65_LS_AO22X9 U198 ( .A(wr_data[3]), .B(n159), .C(n156), .D(\mem[2][3] ), 
        .Z(n253) );
  HS65_LS_AO22X9 U199 ( .A(wr_data[4]), .B(n159), .C(n156), .D(\mem[2][4] ), 
        .Z(n252) );
  HS65_LS_AO22X9 U200 ( .A(wr_data[5]), .B(n159), .C(n156), .D(\mem[2][5] ), 
        .Z(n251) );
  HS65_LS_AO22X9 U201 ( .A(wr_data[6]), .B(n159), .C(n156), .D(\mem[2][6] ), 
        .Z(n250) );
  HS65_LS_AO22X9 U202 ( .A(wr_data[7]), .B(n159), .C(n156), .D(\mem[2][7] ), 
        .Z(n249) );
  HS65_LS_AO22X9 U203 ( .A(wr_data[8]), .B(n159), .C(n156), .D(\mem[2][8] ), 
        .Z(n248) );
  HS65_LS_AO22X9 U204 ( .A(wr_data[9]), .B(n159), .C(n156), .D(\mem[2][9] ), 
        .Z(n247) );
  HS65_LS_AO22X9 U205 ( .A(wr_data[10]), .B(n159), .C(n156), .D(\mem[2][10] ), 
        .Z(n246) );
  HS65_LS_AO22X9 U206 ( .A(wr_data[11]), .B(n158), .C(n156), .D(\mem[2][11] ), 
        .Z(n245) );
  HS65_LS_AO22X9 U207 ( .A(wr_data[12]), .B(n158), .C(n156), .D(\mem[2][12] ), 
        .Z(n244) );
  HS65_LS_AO22X9 U208 ( .A(wr_data[13]), .B(n158), .C(n156), .D(\mem[2][13] ), 
        .Z(n243) );
  HS65_LS_AO22X9 U209 ( .A(wr_data[14]), .B(n158), .C(n156), .D(\mem[2][14] ), 
        .Z(n242) );
  HS65_LS_AO22X9 U210 ( .A(wr_data[15]), .B(n158), .C(n156), .D(\mem[2][15] ), 
        .Z(n241) );
  HS65_LS_AO22X9 U211 ( .A(wr_data[16]), .B(n158), .C(n156), .D(\mem[2][16] ), 
        .Z(n240) );
  HS65_LS_AO22X9 U212 ( .A(wr_data[17]), .B(n158), .C(n156), .D(\mem[2][17] ), 
        .Z(n239) );
  HS65_LS_AO22X9 U213 ( .A(wr_data[18]), .B(n158), .C(n156), .D(\mem[2][18] ), 
        .Z(n238) );
  HS65_LS_AO22X9 U214 ( .A(wr_data[19]), .B(n158), .C(n156), .D(\mem[2][19] ), 
        .Z(n237) );
  HS65_LS_AO22X9 U215 ( .A(wr_data[20]), .B(n158), .C(n326), .D(\mem[2][20] ), 
        .Z(n236) );
  HS65_LS_AO22X9 U216 ( .A(wr_data[21]), .B(n158), .C(n326), .D(\mem[2][21] ), 
        .Z(n235) );
  HS65_LS_AO22X9 U217 ( .A(wr_data[22]), .B(n158), .C(n326), .D(\mem[2][22] ), 
        .Z(n234) );
  HS65_LS_AO22X9 U218 ( .A(wr_data[23]), .B(n158), .C(n326), .D(\mem[2][23] ), 
        .Z(n233) );
  HS65_LS_AO22X9 U219 ( .A(wr_data[24]), .B(n158), .C(n326), .D(\mem[2][24] ), 
        .Z(n232) );
  HS65_LS_AO22X9 U220 ( .A(wr_data[25]), .B(n158), .C(n326), .D(\mem[2][25] ), 
        .Z(n231) );
  HS65_LS_AO22X9 U221 ( .A(wr_data[26]), .B(n158), .C(n326), .D(\mem[2][26] ), 
        .Z(n230) );
  HS65_LS_AO22X9 U222 ( .A(wr_data[27]), .B(n158), .C(n326), .D(\mem[2][27] ), 
        .Z(n229) );
  HS65_LS_AO22X9 U223 ( .A(wr_data[28]), .B(n158), .C(n326), .D(\mem[2][28] ), 
        .Z(n228) );
  HS65_LS_AO22X9 U224 ( .A(wr_data[29]), .B(n158), .C(n326), .D(\mem[2][29] ), 
        .Z(n227) );
  HS65_LS_AO22X9 U225 ( .A(wr_data[30]), .B(n158), .C(n326), .D(\mem[2][30] ), 
        .Z(n226) );
  HS65_LS_AO22X9 U226 ( .A(wr_data[31]), .B(n157), .C(n326), .D(\mem[2][31] ), 
        .Z(n225) );
endmodule


module bram_DATA16_ADDR2_5 ( clk, reset, rd_addr, wr_addr, wr_data, wr_ena, 
        rd_data );
  input [1:0] rd_addr;
  input [1:0] wr_addr;
  input [15:0] wr_data;
  output [15:0] rd_data;
  input clk, reset, wr_ena;
  wire   \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] ,
         \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][15] , \mem[1][14] , \mem[1][13] ,
         \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] , \mem[1][8] ,
         \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] ,
         \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][15] , \mem[0][14] ,
         \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] ,
         \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] ,
         \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, n1,
         n2, n3, n4, n5, n6, n7, n8, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162;

  HS65_LS_DFPRQX9 \mem_reg[3][15]  ( .D(n91), .CP(clk), .RN(n1), .Q(
        \mem[3][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][14]  ( .D(n92), .CP(clk), .RN(n1), .Q(
        \mem[3][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][13]  ( .D(n93), .CP(clk), .RN(n1), .Q(
        \mem[3][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][12]  ( .D(n94), .CP(clk), .RN(n1), .Q(
        \mem[3][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][11]  ( .D(n95), .CP(clk), .RN(n1), .Q(
        \mem[3][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][10]  ( .D(n96), .CP(clk), .RN(n1), .Q(
        \mem[3][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][9]  ( .D(n97), .CP(clk), .RN(n1), .Q(\mem[3][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][8]  ( .D(n98), .CP(clk), .RN(n1), .Q(\mem[3][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][7]  ( .D(n99), .CP(clk), .RN(n1), .Q(\mem[3][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][6]  ( .D(n100), .CP(clk), .RN(n1), .Q(
        \mem[3][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][5]  ( .D(n101), .CP(clk), .RN(n1), .Q(
        \mem[3][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][4]  ( .D(n102), .CP(clk), .RN(n1), .Q(
        \mem[3][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][3]  ( .D(n103), .CP(clk), .RN(n1), .Q(
        \mem[3][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][2]  ( .D(n104), .CP(clk), .RN(n2), .Q(
        \mem[3][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][1]  ( .D(n105), .CP(clk), .RN(n2), .Q(
        \mem[3][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][0]  ( .D(n106), .CP(clk), .RN(n2), .Q(
        \mem[3][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][15]  ( .D(n107), .CP(clk), .RN(n2), .Q(
        \mem[2][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][14]  ( .D(n108), .CP(clk), .RN(n2), .Q(
        \mem[2][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][13]  ( .D(n109), .CP(clk), .RN(n2), .Q(
        \mem[2][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][12]  ( .D(n110), .CP(clk), .RN(n2), .Q(
        \mem[2][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][11]  ( .D(n111), .CP(clk), .RN(n2), .Q(
        \mem[2][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][10]  ( .D(n112), .CP(clk), .RN(n2), .Q(
        \mem[2][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][9]  ( .D(n113), .CP(clk), .RN(n2), .Q(
        \mem[2][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][8]  ( .D(n114), .CP(clk), .RN(n2), .Q(
        \mem[2][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][7]  ( .D(n115), .CP(clk), .RN(n2), .Q(
        \mem[2][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][6]  ( .D(n116), .CP(clk), .RN(n2), .Q(
        \mem[2][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][5]  ( .D(n117), .CP(clk), .RN(n3), .Q(
        \mem[2][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][4]  ( .D(n118), .CP(clk), .RN(n3), .Q(
        \mem[2][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][3]  ( .D(n119), .CP(clk), .RN(n3), .Q(
        \mem[2][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][2]  ( .D(n120), .CP(clk), .RN(n3), .Q(
        \mem[2][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][1]  ( .D(n121), .CP(clk), .RN(n3), .Q(
        \mem[2][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][0]  ( .D(n122), .CP(clk), .RN(n3), .Q(
        \mem[2][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][15]  ( .D(n123), .CP(clk), .RN(n3), .Q(
        \mem[1][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][14]  ( .D(n124), .CP(clk), .RN(n3), .Q(
        \mem[1][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][13]  ( .D(n125), .CP(clk), .RN(n3), .Q(
        \mem[1][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][12]  ( .D(n126), .CP(clk), .RN(n3), .Q(
        \mem[1][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][11]  ( .D(n127), .CP(clk), .RN(n3), .Q(
        \mem[1][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][10]  ( .D(n128), .CP(clk), .RN(n3), .Q(
        \mem[1][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][9]  ( .D(n129), .CP(clk), .RN(n3), .Q(
        \mem[1][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][8]  ( .D(n130), .CP(clk), .RN(n4), .Q(
        \mem[1][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][7]  ( .D(n131), .CP(clk), .RN(n4), .Q(
        \mem[1][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][6]  ( .D(n132), .CP(clk), .RN(n4), .Q(
        \mem[1][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][5]  ( .D(n133), .CP(clk), .RN(n4), .Q(
        \mem[1][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][4]  ( .D(n134), .CP(clk), .RN(n4), .Q(
        \mem[1][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][3]  ( .D(n135), .CP(clk), .RN(n4), .Q(
        \mem[1][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][2]  ( .D(n136), .CP(clk), .RN(n4), .Q(
        \mem[1][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][1]  ( .D(n137), .CP(clk), .RN(n4), .Q(
        \mem[1][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][0]  ( .D(n138), .CP(clk), .RN(n4), .Q(
        \mem[1][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][15]  ( .D(n139), .CP(clk), .RN(n4), .Q(
        \mem[0][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][14]  ( .D(n140), .CP(clk), .RN(n4), .Q(
        \mem[0][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][13]  ( .D(n141), .CP(clk), .RN(n4), .Q(
        \mem[0][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][12]  ( .D(n142), .CP(clk), .RN(n4), .Q(
        \mem[0][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][11]  ( .D(n143), .CP(clk), .RN(n5), .Q(
        \mem[0][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][10]  ( .D(n144), .CP(clk), .RN(n5), .Q(
        \mem[0][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][9]  ( .D(n145), .CP(clk), .RN(n5), .Q(
        \mem[0][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][8]  ( .D(n146), .CP(clk), .RN(n5), .Q(
        \mem[0][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][7]  ( .D(n147), .CP(clk), .RN(n5), .Q(
        \mem[0][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][6]  ( .D(n148), .CP(clk), .RN(n5), .Q(
        \mem[0][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][5]  ( .D(n149), .CP(clk), .RN(n5), .Q(
        \mem[0][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][4]  ( .D(n150), .CP(clk), .RN(n5), .Q(
        \mem[0][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][3]  ( .D(n151), .CP(clk), .RN(n5), .Q(
        \mem[0][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][2]  ( .D(n152), .CP(clk), .RN(n5), .Q(
        \mem[0][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][1]  ( .D(n153), .CP(clk), .RN(n5), .Q(
        \mem[0][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][0]  ( .D(n154), .CP(clk), .RN(n5), .Q(
        \mem[0][0] ) );
  HS65_LS_DFPRQX9 \rd_data_reg[15]  ( .D(N17), .CP(clk), .RN(n5), .Q(
        rd_data[15]) );
  HS65_LS_DFPRQX9 \rd_data_reg[14]  ( .D(N18), .CP(clk), .RN(n6), .Q(
        rd_data[14]) );
  HS65_LS_DFPRQX9 \rd_data_reg[13]  ( .D(N19), .CP(clk), .RN(n6), .Q(
        rd_data[13]) );
  HS65_LS_DFPRQX9 \rd_data_reg[12]  ( .D(N20), .CP(clk), .RN(n6), .Q(
        rd_data[12]) );
  HS65_LS_DFPRQX9 \rd_data_reg[11]  ( .D(N21), .CP(clk), .RN(n6), .Q(
        rd_data[11]) );
  HS65_LS_DFPRQX9 \rd_data_reg[10]  ( .D(N22), .CP(clk), .RN(n6), .Q(
        rd_data[10]) );
  HS65_LS_DFPRQX9 \rd_data_reg[9]  ( .D(N23), .CP(clk), .RN(n6), .Q(rd_data[9]) );
  HS65_LS_DFPRQX9 \rd_data_reg[8]  ( .D(N24), .CP(clk), .RN(n6), .Q(rd_data[8]) );
  HS65_LS_DFPRQX9 \rd_data_reg[7]  ( .D(N25), .CP(clk), .RN(n6), .Q(rd_data[7]) );
  HS65_LS_DFPRQX9 \rd_data_reg[6]  ( .D(N26), .CP(clk), .RN(n6), .Q(rd_data[6]) );
  HS65_LS_DFPRQX9 \rd_data_reg[5]  ( .D(N27), .CP(clk), .RN(n6), .Q(rd_data[5]) );
  HS65_LS_DFPRQX9 \rd_data_reg[4]  ( .D(N28), .CP(clk), .RN(n6), .Q(rd_data[4]) );
  HS65_LS_DFPRQX9 \rd_data_reg[3]  ( .D(N29), .CP(clk), .RN(n6), .Q(rd_data[3]) );
  HS65_LS_DFPRQX9 \rd_data_reg[2]  ( .D(N30), .CP(clk), .RN(n6), .Q(rd_data[2]) );
  HS65_LS_DFPRQX9 \rd_data_reg[1]  ( .D(N31), .CP(clk), .RN(n7), .Q(rd_data[1]) );
  HS65_LS_DFPRQX9 \rd_data_reg[0]  ( .D(N32), .CP(clk), .RN(n7), .Q(rd_data[0]) );
  HS65_LS_BFX9 U3 ( .A(n81), .Z(n4) );
  HS65_LS_BFX9 U4 ( .A(n81), .Z(n3) );
  HS65_LS_BFX9 U5 ( .A(n81), .Z(n2) );
  HS65_LS_BFX9 U6 ( .A(n83), .Z(n81) );
  HS65_LS_BFX9 U7 ( .A(n8), .Z(n6) );
  HS65_LS_BFX9 U8 ( .A(n8), .Z(n5) );
  HS65_LS_BFX9 U9 ( .A(n82), .Z(n1) );
  HS65_LS_BFX9 U10 ( .A(n83), .Z(n82) );
  HS65_LS_BFX9 U11 ( .A(n8), .Z(n7) );
  HS65_LS_BFX9 U12 ( .A(n83), .Z(n8) );
  HS65_LS_IVX9 U13 ( .A(reset), .Z(n83) );
  HS65_LS_IVX9 U14 ( .A(n161), .Z(n85) );
  HS65_LS_IVX9 U15 ( .A(n162), .Z(n84) );
  HS65_LS_NAND3X5 U16 ( .A(wr_ena), .B(n86), .C(wr_addr[0]), .Z(n161) );
  HS65_LS_IVX9 U17 ( .A(wr_addr[0]), .Z(n89) );
  HS65_LS_NAND3X5 U18 ( .A(n89), .B(n86), .C(wr_ena), .Z(n162) );
  HS65_LS_IVX9 U19 ( .A(n160), .Z(n88) );
  HS65_LS_IVX9 U20 ( .A(n159), .Z(n87) );
  HS65_LS_NAND3X5 U21 ( .A(wr_ena), .B(n89), .C(wr_addr[1]), .Z(n160) );
  HS65_LS_NOR2X6 U22 ( .A(n90), .B(rd_addr[1]), .Z(n157) );
  HS65_LS_NOR2X6 U23 ( .A(rd_addr[0]), .B(rd_addr[1]), .Z(n158) );
  HS65_LS_IVX9 U24 ( .A(wr_addr[1]), .Z(n86) );
  HS65_LS_NAND3X5 U25 ( .A(wr_addr[0]), .B(wr_ena), .C(wr_addr[1]), .Z(n159)
         );
  HS65_LS_AND2X4 U26 ( .A(rd_addr[1]), .B(n90), .Z(n156) );
  HS65_LS_AND2X4 U27 ( .A(rd_addr[1]), .B(rd_addr[0]), .Z(n155) );
  HS65_LS_IVX9 U28 ( .A(rd_addr[0]), .Z(n90) );
  HS65_LS_MX41X7 U29 ( .D0(n158), .S0(\mem[0][0] ), .D1(n157), .S1(\mem[1][0] ), .D2(n156), .S2(\mem[2][0] ), .D3(n155), .S3(\mem[3][0] ), .Z(N32) );
  HS65_LS_MX41X7 U30 ( .D0(n158), .S0(\mem[0][1] ), .D1(n157), .S1(\mem[1][1] ), .D2(n156), .S2(\mem[2][1] ), .D3(n155), .S3(\mem[3][1] ), .Z(N31) );
  HS65_LS_MX41X7 U31 ( .D0(n158), .S0(\mem[0][2] ), .D1(n157), .S1(\mem[1][2] ), .D2(n156), .S2(\mem[2][2] ), .D3(n155), .S3(\mem[3][2] ), .Z(N30) );
  HS65_LS_MX41X7 U32 ( .D0(n158), .S0(\mem[0][3] ), .D1(n157), .S1(\mem[1][3] ), .D2(n156), .S2(\mem[2][3] ), .D3(n155), .S3(\mem[3][3] ), .Z(N29) );
  HS65_LS_MX41X7 U33 ( .D0(n158), .S0(\mem[0][4] ), .D1(n157), .S1(\mem[1][4] ), .D2(n156), .S2(\mem[2][4] ), .D3(n155), .S3(\mem[3][4] ), .Z(N28) );
  HS65_LS_MX41X7 U34 ( .D0(n158), .S0(\mem[0][5] ), .D1(n157), .S1(\mem[1][5] ), .D2(n156), .S2(\mem[2][5] ), .D3(n155), .S3(\mem[3][5] ), .Z(N27) );
  HS65_LS_MX41X7 U35 ( .D0(n158), .S0(\mem[0][6] ), .D1(n157), .S1(\mem[1][6] ), .D2(n156), .S2(\mem[2][6] ), .D3(n155), .S3(\mem[3][6] ), .Z(N26) );
  HS65_LS_MX41X7 U36 ( .D0(n158), .S0(\mem[0][7] ), .D1(n157), .S1(\mem[1][7] ), .D2(n156), .S2(\mem[2][7] ), .D3(n155), .S3(\mem[3][7] ), .Z(N25) );
  HS65_LS_MX41X7 U37 ( .D0(n158), .S0(\mem[0][8] ), .D1(n157), .S1(\mem[1][8] ), .D2(n156), .S2(\mem[2][8] ), .D3(n155), .S3(\mem[3][8] ), .Z(N24) );
  HS65_LS_MX41X7 U38 ( .D0(n158), .S0(\mem[0][9] ), .D1(n157), .S1(\mem[1][9] ), .D2(n156), .S2(\mem[2][9] ), .D3(n155), .S3(\mem[3][9] ), .Z(N23) );
  HS65_LS_MX41X7 U39 ( .D0(n158), .S0(\mem[0][10] ), .D1(n157), .S1(
        \mem[1][10] ), .D2(n156), .S2(\mem[2][10] ), .D3(n155), .S3(
        \mem[3][10] ), .Z(N22) );
  HS65_LS_MX41X7 U40 ( .D0(n158), .S0(\mem[0][11] ), .D1(n157), .S1(
        \mem[1][11] ), .D2(n156), .S2(\mem[2][11] ), .D3(n155), .S3(
        \mem[3][11] ), .Z(N21) );
  HS65_LS_MX41X7 U41 ( .D0(n158), .S0(\mem[0][12] ), .D1(n157), .S1(
        \mem[1][12] ), .D2(n156), .S2(\mem[2][12] ), .D3(n155), .S3(
        \mem[3][12] ), .Z(N20) );
  HS65_LS_MX41X7 U42 ( .D0(n158), .S0(\mem[0][13] ), .D1(n157), .S1(
        \mem[1][13] ), .D2(n156), .S2(\mem[2][13] ), .D3(n155), .S3(
        \mem[3][13] ), .Z(N19) );
  HS65_LS_MX41X7 U43 ( .D0(n158), .S0(\mem[0][14] ), .D1(n157), .S1(
        \mem[1][14] ), .D2(n156), .S2(\mem[2][14] ), .D3(n155), .S3(
        \mem[3][14] ), .Z(N18) );
  HS65_LS_MX41X7 U44 ( .D0(n158), .S0(\mem[0][15] ), .D1(n157), .S1(
        \mem[1][15] ), .D2(n156), .S2(\mem[2][15] ), .D3(n155), .S3(
        \mem[3][15] ), .Z(N17) );
  HS65_LS_AO22X9 U45 ( .A(wr_data[0]), .B(n85), .C(n161), .D(\mem[1][0] ), .Z(
        n138) );
  HS65_LS_AO22X9 U46 ( .A(wr_data[1]), .B(n85), .C(n161), .D(\mem[1][1] ), .Z(
        n137) );
  HS65_LS_AO22X9 U47 ( .A(wr_data[2]), .B(n85), .C(n161), .D(\mem[1][2] ), .Z(
        n136) );
  HS65_LS_AO22X9 U48 ( .A(wr_data[3]), .B(n85), .C(n161), .D(\mem[1][3] ), .Z(
        n135) );
  HS65_LS_AO22X9 U49 ( .A(wr_data[4]), .B(n85), .C(n161), .D(\mem[1][4] ), .Z(
        n134) );
  HS65_LS_AO22X9 U50 ( .A(wr_data[5]), .B(n85), .C(n161), .D(\mem[1][5] ), .Z(
        n133) );
  HS65_LS_AO22X9 U51 ( .A(wr_data[6]), .B(n85), .C(n161), .D(\mem[1][6] ), .Z(
        n132) );
  HS65_LS_AO22X9 U52 ( .A(wr_data[7]), .B(n85), .C(n161), .D(\mem[1][7] ), .Z(
        n131) );
  HS65_LS_AO22X9 U53 ( .A(wr_data[8]), .B(n85), .C(n161), .D(\mem[1][8] ), .Z(
        n130) );
  HS65_LS_AO22X9 U54 ( .A(wr_data[9]), .B(n85), .C(n161), .D(\mem[1][9] ), .Z(
        n129) );
  HS65_LS_AO22X9 U55 ( .A(wr_data[10]), .B(n85), .C(n161), .D(\mem[1][10] ), 
        .Z(n128) );
  HS65_LS_AO22X9 U56 ( .A(wr_data[11]), .B(n85), .C(n161), .D(\mem[1][11] ), 
        .Z(n127) );
  HS65_LS_AO22X9 U57 ( .A(wr_data[12]), .B(n85), .C(n161), .D(\mem[1][12] ), 
        .Z(n126) );
  HS65_LS_AO22X9 U58 ( .A(wr_data[13]), .B(n85), .C(n161), .D(\mem[1][13] ), 
        .Z(n125) );
  HS65_LS_AO22X9 U59 ( .A(wr_data[14]), .B(n85), .C(n161), .D(\mem[1][14] ), 
        .Z(n124) );
  HS65_LS_AO22X9 U60 ( .A(wr_data[15]), .B(n85), .C(n161), .D(\mem[1][15] ), 
        .Z(n123) );
  HS65_LS_AO22X9 U61 ( .A(wr_data[0]), .B(n88), .C(n160), .D(\mem[2][0] ), .Z(
        n122) );
  HS65_LS_AO22X9 U62 ( .A(wr_data[1]), .B(n88), .C(n160), .D(\mem[2][1] ), .Z(
        n121) );
  HS65_LS_AO22X9 U63 ( .A(wr_data[2]), .B(n88), .C(n160), .D(\mem[2][2] ), .Z(
        n120) );
  HS65_LS_AO22X9 U64 ( .A(wr_data[3]), .B(n88), .C(n160), .D(\mem[2][3] ), .Z(
        n119) );
  HS65_LS_AO22X9 U65 ( .A(wr_data[4]), .B(n88), .C(n160), .D(\mem[2][4] ), .Z(
        n118) );
  HS65_LS_AO22X9 U66 ( .A(wr_data[5]), .B(n88), .C(n160), .D(\mem[2][5] ), .Z(
        n117) );
  HS65_LS_AO22X9 U67 ( .A(wr_data[6]), .B(n88), .C(n160), .D(\mem[2][6] ), .Z(
        n116) );
  HS65_LS_AO22X9 U68 ( .A(wr_data[7]), .B(n88), .C(n160), .D(\mem[2][7] ), .Z(
        n115) );
  HS65_LS_AO22X9 U69 ( .A(wr_data[8]), .B(n88), .C(n160), .D(\mem[2][8] ), .Z(
        n114) );
  HS65_LS_AO22X9 U70 ( .A(wr_data[9]), .B(n88), .C(n160), .D(\mem[2][9] ), .Z(
        n113) );
  HS65_LS_AO22X9 U71 ( .A(wr_data[10]), .B(n88), .C(n160), .D(\mem[2][10] ), 
        .Z(n112) );
  HS65_LS_AO22X9 U72 ( .A(wr_data[11]), .B(n88), .C(n160), .D(\mem[2][11] ), 
        .Z(n111) );
  HS65_LS_AO22X9 U73 ( .A(wr_data[12]), .B(n88), .C(n160), .D(\mem[2][12] ), 
        .Z(n110) );
  HS65_LS_AO22X9 U74 ( .A(wr_data[13]), .B(n88), .C(n160), .D(\mem[2][13] ), 
        .Z(n109) );
  HS65_LS_AO22X9 U75 ( .A(wr_data[14]), .B(n88), .C(n160), .D(\mem[2][14] ), 
        .Z(n108) );
  HS65_LS_AO22X9 U76 ( .A(wr_data[15]), .B(n88), .C(n160), .D(\mem[2][15] ), 
        .Z(n107) );
  HS65_LS_AO22X9 U77 ( .A(n84), .B(wr_data[0]), .C(n162), .D(\mem[0][0] ), .Z(
        n154) );
  HS65_LS_AO22X9 U78 ( .A(n84), .B(wr_data[1]), .C(n162), .D(\mem[0][1] ), .Z(
        n153) );
  HS65_LS_AO22X9 U79 ( .A(n84), .B(wr_data[2]), .C(n162), .D(\mem[0][2] ), .Z(
        n152) );
  HS65_LS_AO22X9 U80 ( .A(n84), .B(wr_data[3]), .C(n162), .D(\mem[0][3] ), .Z(
        n151) );
  HS65_LS_AO22X9 U81 ( .A(n84), .B(wr_data[4]), .C(n162), .D(\mem[0][4] ), .Z(
        n150) );
  HS65_LS_AO22X9 U82 ( .A(n84), .B(wr_data[5]), .C(n162), .D(\mem[0][5] ), .Z(
        n149) );
  HS65_LS_AO22X9 U83 ( .A(n84), .B(wr_data[6]), .C(n162), .D(\mem[0][6] ), .Z(
        n148) );
  HS65_LS_AO22X9 U84 ( .A(n84), .B(wr_data[7]), .C(n162), .D(\mem[0][7] ), .Z(
        n147) );
  HS65_LS_AO22X9 U85 ( .A(n84), .B(wr_data[8]), .C(n162), .D(\mem[0][8] ), .Z(
        n146) );
  HS65_LS_AO22X9 U86 ( .A(n84), .B(wr_data[9]), .C(n162), .D(\mem[0][9] ), .Z(
        n145) );
  HS65_LS_AO22X9 U87 ( .A(n84), .B(wr_data[10]), .C(n162), .D(\mem[0][10] ), 
        .Z(n144) );
  HS65_LS_AO22X9 U88 ( .A(n84), .B(wr_data[11]), .C(n162), .D(\mem[0][11] ), 
        .Z(n143) );
  HS65_LS_AO22X9 U89 ( .A(n84), .B(wr_data[12]), .C(n162), .D(\mem[0][12] ), 
        .Z(n142) );
  HS65_LS_AO22X9 U90 ( .A(n84), .B(wr_data[13]), .C(n162), .D(\mem[0][13] ), 
        .Z(n141) );
  HS65_LS_AO22X9 U91 ( .A(n84), .B(wr_data[14]), .C(n162), .D(\mem[0][14] ), 
        .Z(n140) );
  HS65_LS_AO22X9 U92 ( .A(n84), .B(wr_data[15]), .C(n162), .D(\mem[0][15] ), 
        .Z(n139) );
  HS65_LS_AO22X9 U93 ( .A(wr_data[0]), .B(n87), .C(n159), .D(\mem[3][0] ), .Z(
        n106) );
  HS65_LS_AO22X9 U94 ( .A(wr_data[1]), .B(n87), .C(n159), .D(\mem[3][1] ), .Z(
        n105) );
  HS65_LS_AO22X9 U95 ( .A(wr_data[2]), .B(n87), .C(n159), .D(\mem[3][2] ), .Z(
        n104) );
  HS65_LS_AO22X9 U96 ( .A(wr_data[3]), .B(n87), .C(n159), .D(\mem[3][3] ), .Z(
        n103) );
  HS65_LS_AO22X9 U97 ( .A(wr_data[4]), .B(n87), .C(n159), .D(\mem[3][4] ), .Z(
        n102) );
  HS65_LS_AO22X9 U98 ( .A(wr_data[5]), .B(n87), .C(n159), .D(\mem[3][5] ), .Z(
        n101) );
  HS65_LS_AO22X9 U99 ( .A(wr_data[6]), .B(n87), .C(n159), .D(\mem[3][6] ), .Z(
        n100) );
  HS65_LS_AO22X9 U100 ( .A(wr_data[7]), .B(n87), .C(n159), .D(\mem[3][7] ), 
        .Z(n99) );
  HS65_LS_AO22X9 U101 ( .A(wr_data[8]), .B(n87), .C(n159), .D(\mem[3][8] ), 
        .Z(n98) );
  HS65_LS_AO22X9 U102 ( .A(wr_data[9]), .B(n87), .C(n159), .D(\mem[3][9] ), 
        .Z(n97) );
  HS65_LS_AO22X9 U103 ( .A(wr_data[10]), .B(n87), .C(n159), .D(\mem[3][10] ), 
        .Z(n96) );
  HS65_LS_AO22X9 U104 ( .A(wr_data[11]), .B(n87), .C(n159), .D(\mem[3][11] ), 
        .Z(n95) );
  HS65_LS_AO22X9 U105 ( .A(wr_data[12]), .B(n87), .C(n159), .D(\mem[3][12] ), 
        .Z(n94) );
  HS65_LS_AO22X9 U106 ( .A(wr_data[13]), .B(n87), .C(n159), .D(\mem[3][13] ), 
        .Z(n93) );
  HS65_LS_AO22X9 U107 ( .A(wr_data[14]), .B(n87), .C(n159), .D(\mem[3][14] ), 
        .Z(n92) );
  HS65_LS_AO22X9 U108 ( .A(wr_data[15]), .B(n87), .C(n159), .D(\mem[3][15] ), 
        .Z(n91) );
endmodule


module dma_sdp_DATA64_ADDR2_3 ( clk, reset, ren, wen, waddr, wdata, raddr, 
        rdata );
  input [2:0] ren;
  input [2:0] wen;
  input [1:0] waddr;
  input [63:0] wdata;
  input [1:0] raddr;
  output [63:0] rdata;
  input clk, reset;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n41, n42, n43, n44, n45, n46, n47, n48;
  wire   [2:0] sel_out;
  wire   [15:0] rdata0;
  wire   [31:0] rdata1;
  wire   [15:0] rdata2;

  HS65_LS_DFPRQX9 \sel_out_reg[2]  ( .D(ren[2]), .CP(clk), .RN(n5), .Q(
        sel_out[2]) );
  HS65_LS_DFPRQX9 \sel_out_reg[1]  ( .D(ren[1]), .CP(clk), .RN(n5), .Q(
        sel_out[1]) );
  HS65_LS_DFPRQX9 \sel_out_reg[0]  ( .D(ren[0]), .CP(clk), .RN(n5), .Q(
        sel_out[0]) );
  bram_DATA16_ADDR2_6 dma0 ( .clk(clk), .reset(reset), .rd_addr(raddr), 
        .wr_addr(waddr), .wr_data(wdata[63:48]), .wr_ena(wen[2]), .rd_data(
        rdata0) );
  bram_DATA32_ADDR2_3 dma1 ( .clk(clk), .reset(reset), .rd_addr(raddr), 
        .wr_addr(waddr), .wr_data(wdata[47:16]), .wr_ena(wen[1]), .rd_data(
        rdata1) );
  bram_DATA16_ADDR2_5 dma2 ( .clk(clk), .reset(reset), .rd_addr(raddr), 
        .wr_addr(waddr), .wr_data(wdata[15:0]), .wr_ena(wen[0]), .rd_data(
        rdata2) );
  HS65_LS_NAND3X5 U3 ( .A(sel_out[2]), .B(sel_out[1]), .C(sel_out[0]), .Z(n46)
         );
  HS65_LS_IVX9 U4 ( .A(reset), .Z(n5) );
  HS65_LS_NOR2X6 U5 ( .A(n2), .B(n13), .Z(rdata[40]) );
  HS65_LS_NOR2X6 U6 ( .A(n2), .B(n12), .Z(rdata[41]) );
  HS65_LS_NOR2X6 U7 ( .A(n2), .B(n11), .Z(rdata[42]) );
  HS65_LS_NOR2X6 U8 ( .A(n2), .B(n10), .Z(rdata[43]) );
  HS65_LS_NOR2X6 U9 ( .A(n2), .B(n9), .Z(rdata[44]) );
  HS65_LS_NOR2X6 U10 ( .A(n2), .B(n8), .Z(rdata[45]) );
  HS65_LS_NOR2X6 U11 ( .A(n2), .B(n7), .Z(rdata[46]) );
  HS65_LS_NOR2X6 U12 ( .A(n2), .B(n14), .Z(rdata[39]) );
  HS65_LS_BFX9 U13 ( .A(n46), .Z(n2) );
  HS65_LS_NOR2X6 U14 ( .A(n2), .B(n15), .Z(rdata[38]) );
  HS65_LS_NOR2X6 U15 ( .A(n3), .B(n19), .Z(rdata[34]) );
  HS65_LS_NOR2X6 U16 ( .A(n2), .B(n18), .Z(rdata[35]) );
  HS65_LS_NOR2X6 U17 ( .A(n3), .B(n17), .Z(rdata[36]) );
  HS65_LS_NOR2X6 U18 ( .A(n2), .B(n16), .Z(rdata[37]) );
  HS65_LS_NOR2X6 U19 ( .A(n3), .B(n20), .Z(rdata[33]) );
  HS65_LS_BFX9 U20 ( .A(n46), .Z(n3) );
  HS65_LS_BFX9 U21 ( .A(n46), .Z(n1) );
  HS65_LS_BFX9 U22 ( .A(n46), .Z(n4) );
  HS65_LS_IVX9 U23 ( .A(n45), .Z(n42) );
  HS65_LS_NOR2X6 U24 ( .A(n2), .B(n6), .Z(rdata[47]) );
  HS65_LS_NAND3X5 U25 ( .A(n44), .B(n43), .C(sel_out[1]), .Z(n45) );
  HS65_LS_IVX9 U26 ( .A(sel_out[0]), .Z(n44) );
  HS65_LS_IVX9 U27 ( .A(sel_out[2]), .Z(n43) );
  HS65_LS_OAI22X6 U28 ( .A(n45), .B(n19), .C(n1), .D(n35), .Z(rdata[18]) );
  HS65_LS_IVX9 U29 ( .A(rdata1[2]), .Z(n35) );
  HS65_LS_OAI22X6 U30 ( .A(n45), .B(n18), .C(n1), .D(n34), .Z(rdata[19]) );
  HS65_LS_IVX9 U31 ( .A(rdata1[3]), .Z(n34) );
  HS65_LS_OAI22X6 U32 ( .A(n45), .B(n17), .C(n1), .D(n33), .Z(rdata[20]) );
  HS65_LS_IVX9 U33 ( .A(rdata1[4]), .Z(n33) );
  HS65_LS_OAI22X6 U34 ( .A(n45), .B(n16), .C(n1), .D(n32), .Z(rdata[21]) );
  HS65_LS_IVX9 U35 ( .A(rdata1[5]), .Z(n32) );
  HS65_LS_OAI22X6 U36 ( .A(n45), .B(n15), .C(n31), .D(n3), .Z(rdata[22]) );
  HS65_LS_IVX9 U37 ( .A(rdata1[6]), .Z(n31) );
  HS65_LS_OAI22X6 U38 ( .A(n45), .B(n14), .C(n30), .D(n3), .Z(rdata[23]) );
  HS65_LS_IVX9 U39 ( .A(rdata1[7]), .Z(n30) );
  HS65_LS_OAI22X6 U40 ( .A(n45), .B(n13), .C(n29), .D(n3), .Z(rdata[24]) );
  HS65_LS_IVX9 U41 ( .A(rdata1[8]), .Z(n29) );
  HS65_LS_OAI22X6 U42 ( .A(n45), .B(n12), .C(n28), .D(n3), .Z(rdata[25]) );
  HS65_LS_IVX9 U43 ( .A(rdata1[9]), .Z(n28) );
  HS65_LS_OAI22X6 U44 ( .A(n45), .B(n11), .C(n1), .D(n27), .Z(rdata[26]) );
  HS65_LS_IVX9 U45 ( .A(rdata1[10]), .Z(n27) );
  HS65_LS_OAI22X6 U46 ( .A(n45), .B(n10), .C(n1), .D(n26), .Z(rdata[27]) );
  HS65_LS_IVX9 U47 ( .A(rdata1[11]), .Z(n26) );
  HS65_LS_OAI22X6 U48 ( .A(n45), .B(n20), .C(n1), .D(n36), .Z(rdata[17]) );
  HS65_LS_IVX9 U49 ( .A(rdata1[1]), .Z(n36) );
  HS65_LS_NOR2X6 U50 ( .A(n3), .B(n21), .Z(rdata[32]) );
  HS65_LS_NOR2AX3 U51 ( .A(rdata0[15]), .B(n3), .Z(rdata[63]) );
  HS65_LS_IVX9 U52 ( .A(rdata1[18]), .Z(n19) );
  HS65_LS_IVX9 U53 ( .A(rdata1[19]), .Z(n18) );
  HS65_LS_IVX9 U54 ( .A(rdata1[17]), .Z(n20) );
  HS65_LS_NOR2AX3 U55 ( .A(rdata0[3]), .B(n3), .Z(rdata[51]) );
  HS65_LS_NOR2AX3 U56 ( .A(rdata0[4]), .B(n4), .Z(rdata[52]) );
  HS65_LS_NOR2AX3 U57 ( .A(rdata0[7]), .B(n4), .Z(rdata[55]) );
  HS65_LS_NOR2AX3 U58 ( .A(rdata0[8]), .B(n4), .Z(rdata[56]) );
  HS65_LS_NOR2AX3 U59 ( .A(rdata0[10]), .B(n4), .Z(rdata[58]) );
  HS65_LS_NOR2AX3 U60 ( .A(rdata0[12]), .B(n4), .Z(rdata[60]) );
  HS65_LS_NOR2AX3 U61 ( .A(rdata0[1]), .B(n3), .Z(rdata[49]) );
  HS65_LS_NOR2AX3 U62 ( .A(rdata0[2]), .B(n3), .Z(rdata[50]) );
  HS65_LS_NOR2AX3 U63 ( .A(rdata0[5]), .B(n4), .Z(rdata[53]) );
  HS65_LS_NOR2AX3 U64 ( .A(rdata0[6]), .B(n4), .Z(rdata[54]) );
  HS65_LS_NOR2AX3 U65 ( .A(rdata0[9]), .B(n4), .Z(rdata[57]) );
  HS65_LS_NOR2AX3 U66 ( .A(rdata0[11]), .B(n4), .Z(rdata[59]) );
  HS65_LS_NOR2AX3 U67 ( .A(rdata0[14]), .B(n4), .Z(rdata[62]) );
  HS65_LS_OAI31X5 U68 ( .A(n44), .B(sel_out[2]), .C(sel_out[1]), .D(n2), .Z(
        n47) );
  HS65_LS_NOR3X4 U69 ( .A(sel_out[0]), .B(sel_out[1]), .C(n43), .Z(n48) );
  HS65_LS_OAI22X6 U70 ( .A(n45), .B(n9), .C(n1), .D(n25), .Z(rdata[28]) );
  HS65_LS_IVX9 U71 ( .A(rdata1[12]), .Z(n25) );
  HS65_LS_OAI22X6 U72 ( .A(n45), .B(n8), .C(n1), .D(n24), .Z(rdata[29]) );
  HS65_LS_IVX9 U73 ( .A(rdata1[13]), .Z(n24) );
  HS65_LS_OAI22X6 U74 ( .A(n45), .B(n7), .C(n1), .D(n23), .Z(rdata[30]) );
  HS65_LS_IVX9 U75 ( .A(rdata1[14]), .Z(n23) );
  HS65_LS_OAI22X6 U76 ( .A(n45), .B(n6), .C(n1), .D(n22), .Z(rdata[31]) );
  HS65_LS_IVX9 U77 ( .A(rdata1[15]), .Z(n22) );
  HS65_LS_OAI22X6 U78 ( .A(n45), .B(n21), .C(n1), .D(n41), .Z(rdata[16]) );
  HS65_LS_IVX9 U79 ( .A(rdata1[0]), .Z(n41) );
  HS65_LS_NOR2AX3 U80 ( .A(rdata0[0]), .B(n3), .Z(rdata[48]) );
  HS65_LS_IVX9 U81 ( .A(rdata1[20]), .Z(n17) );
  HS65_LS_IVX9 U82 ( .A(rdata1[21]), .Z(n16) );
  HS65_LS_IVX9 U83 ( .A(rdata1[22]), .Z(n15) );
  HS65_LS_IVX9 U84 ( .A(rdata1[23]), .Z(n14) );
  HS65_LS_IVX9 U85 ( .A(rdata1[24]), .Z(n13) );
  HS65_LS_IVX9 U86 ( .A(rdata1[25]), .Z(n12) );
  HS65_LS_IVX9 U87 ( .A(rdata1[26]), .Z(n11) );
  HS65_LS_IVX9 U88 ( .A(rdata1[27]), .Z(n10) );
  HS65_LS_IVX9 U89 ( .A(rdata1[28]), .Z(n9) );
  HS65_LS_IVX9 U90 ( .A(rdata1[29]), .Z(n8) );
  HS65_LS_IVX9 U91 ( .A(rdata1[30]), .Z(n7) );
  HS65_LS_IVX9 U92 ( .A(rdata1[31]), .Z(n6) );
  HS65_LS_IVX9 U93 ( .A(rdata1[16]), .Z(n21) );
  HS65_LS_AO222X4 U94 ( .A(rdata0[0]), .B(n48), .C(rdata1[0]), .D(n42), .E(
        rdata2[0]), .F(n47), .Z(rdata[0]) );
  HS65_LS_AO222X4 U95 ( .A(rdata0[1]), .B(n48), .C(rdata1[1]), .D(n42), .E(
        rdata2[1]), .F(n47), .Z(rdata[1]) );
  HS65_LS_AO222X4 U96 ( .A(rdata0[2]), .B(n48), .C(rdata1[2]), .D(n42), .E(
        rdata2[2]), .F(n47), .Z(rdata[2]) );
  HS65_LS_AO222X4 U97 ( .A(rdata0[3]), .B(n48), .C(rdata1[3]), .D(n42), .E(
        rdata2[3]), .F(n47), .Z(rdata[3]) );
  HS65_LS_AO222X4 U98 ( .A(rdata0[4]), .B(n48), .C(rdata1[4]), .D(n42), .E(
        rdata2[4]), .F(n47), .Z(rdata[4]) );
  HS65_LS_AO222X4 U99 ( .A(rdata0[5]), .B(n48), .C(rdata1[5]), .D(n42), .E(
        rdata2[5]), .F(n47), .Z(rdata[5]) );
  HS65_LS_AO222X4 U100 ( .A(rdata0[6]), .B(n48), .C(rdata1[6]), .D(n42), .E(
        rdata2[6]), .F(n47), .Z(rdata[6]) );
  HS65_LS_AO222X4 U101 ( .A(rdata0[7]), .B(n48), .C(rdata1[7]), .D(n42), .E(
        rdata2[7]), .F(n47), .Z(rdata[7]) );
  HS65_LS_AO222X4 U102 ( .A(rdata0[8]), .B(n48), .C(rdata1[8]), .D(n42), .E(
        rdata2[8]), .F(n47), .Z(rdata[8]) );
  HS65_LS_AO222X4 U103 ( .A(rdata0[9]), .B(n48), .C(rdata1[9]), .D(n42), .E(
        rdata2[9]), .F(n47), .Z(rdata[9]) );
  HS65_LS_AO222X4 U104 ( .A(rdata0[10]), .B(n48), .C(rdata1[10]), .D(n42), .E(
        rdata2[10]), .F(n47), .Z(rdata[10]) );
  HS65_LS_AO222X4 U105 ( .A(rdata0[11]), .B(n48), .C(rdata1[11]), .D(n42), .E(
        rdata2[11]), .F(n47), .Z(rdata[11]) );
  HS65_LS_AO222X4 U106 ( .A(rdata0[12]), .B(n48), .C(rdata1[12]), .D(n42), .E(
        rdata2[12]), .F(n47), .Z(rdata[12]) );
  HS65_LS_AO222X4 U107 ( .A(rdata0[13]), .B(n48), .C(rdata1[13]), .D(n42), .E(
        rdata2[13]), .F(n47), .Z(rdata[13]) );
  HS65_LS_AO222X4 U108 ( .A(rdata0[14]), .B(n48), .C(rdata1[14]), .D(n42), .E(
        rdata2[14]), .F(n47), .Z(rdata[14]) );
  HS65_LS_AO222X4 U109 ( .A(rdata0[15]), .B(n48), .C(rdata1[15]), .D(n42), .E(
        rdata2[15]), .F(n47), .Z(rdata[15]) );
  HS65_LS_NOR2AX3 U110 ( .A(rdata0[13]), .B(n4), .Z(rdata[61]) );
endmodule


module bram_DATA5_ADDR3_3 ( clk, reset, rd_addr, wr_addr, wr_data, wr_ena, 
        rd_data );
  input [2:0] rd_addr;
  input [2:0] wr_addr;
  input [4:0] wr_data;
  output [4:0] rd_data;
  input clk, reset, wr_ena;
  wire   \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N34,
         N35, N36, N37, N38, n1, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218;

  HS65_LS_DFPRQX9 \mem_reg[5][4]  ( .D(n131), .CP(clk), .RN(n1), .Q(
        \mem[5][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[5][3]  ( .D(n132), .CP(clk), .RN(n1), .Q(
        \mem[5][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[5][2]  ( .D(n133), .CP(clk), .RN(n1), .Q(
        \mem[5][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[5][1]  ( .D(n134), .CP(clk), .RN(n1), .Q(
        \mem[5][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[5][0]  ( .D(n135), .CP(clk), .RN(n22), .Q(
        \mem[5][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[4][4]  ( .D(n136), .CP(clk), .RN(n22), .Q(
        \mem[4][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[4][3]  ( .D(n137), .CP(clk), .RN(n22), .Q(
        \mem[4][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[4][2]  ( .D(n138), .CP(clk), .RN(n22), .Q(
        \mem[4][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[4][1]  ( .D(n139), .CP(clk), .RN(n22), .Q(
        \mem[4][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[4][0]  ( .D(n140), .CP(clk), .RN(n22), .Q(
        \mem[4][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][4]  ( .D(n151), .CP(clk), .RN(n22), .Q(
        \mem[1][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][3]  ( .D(n152), .CP(clk), .RN(n22), .Q(
        \mem[1][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][2]  ( .D(n153), .CP(clk), .RN(n22), .Q(
        \mem[1][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][1]  ( .D(n154), .CP(clk), .RN(n22), .Q(
        \mem[1][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][0]  ( .D(n155), .CP(clk), .RN(n22), .Q(
        \mem[1][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][4]  ( .D(n156), .CP(clk), .RN(n22), .Q(
        \mem[0][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][3]  ( .D(n157), .CP(clk), .RN(n1), .Q(
        \mem[0][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][2]  ( .D(n158), .CP(clk), .RN(n1), .Q(
        \mem[0][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][1]  ( .D(n159), .CP(clk), .RN(n1), .Q(
        \mem[0][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][0]  ( .D(n160), .CP(clk), .RN(n1), .Q(
        \mem[0][0] ) );
  HS65_LS_DFPRQX9 \rd_data_reg[4]  ( .D(N34), .CP(clk), .RN(n1), .Q(rd_data[4]) );
  HS65_LS_DFPRQX9 \rd_data_reg[3]  ( .D(N35), .CP(clk), .RN(n1), .Q(rd_data[3]) );
  HS65_LS_DFPRQX9 \rd_data_reg[2]  ( .D(N36), .CP(clk), .RN(n1), .Q(rd_data[2]) );
  HS65_LS_DFPRQX9 \rd_data_reg[1]  ( .D(N37), .CP(clk), .RN(n1), .Q(rd_data[1]) );
  HS65_LS_DFPRQX9 \rd_data_reg[0]  ( .D(N38), .CP(clk), .RN(n1), .Q(rd_data[0]) );
  HS65_LS_DFPRQNX9 \mem_reg[7][4]  ( .D(n121), .CP(clk), .RN(n23), .QN(n218)
         );
  HS65_LS_DFPRQNX9 \mem_reg[7][3]  ( .D(n122), .CP(clk), .RN(n22), .QN(n217)
         );
  HS65_LS_DFPRQNX9 \mem_reg[7][2]  ( .D(n123), .CP(clk), .RN(n24), .QN(n216)
         );
  HS65_LS_DFPRQNX9 \mem_reg[7][1]  ( .D(n124), .CP(clk), .RN(n24), .QN(n215)
         );
  HS65_LS_DFPRQNX9 \mem_reg[7][0]  ( .D(n125), .CP(clk), .RN(n24), .QN(n214)
         );
  HS65_LS_DFPRQNX9 \mem_reg[3][4]  ( .D(n141), .CP(clk), .RN(n23), .QN(n208)
         );
  HS65_LS_DFPRQNX9 \mem_reg[3][3]  ( .D(n142), .CP(clk), .RN(n23), .QN(n207)
         );
  HS65_LS_DFPRQNX9 \mem_reg[3][2]  ( .D(n143), .CP(clk), .RN(n23), .QN(n206)
         );
  HS65_LS_DFPRQNX9 \mem_reg[3][1]  ( .D(n144), .CP(clk), .RN(n23), .QN(n205)
         );
  HS65_LS_DFPRQNX9 \mem_reg[3][0]  ( .D(n145), .CP(clk), .RN(n23), .QN(n204)
         );
  HS65_LS_DFPRQNX9 \mem_reg[6][4]  ( .D(n126), .CP(clk), .RN(n24), .QN(n213)
         );
  HS65_LS_DFPRQNX9 \mem_reg[6][3]  ( .D(n127), .CP(clk), .RN(n24), .QN(n212)
         );
  HS65_LS_DFPRQNX9 \mem_reg[6][2]  ( .D(n128), .CP(clk), .RN(n23), .QN(n211)
         );
  HS65_LS_DFPRQNX9 \mem_reg[6][1]  ( .D(n129), .CP(clk), .RN(n23), .QN(n210)
         );
  HS65_LS_DFPRQNX9 \mem_reg[6][0]  ( .D(n130), .CP(clk), .RN(n23), .QN(n209)
         );
  HS65_LS_DFPRQNX9 \mem_reg[2][4]  ( .D(n146), .CP(clk), .RN(n23), .QN(n203)
         );
  HS65_LS_DFPRQNX9 \mem_reg[2][3]  ( .D(n147), .CP(clk), .RN(n23), .QN(n202)
         );
  HS65_LS_DFPRQNX9 \mem_reg[2][2]  ( .D(n148), .CP(clk), .RN(n23), .QN(n201)
         );
  HS65_LS_DFPRQNX9 \mem_reg[2][1]  ( .D(n149), .CP(clk), .RN(n23), .QN(n200)
         );
  HS65_LS_DFPRQNX9 \mem_reg[2][0]  ( .D(n150), .CP(clk), .RN(n23), .QN(n199)
         );
  HS65_LS_BFX9 U3 ( .A(n25), .Z(n1) );
  HS65_LS_BFX9 U4 ( .A(n25), .Z(n22) );
  HS65_LS_BFX9 U5 ( .A(n25), .Z(n23) );
  HS65_LS_BFX9 U6 ( .A(n25), .Z(n24) );
  HS65_LS_IVX9 U7 ( .A(reset), .Z(n25) );
  HS65_LS_IVX9 U8 ( .A(n198), .Z(n35) );
  HS65_LS_IVX9 U9 ( .A(n193), .Z(n31) );
  HS65_LS_IVX9 U10 ( .A(n194), .Z(n32) );
  HS65_LS_IVX9 U11 ( .A(n190), .Z(n29) );
  HS65_LS_IVX9 U12 ( .A(n189), .Z(n28) );
  HS65_LS_IVX9 U13 ( .A(n195), .Z(n33) );
  HS65_LS_NAND3X5 U14 ( .A(n37), .B(n36), .C(n197), .Z(n198) );
  HS65_LS_NAND3X5 U15 ( .A(n37), .B(n36), .C(n192), .Z(n193) );
  HS65_LS_IVX9 U16 ( .A(n191), .Z(n30) );
  HS65_LS_IVX9 U17 ( .A(n196), .Z(n34) );
  HS65_LS_NOR3X4 U18 ( .A(n26), .B(rd_addr[1]), .C(n27), .Z(n186) );
  HS65_LS_NOR3X4 U19 ( .A(rd_addr[1]), .B(rd_addr[2]), .C(n26), .Z(n181) );
  HS65_LS_NOR3X4 U20 ( .A(rd_addr[1]), .B(rd_addr[2]), .C(rd_addr[0]), .Z(n180) );
  HS65_LS_NOR3X4 U21 ( .A(rd_addr[0]), .B(rd_addr[1]), .C(n27), .Z(n185) );
  HS65_LS_NAND3X5 U22 ( .A(n26), .B(n27), .C(rd_addr[1]), .Z(n178) );
  HS65_LS_NAND3X5 U23 ( .A(rd_addr[0]), .B(n27), .C(rd_addr[1]), .Z(n177) );
  HS65_LS_NAND3X5 U24 ( .A(rd_addr[1]), .B(n26), .C(rd_addr[2]), .Z(n183) );
  HS65_LS_NAND3X5 U25 ( .A(rd_addr[1]), .B(rd_addr[0]), .C(rd_addr[2]), .Z(
        n182) );
  HS65_LS_OAI22X6 U26 ( .A(n199), .B(n178), .C(n204), .D(n177), .Z(n179) );
  HS65_LS_OAI22X6 U27 ( .A(n200), .B(n178), .C(n205), .D(n177), .Z(n173) );
  HS65_LS_OAI22X6 U28 ( .A(n201), .B(n178), .C(n206), .D(n177), .Z(n169) );
  HS65_LS_OAI22X6 U29 ( .A(n202), .B(n178), .C(n207), .D(n177), .Z(n165) );
  HS65_LS_OAI22X6 U30 ( .A(n203), .B(n178), .C(n208), .D(n177), .Z(n161) );
  HS65_LS_IVX9 U31 ( .A(rd_addr[0]), .Z(n26) );
  HS65_LS_IVX9 U32 ( .A(rd_addr[2]), .Z(n27) );
  HS65_LS_OAI22X6 U33 ( .A(n120), .B(n194), .C(n32), .D(n204), .Z(n145) );
  HS65_LS_OAI22X6 U34 ( .A(n119), .B(n194), .C(n32), .D(n205), .Z(n144) );
  HS65_LS_OAI22X6 U35 ( .A(n118), .B(n194), .C(n32), .D(n206), .Z(n143) );
  HS65_LS_OAI22X6 U36 ( .A(n117), .B(n194), .C(n32), .D(n207), .Z(n142) );
  HS65_LS_OAI22X6 U37 ( .A(n38), .B(n194), .C(n32), .D(n208), .Z(n141) );
  HS65_LS_OAI22X6 U38 ( .A(n120), .B(n190), .C(n29), .D(n209), .Z(n130) );
  HS65_LS_OAI22X6 U39 ( .A(n119), .B(n190), .C(n29), .D(n210), .Z(n129) );
  HS65_LS_OAI22X6 U40 ( .A(n118), .B(n190), .C(n29), .D(n211), .Z(n128) );
  HS65_LS_OAI22X6 U41 ( .A(n117), .B(n190), .C(n29), .D(n212), .Z(n127) );
  HS65_LS_OAI22X6 U42 ( .A(n38), .B(n190), .C(n29), .D(n213), .Z(n126) );
  HS65_LS_OAI22X6 U43 ( .A(n120), .B(n189), .C(n28), .D(n214), .Z(n125) );
  HS65_LS_OAI22X6 U44 ( .A(n119), .B(n189), .C(n28), .D(n215), .Z(n124) );
  HS65_LS_OAI22X6 U45 ( .A(n118), .B(n189), .C(n28), .D(n216), .Z(n123) );
  HS65_LS_OAI22X6 U46 ( .A(n117), .B(n189), .C(n28), .D(n217), .Z(n122) );
  HS65_LS_OAI22X6 U47 ( .A(n38), .B(n189), .C(n28), .D(n218), .Z(n121) );
  HS65_LS_OAI22X6 U48 ( .A(n120), .B(n195), .C(n33), .D(n199), .Z(n150) );
  HS65_LS_OAI22X6 U49 ( .A(n119), .B(n195), .C(n33), .D(n200), .Z(n149) );
  HS65_LS_OAI22X6 U50 ( .A(n118), .B(n195), .C(n33), .D(n201), .Z(n148) );
  HS65_LS_OAI22X6 U51 ( .A(n117), .B(n195), .C(n33), .D(n202), .Z(n147) );
  HS65_LS_OAI22X6 U52 ( .A(n38), .B(n195), .C(n33), .D(n203), .Z(n146) );
  HS65_LS_NAND2X7 U53 ( .A(n188), .B(n187), .Z(N38) );
  HS65_LS_AOI212X4 U54 ( .A(n186), .B(\mem[5][0] ), .C(n185), .D(\mem[4][0] ), 
        .E(n184), .Z(n187) );
  HS65_LS_AOI212X4 U55 ( .A(n181), .B(\mem[1][0] ), .C(n180), .D(\mem[0][0] ), 
        .E(n179), .Z(n188) );
  HS65_LS_OAI22X6 U56 ( .A(n209), .B(n183), .C(n214), .D(n182), .Z(n184) );
  HS65_LS_NAND2X7 U57 ( .A(n176), .B(n175), .Z(N37) );
  HS65_LS_AOI212X4 U58 ( .A(n186), .B(\mem[5][1] ), .C(n185), .D(\mem[4][1] ), 
        .E(n174), .Z(n175) );
  HS65_LS_AOI212X4 U59 ( .A(n181), .B(\mem[1][1] ), .C(n180), .D(\mem[0][1] ), 
        .E(n173), .Z(n176) );
  HS65_LS_OAI22X6 U60 ( .A(n210), .B(n183), .C(n215), .D(n182), .Z(n174) );
  HS65_LS_NAND2X7 U61 ( .A(n172), .B(n171), .Z(N36) );
  HS65_LS_AOI212X4 U62 ( .A(n186), .B(\mem[5][2] ), .C(n185), .D(\mem[4][2] ), 
        .E(n170), .Z(n171) );
  HS65_LS_AOI212X4 U63 ( .A(n181), .B(\mem[1][2] ), .C(n180), .D(\mem[0][2] ), 
        .E(n169), .Z(n172) );
  HS65_LS_OAI22X6 U64 ( .A(n211), .B(n183), .C(n216), .D(n182), .Z(n170) );
  HS65_LS_NAND2X7 U65 ( .A(n168), .B(n167), .Z(N35) );
  HS65_LS_AOI212X4 U66 ( .A(n186), .B(\mem[5][3] ), .C(n185), .D(\mem[4][3] ), 
        .E(n166), .Z(n167) );
  HS65_LS_AOI212X4 U67 ( .A(n181), .B(\mem[1][3] ), .C(n180), .D(\mem[0][3] ), 
        .E(n165), .Z(n168) );
  HS65_LS_OAI22X6 U68 ( .A(n212), .B(n183), .C(n217), .D(n182), .Z(n166) );
  HS65_LS_NAND2X7 U69 ( .A(n164), .B(n163), .Z(N34) );
  HS65_LS_AOI212X4 U70 ( .A(n186), .B(\mem[5][4] ), .C(n185), .D(\mem[4][4] ), 
        .E(n162), .Z(n163) );
  HS65_LS_AOI212X4 U71 ( .A(n181), .B(\mem[1][4] ), .C(n180), .D(\mem[0][4] ), 
        .E(n161), .Z(n164) );
  HS65_LS_OAI22X6 U72 ( .A(n213), .B(n183), .C(n218), .D(n182), .Z(n162) );
  HS65_LS_AO22X9 U73 ( .A(n35), .B(wr_data[0]), .C(n198), .D(\mem[0][0] ), .Z(
        n160) );
  HS65_LS_AO22X9 U74 ( .A(n35), .B(wr_data[1]), .C(n198), .D(\mem[0][1] ), .Z(
        n159) );
  HS65_LS_AO22X9 U75 ( .A(n35), .B(wr_data[2]), .C(n198), .D(\mem[0][2] ), .Z(
        n158) );
  HS65_LS_AO22X9 U76 ( .A(n35), .B(wr_data[3]), .C(n198), .D(\mem[0][3] ), .Z(
        n157) );
  HS65_LS_AO22X9 U77 ( .A(n35), .B(wr_data[4]), .C(n198), .D(\mem[0][4] ), .Z(
        n156) );
  HS65_LS_AO22X9 U78 ( .A(wr_data[0]), .B(n31), .C(n193), .D(\mem[4][0] ), .Z(
        n140) );
  HS65_LS_AO22X9 U79 ( .A(wr_data[1]), .B(n31), .C(n193), .D(\mem[4][1] ), .Z(
        n139) );
  HS65_LS_AO22X9 U80 ( .A(wr_data[2]), .B(n31), .C(n193), .D(\mem[4][2] ), .Z(
        n138) );
  HS65_LS_AO22X9 U81 ( .A(wr_data[3]), .B(n31), .C(n193), .D(\mem[4][3] ), .Z(
        n137) );
  HS65_LS_AO22X9 U82 ( .A(wr_data[4]), .B(n31), .C(n193), .D(\mem[4][4] ), .Z(
        n136) );
  HS65_LS_AO22X9 U83 ( .A(wr_data[0]), .B(n30), .C(n191), .D(\mem[5][0] ), .Z(
        n135) );
  HS65_LS_AO22X9 U84 ( .A(wr_data[1]), .B(n30), .C(n191), .D(\mem[5][1] ), .Z(
        n134) );
  HS65_LS_AO22X9 U85 ( .A(wr_data[2]), .B(n30), .C(n191), .D(\mem[5][2] ), .Z(
        n133) );
  HS65_LS_AO22X9 U86 ( .A(wr_data[3]), .B(n30), .C(n191), .D(\mem[5][3] ), .Z(
        n132) );
  HS65_LS_AO22X9 U87 ( .A(wr_data[4]), .B(n30), .C(n191), .D(\mem[5][4] ), .Z(
        n131) );
  HS65_LS_AO22X9 U88 ( .A(wr_data[0]), .B(n34), .C(n196), .D(\mem[1][0] ), .Z(
        n155) );
  HS65_LS_AO22X9 U89 ( .A(wr_data[1]), .B(n34), .C(n196), .D(\mem[1][1] ), .Z(
        n154) );
  HS65_LS_AO22X9 U90 ( .A(wr_data[2]), .B(n34), .C(n196), .D(\mem[1][2] ), .Z(
        n153) );
  HS65_LS_AO22X9 U91 ( .A(wr_data[3]), .B(n34), .C(n196), .D(\mem[1][3] ), .Z(
        n152) );
  HS65_LS_AO22X9 U92 ( .A(wr_data[4]), .B(n34), .C(n196), .D(\mem[1][4] ), .Z(
        n151) );
  HS65_LS_NAND3X5 U93 ( .A(wr_addr[0]), .B(n197), .C(wr_addr[1]), .Z(n194) );
  HS65_LS_NAND3X5 U94 ( .A(wr_addr[1]), .B(n37), .C(n192), .Z(n190) );
  HS65_LS_NAND3X5 U95 ( .A(wr_addr[1]), .B(wr_addr[0]), .C(n192), .Z(n189) );
  HS65_LS_NAND3X5 U96 ( .A(n197), .B(n37), .C(wr_addr[1]), .Z(n195) );
  HS65_LS_NOR2AX3 U97 ( .A(wr_ena), .B(wr_addr[2]), .Z(n197) );
  HS65_LS_NAND3X5 U98 ( .A(wr_addr[0]), .B(n36), .C(n192), .Z(n191) );
  HS65_LS_NAND3X5 U99 ( .A(n197), .B(n36), .C(wr_addr[0]), .Z(n196) );
  HS65_LS_IVX9 U100 ( .A(wr_addr[0]), .Z(n37) );
  HS65_LS_IVX9 U101 ( .A(wr_data[0]), .Z(n120) );
  HS65_LS_IVX9 U102 ( .A(wr_data[1]), .Z(n119) );
  HS65_LS_IVX9 U103 ( .A(wr_data[2]), .Z(n118) );
  HS65_LS_IVX9 U104 ( .A(wr_data[3]), .Z(n117) );
  HS65_LS_IVX9 U105 ( .A(wr_data[4]), .Z(n38) );
  HS65_LS_IVX9 U106 ( .A(wr_addr[1]), .Z(n36) );
  HS65_LS_AND2X4 U107 ( .A(wr_addr[2]), .B(wr_ena), .Z(n192) );
endmodule


module nAdapter_3 ( na_clk, na_reset, .proc_in({\proc_in[MCMD][1] , 
        \proc_in[MCMD][0] , \proc_in[MADDR][31] , \proc_in[MADDR][30] , 
        \proc_in[MADDR][29] , \proc_in[MADDR][28] , \proc_in[MADDR][27] , 
        \proc_in[MADDR][26] , \proc_in[MADDR][25] , \proc_in[MADDR][24] , 
        \proc_in[MADDR][23] , \proc_in[MADDR][22] , \proc_in[MADDR][21] , 
        \proc_in[MADDR][20] , \proc_in[MADDR][19] , \proc_in[MADDR][18] , 
        \proc_in[MADDR][17] , \proc_in[MADDR][16] , \proc_in[MADDR][15] , 
        \proc_in[MADDR][14] , \proc_in[MADDR][13] , \proc_in[MADDR][12] , 
        \proc_in[MADDR][11] , \proc_in[MADDR][10] , \proc_in[MADDR][9] , 
        \proc_in[MADDR][8] , \proc_in[MADDR][7] , \proc_in[MADDR][6] , 
        \proc_in[MADDR][5] , \proc_in[MADDR][4] , \proc_in[MADDR][3] , 
        \proc_in[MADDR][2] , \proc_in[MADDR][1] , \proc_in[MADDR][0] , 
        \proc_in[MDATA][31] , \proc_in[MDATA][30] , \proc_in[MDATA][29] , 
        \proc_in[MDATA][28] , \proc_in[MDATA][27] , \proc_in[MDATA][26] , 
        \proc_in[MDATA][25] , \proc_in[MDATA][24] , \proc_in[MDATA][23] , 
        \proc_in[MDATA][22] , \proc_in[MDATA][21] , \proc_in[MDATA][20] , 
        \proc_in[MDATA][19] , \proc_in[MDATA][18] , \proc_in[MDATA][17] , 
        \proc_in[MDATA][16] , \proc_in[MDATA][15] , \proc_in[MDATA][14] , 
        \proc_in[MDATA][13] , \proc_in[MDATA][12] , \proc_in[MDATA][11] , 
        \proc_in[MDATA][10] , \proc_in[MDATA][9] , \proc_in[MDATA][8] , 
        \proc_in[MDATA][7] , \proc_in[MDATA][6] , \proc_in[MDATA][5] , 
        \proc_in[MDATA][4] , \proc_in[MDATA][3] , \proc_in[MDATA][2] , 
        \proc_in[MDATA][1] , \proc_in[MDATA][0] }), .proc_out({
        \proc_out[SCMDACCEPT] , \proc_out[SRESP] , \proc_out[SDATA][31] , 
        \proc_out[SDATA][30] , \proc_out[SDATA][29] , \proc_out[SDATA][28] , 
        \proc_out[SDATA][27] , \proc_out[SDATA][26] , \proc_out[SDATA][25] , 
        \proc_out[SDATA][24] , \proc_out[SDATA][23] , \proc_out[SDATA][22] , 
        \proc_out[SDATA][21] , \proc_out[SDATA][20] , \proc_out[SDATA][19] , 
        \proc_out[SDATA][18] , \proc_out[SDATA][17] , \proc_out[SDATA][16] , 
        \proc_out[SDATA][15] , \proc_out[SDATA][14] , \proc_out[SDATA][13] , 
        \proc_out[SDATA][12] , \proc_out[SDATA][11] , \proc_out[SDATA][10] , 
        \proc_out[SDATA][9] , \proc_out[SDATA][8] , \proc_out[SDATA][7] , 
        \proc_out[SDATA][6] , \proc_out[SDATA][5] , \proc_out[SDATA][4] , 
        \proc_out[SDATA][3] , \proc_out[SDATA][2] , \proc_out[SDATA][1] , 
        \proc_out[SDATA][0] }), .spm_in({\spm_in[SCMDACCEPT] , \spm_in[SRESP] , 
        \spm_in[SDATA][63] , \spm_in[SDATA][62] , \spm_in[SDATA][61] , 
        \spm_in[SDATA][60] , \spm_in[SDATA][59] , \spm_in[SDATA][58] , 
        \spm_in[SDATA][57] , \spm_in[SDATA][56] , \spm_in[SDATA][55] , 
        \spm_in[SDATA][54] , \spm_in[SDATA][53] , \spm_in[SDATA][52] , 
        \spm_in[SDATA][51] , \spm_in[SDATA][50] , \spm_in[SDATA][49] , 
        \spm_in[SDATA][48] , \spm_in[SDATA][47] , \spm_in[SDATA][46] , 
        \spm_in[SDATA][45] , \spm_in[SDATA][44] , \spm_in[SDATA][43] , 
        \spm_in[SDATA][42] , \spm_in[SDATA][41] , \spm_in[SDATA][40] , 
        \spm_in[SDATA][39] , \spm_in[SDATA][38] , \spm_in[SDATA][37] , 
        \spm_in[SDATA][36] , \spm_in[SDATA][35] , \spm_in[SDATA][34] , 
        \spm_in[SDATA][33] , \spm_in[SDATA][32] , \spm_in[SDATA][31] , 
        \spm_in[SDATA][30] , \spm_in[SDATA][29] , \spm_in[SDATA][28] , 
        \spm_in[SDATA][27] , \spm_in[SDATA][26] , \spm_in[SDATA][25] , 
        \spm_in[SDATA][24] , \spm_in[SDATA][23] , \spm_in[SDATA][22] , 
        \spm_in[SDATA][21] , \spm_in[SDATA][20] , \spm_in[SDATA][19] , 
        \spm_in[SDATA][18] , \spm_in[SDATA][17] , \spm_in[SDATA][16] , 
        \spm_in[SDATA][15] , \spm_in[SDATA][14] , \spm_in[SDATA][13] , 
        \spm_in[SDATA][12] , \spm_in[SDATA][11] , \spm_in[SDATA][10] , 
        \spm_in[SDATA][9] , \spm_in[SDATA][8] , \spm_in[SDATA][7] , 
        \spm_in[SDATA][6] , \spm_in[SDATA][5] , \spm_in[SDATA][4] , 
        \spm_in[SDATA][3] , \spm_in[SDATA][2] , \spm_in[SDATA][1] , 
        \spm_in[SDATA][0] }), .spm_out({\spm_out[MCMD][1] , \spm_out[MCMD][0] , 
        \spm_out[MADDR][31] , \spm_out[MADDR][30] , \spm_out[MADDR][29] , 
        \spm_out[MADDR][28] , \spm_out[MADDR][27] , \spm_out[MADDR][26] , 
        \spm_out[MADDR][25] , \spm_out[MADDR][24] , \spm_out[MADDR][23] , 
        \spm_out[MADDR][22] , \spm_out[MADDR][21] , \spm_out[MADDR][20] , 
        \spm_out[MADDR][19] , \spm_out[MADDR][18] , \spm_out[MADDR][17] , 
        \spm_out[MADDR][16] , \spm_out[MADDR][15] , \spm_out[MADDR][14] , 
        \spm_out[MADDR][13] , \spm_out[MADDR][12] , \spm_out[MADDR][11] , 
        \spm_out[MADDR][10] , \spm_out[MADDR][9] , \spm_out[MADDR][8] , 
        \spm_out[MADDR][7] , \spm_out[MADDR][6] , \spm_out[MADDR][5] , 
        \spm_out[MADDR][4] , \spm_out[MADDR][3] , \spm_out[MADDR][2] , 
        \spm_out[MADDR][1] , \spm_out[MADDR][0] , \spm_out[MDATA][63] , 
        \spm_out[MDATA][62] , \spm_out[MDATA][61] , \spm_out[MDATA][60] , 
        \spm_out[MDATA][59] , \spm_out[MDATA][58] , \spm_out[MDATA][57] , 
        \spm_out[MDATA][56] , \spm_out[MDATA][55] , \spm_out[MDATA][54] , 
        \spm_out[MDATA][53] , \spm_out[MDATA][52] , \spm_out[MDATA][51] , 
        \spm_out[MDATA][50] , \spm_out[MDATA][49] , \spm_out[MDATA][48] , 
        \spm_out[MDATA][47] , \spm_out[MDATA][46] , \spm_out[MDATA][45] , 
        \spm_out[MDATA][44] , \spm_out[MDATA][43] , \spm_out[MDATA][42] , 
        \spm_out[MDATA][41] , \spm_out[MDATA][40] , \spm_out[MDATA][39] , 
        \spm_out[MDATA][38] , \spm_out[MDATA][37] , \spm_out[MDATA][36] , 
        \spm_out[MDATA][35] , \spm_out[MDATA][34] , \spm_out[MDATA][33] , 
        \spm_out[MDATA][32] , \spm_out[MDATA][31] , \spm_out[MDATA][30] , 
        \spm_out[MDATA][29] , \spm_out[MDATA][28] , \spm_out[MDATA][27] , 
        \spm_out[MDATA][26] , \spm_out[MDATA][25] , \spm_out[MDATA][24] , 
        \spm_out[MDATA][23] , \spm_out[MDATA][22] , \spm_out[MDATA][21] , 
        \spm_out[MDATA][20] , \spm_out[MDATA][19] , \spm_out[MDATA][18] , 
        \spm_out[MDATA][17] , \spm_out[MDATA][16] , \spm_out[MDATA][15] , 
        \spm_out[MDATA][14] , \spm_out[MDATA][13] , \spm_out[MDATA][12] , 
        \spm_out[MDATA][11] , \spm_out[MDATA][10] , \spm_out[MDATA][9] , 
        \spm_out[MDATA][8] , \spm_out[MDATA][7] , \spm_out[MDATA][6] , 
        \spm_out[MDATA][5] , \spm_out[MDATA][4] , \spm_out[MDATA][3] , 
        \spm_out[MDATA][2] , \spm_out[MDATA][1] , \spm_out[MDATA][0] }), 
        pkt_in, pkt_out );
  input [34:0] pkt_in;
  output [34:0] pkt_out;
  input na_clk, na_reset, \proc_in[MCMD][1] , \proc_in[MCMD][0] ,
         \proc_in[MADDR][31] , \proc_in[MADDR][30] , \proc_in[MADDR][29] ,
         \proc_in[MADDR][28] , \proc_in[MADDR][27] , \proc_in[MADDR][26] ,
         \proc_in[MADDR][25] , \proc_in[MADDR][24] , \proc_in[MADDR][23] ,
         \proc_in[MADDR][22] , \proc_in[MADDR][21] , \proc_in[MADDR][20] ,
         \proc_in[MADDR][19] , \proc_in[MADDR][18] , \proc_in[MADDR][17] ,
         \proc_in[MADDR][16] , \proc_in[MADDR][15] , \proc_in[MADDR][14] ,
         \proc_in[MADDR][13] , \proc_in[MADDR][12] , \proc_in[MADDR][11] ,
         \proc_in[MADDR][10] , \proc_in[MADDR][9] , \proc_in[MADDR][8] ,
         \proc_in[MADDR][7] , \proc_in[MADDR][6] , \proc_in[MADDR][5] ,
         \proc_in[MADDR][4] , \proc_in[MADDR][3] , \proc_in[MADDR][2] ,
         \proc_in[MADDR][1] , \proc_in[MADDR][0] , \proc_in[MDATA][31] ,
         \proc_in[MDATA][30] , \proc_in[MDATA][29] , \proc_in[MDATA][28] ,
         \proc_in[MDATA][27] , \proc_in[MDATA][26] , \proc_in[MDATA][25] ,
         \proc_in[MDATA][24] , \proc_in[MDATA][23] , \proc_in[MDATA][22] ,
         \proc_in[MDATA][21] , \proc_in[MDATA][20] , \proc_in[MDATA][19] ,
         \proc_in[MDATA][18] , \proc_in[MDATA][17] , \proc_in[MDATA][16] ,
         \proc_in[MDATA][15] , \proc_in[MDATA][14] , \proc_in[MDATA][13] ,
         \proc_in[MDATA][12] , \proc_in[MDATA][11] , \proc_in[MDATA][10] ,
         \proc_in[MDATA][9] , \proc_in[MDATA][8] , \proc_in[MDATA][7] ,
         \proc_in[MDATA][6] , \proc_in[MDATA][5] , \proc_in[MDATA][4] ,
         \proc_in[MDATA][3] , \proc_in[MDATA][2] , \proc_in[MDATA][1] ,
         \proc_in[MDATA][0] , \spm_in[SCMDACCEPT] , \spm_in[SRESP] ,
         \spm_in[SDATA][63] , \spm_in[SDATA][62] , \spm_in[SDATA][61] ,
         \spm_in[SDATA][60] , \spm_in[SDATA][59] , \spm_in[SDATA][58] ,
         \spm_in[SDATA][57] , \spm_in[SDATA][56] , \spm_in[SDATA][55] ,
         \spm_in[SDATA][54] , \spm_in[SDATA][53] , \spm_in[SDATA][52] ,
         \spm_in[SDATA][51] , \spm_in[SDATA][50] , \spm_in[SDATA][49] ,
         \spm_in[SDATA][48] , \spm_in[SDATA][47] , \spm_in[SDATA][46] ,
         \spm_in[SDATA][45] , \spm_in[SDATA][44] , \spm_in[SDATA][43] ,
         \spm_in[SDATA][42] , \spm_in[SDATA][41] , \spm_in[SDATA][40] ,
         \spm_in[SDATA][39] , \spm_in[SDATA][38] , \spm_in[SDATA][37] ,
         \spm_in[SDATA][36] , \spm_in[SDATA][35] , \spm_in[SDATA][34] ,
         \spm_in[SDATA][33] , \spm_in[SDATA][32] , \spm_in[SDATA][31] ,
         \spm_in[SDATA][30] , \spm_in[SDATA][29] , \spm_in[SDATA][28] ,
         \spm_in[SDATA][27] , \spm_in[SDATA][26] , \spm_in[SDATA][25] ,
         \spm_in[SDATA][24] , \spm_in[SDATA][23] , \spm_in[SDATA][22] ,
         \spm_in[SDATA][21] , \spm_in[SDATA][20] , \spm_in[SDATA][19] ,
         \spm_in[SDATA][18] , \spm_in[SDATA][17] , \spm_in[SDATA][16] ,
         \spm_in[SDATA][15] , \spm_in[SDATA][14] , \spm_in[SDATA][13] ,
         \spm_in[SDATA][12] , \spm_in[SDATA][11] , \spm_in[SDATA][10] ,
         \spm_in[SDATA][9] , \spm_in[SDATA][8] , \spm_in[SDATA][7] ,
         \spm_in[SDATA][6] , \spm_in[SDATA][5] , \spm_in[SDATA][4] ,
         \spm_in[SDATA][3] , \spm_in[SDATA][2] , \spm_in[SDATA][1] ,
         \spm_in[SDATA][0] ;
  output \proc_out[SCMDACCEPT] , \proc_out[SRESP] , \proc_out[SDATA][31] ,
         \proc_out[SDATA][30] , \proc_out[SDATA][29] , \proc_out[SDATA][28] ,
         \proc_out[SDATA][27] , \proc_out[SDATA][26] , \proc_out[SDATA][25] ,
         \proc_out[SDATA][24] , \proc_out[SDATA][23] , \proc_out[SDATA][22] ,
         \proc_out[SDATA][21] , \proc_out[SDATA][20] , \proc_out[SDATA][19] ,
         \proc_out[SDATA][18] , \proc_out[SDATA][17] , \proc_out[SDATA][16] ,
         \proc_out[SDATA][15] , \proc_out[SDATA][14] , \proc_out[SDATA][13] ,
         \proc_out[SDATA][12] , \proc_out[SDATA][11] , \proc_out[SDATA][10] ,
         \proc_out[SDATA][9] , \proc_out[SDATA][8] , \proc_out[SDATA][7] ,
         \proc_out[SDATA][6] , \proc_out[SDATA][5] , \proc_out[SDATA][4] ,
         \proc_out[SDATA][3] , \proc_out[SDATA][2] , \proc_out[SDATA][1] ,
         \proc_out[SDATA][0] , \spm_out[MCMD][1] , \spm_out[MCMD][0] ,
         \spm_out[MADDR][31] , \spm_out[MADDR][30] , \spm_out[MADDR][29] ,
         \spm_out[MADDR][28] , \spm_out[MADDR][27] , \spm_out[MADDR][26] ,
         \spm_out[MADDR][25] , \spm_out[MADDR][24] , \spm_out[MADDR][23] ,
         \spm_out[MADDR][22] , \spm_out[MADDR][21] , \spm_out[MADDR][20] ,
         \spm_out[MADDR][19] , \spm_out[MADDR][18] , \spm_out[MADDR][17] ,
         \spm_out[MADDR][16] , \spm_out[MADDR][15] , \spm_out[MADDR][14] ,
         \spm_out[MADDR][13] , \spm_out[MADDR][12] , \spm_out[MADDR][11] ,
         \spm_out[MADDR][10] , \spm_out[MADDR][9] , \spm_out[MADDR][8] ,
         \spm_out[MADDR][7] , \spm_out[MADDR][6] , \spm_out[MADDR][5] ,
         \spm_out[MADDR][4] , \spm_out[MADDR][3] , \spm_out[MADDR][2] ,
         \spm_out[MADDR][1] , \spm_out[MADDR][0] , \spm_out[MDATA][63] ,
         \spm_out[MDATA][62] , \spm_out[MDATA][61] , \spm_out[MDATA][60] ,
         \spm_out[MDATA][59] , \spm_out[MDATA][58] , \spm_out[MDATA][57] ,
         \spm_out[MDATA][56] , \spm_out[MDATA][55] , \spm_out[MDATA][54] ,
         \spm_out[MDATA][53] , \spm_out[MDATA][52] , \spm_out[MDATA][51] ,
         \spm_out[MDATA][50] , \spm_out[MDATA][49] , \spm_out[MDATA][48] ,
         \spm_out[MDATA][47] , \spm_out[MDATA][46] , \spm_out[MDATA][45] ,
         \spm_out[MDATA][44] , \spm_out[MDATA][43] , \spm_out[MDATA][42] ,
         \spm_out[MDATA][41] , \spm_out[MDATA][40] , \spm_out[MDATA][39] ,
         \spm_out[MDATA][38] , \spm_out[MDATA][37] , \spm_out[MDATA][36] ,
         \spm_out[MDATA][35] , \spm_out[MDATA][34] , \spm_out[MDATA][33] ,
         \spm_out[MDATA][32] , \spm_out[MDATA][31] , \spm_out[MDATA][30] ,
         \spm_out[MDATA][29] , \spm_out[MDATA][28] , \spm_out[MDATA][27] ,
         \spm_out[MDATA][26] , \spm_out[MDATA][25] , \spm_out[MDATA][24] ,
         \spm_out[MDATA][23] , \spm_out[MDATA][22] , \spm_out[MDATA][21] ,
         \spm_out[MDATA][20] , \spm_out[MDATA][19] , \spm_out[MDATA][18] ,
         \spm_out[MDATA][17] , \spm_out[MDATA][16] , \spm_out[MDATA][15] ,
         \spm_out[MDATA][14] , \spm_out[MDATA][13] , \spm_out[MDATA][12] ,
         \spm_out[MDATA][11] , \spm_out[MDATA][10] , \spm_out[MDATA][9] ,
         \spm_out[MDATA][8] , \spm_out[MDATA][7] , \spm_out[MDATA][6] ,
         \spm_out[MDATA][5] , \spm_out[MDATA][4] , \spm_out[MDATA][3] ,
         \spm_out[MDATA][2] , \spm_out[MDATA][1] , \spm_out[MDATA][0] ;
  wire   \spm_out[MCMD][0] , \phase_prev[0] , \phase_next[1] , vld_pkt,
         \add_545/A[8] , \add_545/A[9] , \add_545/A[10] , \add_545/A[11] ,
         \add_545/A[12] , \add_545/A[13] , \add_545/A[14] , \add_545/A[15] ,
         \sub_544/A[1] , \sub_544/A[2] , \sub_544/A[3] , \sub_544/A[4] ,
         \sub_544/A[5] , \sub_544/A[6] , \sub_544/A[7] , \sub_544/A[8] ,
         \sub_544/A[9] , \sub_544/A[10] , \sub_544/A[11] , \sub_544/A[12] , n1,
         n2, n3, n4, n5, n6, n15, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n34, n35, n37, n39, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n62, n64, n72, n73, n74, n75, n77, n78, n79, n80, n84, n87,
         n88, n89, n90, n91, n93, n94, n95, n101, n102, n103, n104, n105, n106,
         n108, n109, n111, n112, n113, n114, n116, n117, n118, n120, n122,
         n124, n125, n127, n128, n129, n130, n132, n133, n134, n136, n137,
         n138, n139, n140, n142, n144, n149, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n310, n311,
         n312, n313, n314, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879;
  wire   [2:0] slt_index;
  wire   [2:0] dma_ren;
  wire   [2:0] dma_wen;
  wire   [1:0] dma_waddr;
  wire   [63:0] dma_wdata;
  wire   [1:0] dma_raddr;
  wire   [63:0] dma_rdata;
  wire   [4:0] slt_entry;
  wire   [1:0] state_cnt;
  wire   [4:0] config_reg;
  wire   [70:64] flit_buf;
  wire   [34:0] phitIn;
  wire   [31:0] mux_out;
  wire   [31:0] dOut_l;
  wire   [34:32] phit_togo;
  wire   [34:0] phitOut0;
  wire   [34:0] phitOut1;
  wire   [34:0] phitOut2;
  wire   [13:0] dma_cnt_new;
  wire   [15:0] dma_rp_new;
  wire   [15:0] dma_wp_new;
  wire   [6:0] address;
  wire   [31:0] dIn_h;
  assign \spm_out[MADDR][15]  = 1'b0;
  assign \spm_out[MADDR][16]  = 1'b0;
  assign \spm_out[MADDR][17]  = 1'b0;
  assign \spm_out[MADDR][18]  = 1'b0;
  assign \spm_out[MADDR][19]  = 1'b0;
  assign \spm_out[MADDR][20]  = 1'b0;
  assign \spm_out[MADDR][21]  = 1'b0;
  assign \spm_out[MADDR][22]  = 1'b0;
  assign \spm_out[MADDR][23]  = 1'b0;
  assign \spm_out[MADDR][24]  = 1'b0;
  assign \spm_out[MADDR][25]  = 1'b0;
  assign \spm_out[MADDR][26]  = 1'b0;
  assign \spm_out[MADDR][27]  = 1'b0;
  assign \spm_out[MADDR][28]  = 1'b0;
  assign \spm_out[MADDR][29]  = 1'b0;
  assign \spm_out[MADDR][30]  = 1'b0;
  assign \spm_out[MADDR][31]  = 1'b0;
  assign \spm_out[MCMD][1]  = \spm_out[MCMD][0] ;

  HS65_LS_DFPRQX9 \state_cnt_reg[0]  ( .D(n137), .CP(na_clk), .RN(n337), .Q(
        state_cnt[0]) );
  HS65_LS_DFPRQX9 \state_cnt_reg[1]  ( .D(n598), .CP(na_clk), .RN(n338), .Q(
        state_cnt[1]) );
  HS65_LS_DFPRQX9 \phase_next_reg[1]  ( .D(n677), .CP(na_clk), .RN(n340), .Q(
        \phase_next[1] ) );
  HS65_LS_DFPRQX9 \dOut_l_reg[31]  ( .D(n687), .CP(na_clk), .RN(n350), .Q(
        dOut_l[31]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[30]  ( .D(n688), .CP(na_clk), .RN(n338), .Q(
        dOut_l[30]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[29]  ( .D(n689), .CP(na_clk), .RN(n342), .Q(
        dOut_l[29]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[28]  ( .D(n690), .CP(na_clk), .RN(n349), .Q(
        dOut_l[28]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[27]  ( .D(n691), .CP(na_clk), .RN(n341), .Q(
        dOut_l[27]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[26]  ( .D(n692), .CP(na_clk), .RN(n339), .Q(
        dOut_l[26]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[25]  ( .D(n693), .CP(na_clk), .RN(n340), .Q(
        dOut_l[25]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[24]  ( .D(n694), .CP(na_clk), .RN(n345), .Q(
        dOut_l[24]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[23]  ( .D(n695), .CP(na_clk), .RN(n351), .Q(
        dOut_l[23]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[22]  ( .D(n696), .CP(na_clk), .RN(n339), .Q(
        dOut_l[22]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[21]  ( .D(n697), .CP(na_clk), .RN(n337), .Q(
        dOut_l[21]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[20]  ( .D(n698), .CP(na_clk), .RN(n341), .Q(
        dOut_l[20]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[19]  ( .D(n699), .CP(na_clk), .RN(n338), .Q(
        dOut_l[19]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[18]  ( .D(n700), .CP(na_clk), .RN(n343), .Q(
        dOut_l[18]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[17]  ( .D(n701), .CP(na_clk), .RN(n348), .Q(
        dOut_l[17]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[16]  ( .D(n702), .CP(na_clk), .RN(n338), .Q(
        dOut_l[16]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[15]  ( .D(n703), .CP(na_clk), .RN(n337), .Q(
        dOut_l[15]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[14]  ( .D(n704), .CP(na_clk), .RN(n341), .Q(
        dOut_l[14]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[13]  ( .D(n705), .CP(na_clk), .RN(n343), .Q(
        dOut_l[13]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[12]  ( .D(n706), .CP(na_clk), .RN(n347), .Q(
        dOut_l[12]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[11]  ( .D(n707), .CP(na_clk), .RN(n351), .Q(
        dOut_l[11]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[10]  ( .D(n708), .CP(na_clk), .RN(n342), .Q(
        dOut_l[10]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[9]  ( .D(n709), .CP(na_clk), .RN(n346), .Q(
        dOut_l[9]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[8]  ( .D(n710), .CP(na_clk), .RN(n344), .Q(
        dOut_l[8]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[7]  ( .D(n711), .CP(na_clk), .RN(n349), .Q(
        dOut_l[7]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[6]  ( .D(n712), .CP(na_clk), .RN(n350), .Q(
        dOut_l[6]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[5]  ( .D(n713), .CP(na_clk), .RN(n340), .Q(
        dOut_l[5]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[4]  ( .D(n714), .CP(na_clk), .RN(n345), .Q(
        dOut_l[4]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[3]  ( .D(n715), .CP(na_clk), .RN(n339), .Q(
        dOut_l[3]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[2]  ( .D(n716), .CP(na_clk), .RN(n346), .Q(
        dOut_l[2]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[1]  ( .D(n717), .CP(na_clk), .RN(n346), .Q(
        dOut_l[1]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[0]  ( .D(n718), .CP(na_clk), .RN(n346), .Q(
        dOut_l[0]) );
  HS65_LS_DFPRQX9 \phitIn_reg[34]  ( .D(pkt_in[34]), .CP(na_clk), .RN(n346), 
        .Q(phitIn[34]) );
  HS65_LS_DFPRQX9 \phitIn_reg[33]  ( .D(pkt_in[33]), .CP(na_clk), .RN(n346), 
        .Q(phitIn[33]) );
  HS65_LS_DFPRQX9 vld_pkt_reg ( .D(n680), .CP(na_clk), .RN(n346), .Q(vld_pkt)
         );
  HS65_LS_DFPRQX9 \phitIn_reg[32]  ( .D(pkt_in[32]), .CP(na_clk), .RN(n346), 
        .Q(phitIn[32]) );
  HS65_LS_DFPRQX9 \phitIn_reg[31]  ( .D(pkt_in[31]), .CP(na_clk), .RN(n346), 
        .Q(phitIn[31]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[31]  ( .D(n719), .CP(na_clk), .RN(n346), .Q(
        dIn_h[31]) );
  HS65_LS_DFPRQX9 \phitIn_reg[30]  ( .D(pkt_in[30]), .CP(na_clk), .RN(n346), 
        .Q(phitIn[30]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[30]  ( .D(n720), .CP(na_clk), .RN(n346), .Q(
        dIn_h[30]) );
  HS65_LS_DFPRQX9 \phitIn_reg[29]  ( .D(pkt_in[29]), .CP(na_clk), .RN(n346), 
        .Q(phitIn[29]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[29]  ( .D(n721), .CP(na_clk), .RN(n346), .Q(
        dIn_h[29]) );
  HS65_LS_DFPRQX9 \phitIn_reg[28]  ( .D(pkt_in[28]), .CP(na_clk), .RN(n346), 
        .Q(phitIn[28]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[28]  ( .D(n722), .CP(na_clk), .RN(n346), .Q(
        dIn_h[28]) );
  HS65_LS_DFPRQX9 \phitIn_reg[27]  ( .D(pkt_in[27]), .CP(na_clk), .RN(n347), 
        .Q(phitIn[27]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[27]  ( .D(n723), .CP(na_clk), .RN(n347), .Q(
        dIn_h[27]) );
  HS65_LS_DFPRQX9 \phitIn_reg[26]  ( .D(pkt_in[26]), .CP(na_clk), .RN(n347), 
        .Q(phitIn[26]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[26]  ( .D(n724), .CP(na_clk), .RN(n347), .Q(
        dIn_h[26]) );
  HS65_LS_DFPRQX9 \phitIn_reg[25]  ( .D(pkt_in[25]), .CP(na_clk), .RN(n347), 
        .Q(phitIn[25]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[25]  ( .D(n725), .CP(na_clk), .RN(n347), .Q(
        dIn_h[25]) );
  HS65_LS_DFPRQX9 \phitIn_reg[24]  ( .D(pkt_in[24]), .CP(na_clk), .RN(n347), 
        .Q(phitIn[24]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[24]  ( .D(n726), .CP(na_clk), .RN(n347), .Q(
        dIn_h[24]) );
  HS65_LS_DFPRQX9 \phitIn_reg[23]  ( .D(pkt_in[23]), .CP(na_clk), .RN(n347), 
        .Q(phitIn[23]) );
  HS65_LS_DFPRQX9 \address_reg[6]  ( .D(n727), .CP(na_clk), .RN(n347), .Q(
        address[6]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[23]  ( .D(n728), .CP(na_clk), .RN(n347), .Q(
        dIn_h[23]) );
  HS65_LS_DFPRQX9 \phitIn_reg[22]  ( .D(pkt_in[22]), .CP(na_clk), .RN(n347), 
        .Q(phitIn[22]) );
  HS65_LS_DFPRQX9 \address_reg[5]  ( .D(n729), .CP(na_clk), .RN(n347), .Q(
        address[5]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[22]  ( .D(n730), .CP(na_clk), .RN(n347), .Q(
        dIn_h[22]) );
  HS65_LS_DFPRQX9 \phitIn_reg[21]  ( .D(pkt_in[21]), .CP(na_clk), .RN(n347), 
        .Q(phitIn[21]) );
  HS65_LS_DFPRQX9 \address_reg[4]  ( .D(n731), .CP(na_clk), .RN(n340), .Q(
        address[4]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[21]  ( .D(n732), .CP(na_clk), .RN(n339), .Q(
        dIn_h[21]) );
  HS65_LS_DFPRQX9 \phitIn_reg[20]  ( .D(pkt_in[20]), .CP(na_clk), .RN(n342), 
        .Q(phitIn[20]) );
  HS65_LS_DFPRQX9 \address_reg[3]  ( .D(n733), .CP(na_clk), .RN(n337), .Q(
        address[3]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[20]  ( .D(n734), .CP(na_clk), .RN(n343), .Q(
        dIn_h[20]) );
  HS65_LS_DFPRQX9 \phitIn_reg[19]  ( .D(pkt_in[19]), .CP(na_clk), .RN(n345), 
        .Q(phitIn[19]) );
  HS65_LS_DFPRQX9 \address_reg[2]  ( .D(n735), .CP(na_clk), .RN(n350), .Q(
        address[2]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[19]  ( .D(n736), .CP(na_clk), .RN(n349), .Q(
        dIn_h[19]) );
  HS65_LS_DFPRQX9 \phitIn_reg[18]  ( .D(pkt_in[18]), .CP(na_clk), .RN(n342), 
        .Q(phitIn[18]) );
  HS65_LS_DFPRQX9 \address_reg[1]  ( .D(n737), .CP(na_clk), .RN(n346), .Q(
        address[1]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[18]  ( .D(n738), .CP(na_clk), .RN(n344), .Q(
        dIn_h[18]) );
  HS65_LS_DFPRQX9 \phitIn_reg[17]  ( .D(pkt_in[17]), .CP(na_clk), .RN(n347), 
        .Q(phitIn[17]) );
  HS65_LS_DFPRQX9 \address_reg[0]  ( .D(n739), .CP(na_clk), .RN(n344), .Q(
        address[0]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[17]  ( .D(n740), .CP(na_clk), .RN(n348), .Q(
        dIn_h[17]) );
  HS65_LS_DFPRQX9 \phitIn_reg[16]  ( .D(pkt_in[16]), .CP(na_clk), .RN(n348), 
        .Q(phitIn[16]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[16]  ( .D(n741), .CP(na_clk), .RN(n348), .Q(
        dIn_h[16]) );
  HS65_LS_DFPRQX9 \phitIn_reg[15]  ( .D(pkt_in[15]), .CP(na_clk), .RN(n348), 
        .Q(phitIn[15]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[15]  ( .D(n742), .CP(na_clk), .RN(n348), .Q(
        dIn_h[15]) );
  HS65_LS_DFPRQX9 \phitIn_reg[14]  ( .D(pkt_in[14]), .CP(na_clk), .RN(n348), 
        .Q(phitIn[14]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[14]  ( .D(n743), .CP(na_clk), .RN(n348), .Q(
        dIn_h[14]) );
  HS65_LS_DFPRQX9 \phitIn_reg[13]  ( .D(pkt_in[13]), .CP(na_clk), .RN(n348), 
        .Q(phitIn[13]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[13]  ( .D(n744), .CP(na_clk), .RN(n348), .Q(
        dIn_h[13]) );
  HS65_LS_DFPRQX9 \phitIn_reg[12]  ( .D(pkt_in[12]), .CP(na_clk), .RN(n348), 
        .Q(phitIn[12]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[12]  ( .D(n745), .CP(na_clk), .RN(n348), .Q(
        dIn_h[12]) );
  HS65_LS_DFPRQX9 \phitIn_reg[11]  ( .D(pkt_in[11]), .CP(na_clk), .RN(n348), 
        .Q(phitIn[11]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[11]  ( .D(n746), .CP(na_clk), .RN(n348), .Q(
        dIn_h[11]) );
  HS65_LS_DFPRQX9 \phitIn_reg[10]  ( .D(pkt_in[10]), .CP(na_clk), .RN(n348), 
        .Q(phitIn[10]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[10]  ( .D(n747), .CP(na_clk), .RN(n348), .Q(
        dIn_h[10]) );
  HS65_LS_DFPRQX9 \phitIn_reg[9]  ( .D(pkt_in[9]), .CP(na_clk), .RN(n348), .Q(
        phitIn[9]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[9]  ( .D(n748), .CP(na_clk), .RN(n349), .Q(
        dIn_h[9]) );
  HS65_LS_DFPRQX9 \phitIn_reg[8]  ( .D(pkt_in[8]), .CP(na_clk), .RN(n349), .Q(
        phitIn[8]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[8]  ( .D(n749), .CP(na_clk), .RN(n349), .Q(
        dIn_h[8]) );
  HS65_LS_DFPRQX9 \phitIn_reg[7]  ( .D(pkt_in[7]), .CP(na_clk), .RN(n349), .Q(
        phitIn[7]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[7]  ( .D(n750), .CP(na_clk), .RN(n349), .Q(
        dIn_h[7]) );
  HS65_LS_DFPRQX9 \phitIn_reg[6]  ( .D(pkt_in[6]), .CP(na_clk), .RN(n349), .Q(
        phitIn[6]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[6]  ( .D(n751), .CP(na_clk), .RN(n349), .Q(
        dIn_h[6]) );
  HS65_LS_DFPRQX9 \phitIn_reg[5]  ( .D(pkt_in[5]), .CP(na_clk), .RN(n349), .Q(
        phitIn[5]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[5]  ( .D(n752), .CP(na_clk), .RN(n349), .Q(
        dIn_h[5]) );
  HS65_LS_DFPRQX9 \phitIn_reg[4]  ( .D(pkt_in[4]), .CP(na_clk), .RN(n349), .Q(
        phitIn[4]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[4]  ( .D(n753), .CP(na_clk), .RN(n349), .Q(
        dIn_h[4]) );
  HS65_LS_DFPRQX9 \phitIn_reg[3]  ( .D(pkt_in[3]), .CP(na_clk), .RN(n349), .Q(
        phitIn[3]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[3]  ( .D(n754), .CP(na_clk), .RN(n349), .Q(
        dIn_h[3]) );
  HS65_LS_DFPRQX9 \phitIn_reg[2]  ( .D(pkt_in[2]), .CP(na_clk), .RN(n349), .Q(
        phitIn[2]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[2]  ( .D(n755), .CP(na_clk), .RN(n349), .Q(
        dIn_h[2]) );
  HS65_LS_DFPRQX9 \phitIn_reg[1]  ( .D(pkt_in[1]), .CP(na_clk), .RN(n350), .Q(
        phitIn[1]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[1]  ( .D(n756), .CP(na_clk), .RN(n350), .Q(
        dIn_h[1]) );
  HS65_LS_DFPRQX9 \phitIn_reg[0]  ( .D(pkt_in[0]), .CP(na_clk), .RN(n350), .Q(
        phitIn[0]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[0]  ( .D(n757), .CP(na_clk), .RN(n350), .Q(
        dIn_h[0]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[34]  ( .D(phit_togo[34]), .CP(na_clk), .RN(
        n350), .Q(phitOut0[34]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[33]  ( .D(n329), .CP(na_clk), .RN(n350), .Q(
        phitOut0[33]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[32]  ( .D(phit_togo[32]), .CP(na_clk), .RN(
        n350), .Q(phitOut0[32]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[31]  ( .D(mux_out[31]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[31]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[30]  ( .D(mux_out[30]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[30]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[29]  ( .D(mux_out[29]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[29]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[28]  ( .D(mux_out[28]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[28]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[27]  ( .D(mux_out[27]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[27]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[26]  ( .D(mux_out[26]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[26]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[25]  ( .D(mux_out[25]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[25]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[24]  ( .D(mux_out[24]), .CP(na_clk), .RN(n350), 
        .Q(phitOut0[24]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[23]  ( .D(mux_out[23]), .CP(na_clk), .RN(n351), 
        .Q(phitOut0[23]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[22]  ( .D(mux_out[22]), .CP(na_clk), .RN(n351), 
        .Q(phitOut0[22]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[21]  ( .D(mux_out[21]), .CP(na_clk), .RN(n351), 
        .Q(phitOut0[21]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[20]  ( .D(mux_out[20]), .CP(na_clk), .RN(n351), 
        .Q(phitOut0[20]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[19]  ( .D(mux_out[19]), .CP(na_clk), .RN(n351), 
        .Q(phitOut0[19]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[18]  ( .D(mux_out[18]), .CP(na_clk), .RN(n351), 
        .Q(phitOut0[18]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[17]  ( .D(mux_out[17]), .CP(na_clk), .RN(n351), 
        .Q(phitOut0[17]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[16]  ( .D(mux_out[16]), .CP(na_clk), .RN(n351), 
        .Q(phitOut0[16]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[15]  ( .D(mux_out[15]), .CP(na_clk), .RN(n351), 
        .Q(phitOut0[15]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[14]  ( .D(mux_out[14]), .CP(na_clk), .RN(n351), 
        .Q(phitOut0[14]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[13]  ( .D(mux_out[13]), .CP(na_clk), .RN(n351), 
        .Q(phitOut0[13]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[12]  ( .D(mux_out[12]), .CP(na_clk), .RN(n351), 
        .Q(phitOut0[12]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[11]  ( .D(mux_out[11]), .CP(na_clk), .RN(n351), 
        .Q(phitOut0[11]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[10]  ( .D(mux_out[10]), .CP(na_clk), .RN(n351), 
        .Q(phitOut0[10]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[9]  ( .D(mux_out[9]), .CP(na_clk), .RN(n351), 
        .Q(phitOut0[9]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[8]  ( .D(mux_out[8]), .CP(na_clk), .RN(n351), 
        .Q(phitOut0[8]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[7]  ( .D(mux_out[7]), .CP(na_clk), .RN(n344), 
        .Q(phitOut0[7]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[6]  ( .D(mux_out[6]), .CP(na_clk), .RN(n341), 
        .Q(phitOut0[6]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[5]  ( .D(mux_out[5]), .CP(na_clk), .RN(n338), 
        .Q(phitOut0[5]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[4]  ( .D(mux_out[4]), .CP(na_clk), .RN(n339), 
        .Q(phitOut0[4]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[3]  ( .D(mux_out[3]), .CP(na_clk), .RN(n340), 
        .Q(phitOut0[3]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[2]  ( .D(mux_out[2]), .CP(na_clk), .RN(n342), 
        .Q(phitOut0[2]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[1]  ( .D(mux_out[1]), .CP(na_clk), .RN(n343), 
        .Q(phitOut0[1]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[0]  ( .D(mux_out[0]), .CP(na_clk), .RN(n337), 
        .Q(phitOut0[0]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[34]  ( .D(phitOut0[34]), .CP(na_clk), .RN(n341), .Q(phitOut1[34]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[33]  ( .D(phitOut0[33]), .CP(na_clk), .RN(n337), .Q(phitOut1[33]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[32]  ( .D(phitOut0[32]), .CP(na_clk), .RN(n337), .Q(phitOut1[32]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[31]  ( .D(phitOut0[31]), .CP(na_clk), .RN(n337), .Q(phitOut1[31]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[30]  ( .D(phitOut0[30]), .CP(na_clk), .RN(n337), .Q(phitOut1[30]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[29]  ( .D(phitOut0[29]), .CP(na_clk), .RN(n337), .Q(phitOut1[29]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[28]  ( .D(phitOut0[28]), .CP(na_clk), .RN(n337), .Q(phitOut1[28]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[27]  ( .D(phitOut0[27]), .CP(na_clk), .RN(n337), .Q(phitOut1[27]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[26]  ( .D(phitOut0[26]), .CP(na_clk), .RN(n337), .Q(phitOut1[26]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[25]  ( .D(phitOut0[25]), .CP(na_clk), .RN(n337), .Q(phitOut1[25]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[24]  ( .D(phitOut0[24]), .CP(na_clk), .RN(n337), .Q(phitOut1[24]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[23]  ( .D(phitOut0[23]), .CP(na_clk), .RN(n337), .Q(phitOut1[23]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[22]  ( .D(phitOut0[22]), .CP(na_clk), .RN(n337), .Q(phitOut1[22]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[21]  ( .D(phitOut0[21]), .CP(na_clk), .RN(n337), .Q(phitOut1[21]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[20]  ( .D(phitOut0[20]), .CP(na_clk), .RN(n344), .Q(phitOut1[20]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[19]  ( .D(phitOut0[19]), .CP(na_clk), .RN(n348), .Q(phitOut1[19]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[18]  ( .D(phitOut0[18]), .CP(na_clk), .RN(n349), .Q(phitOut1[18]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[17]  ( .D(phitOut0[17]), .CP(na_clk), .RN(n346), .Q(phitOut1[17]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[16]  ( .D(phitOut0[16]), .CP(na_clk), .RN(n347), .Q(phitOut1[16]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[15]  ( .D(phitOut0[15]), .CP(na_clk), .RN(n350), .Q(phitOut1[15]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[14]  ( .D(phitOut0[14]), .CP(na_clk), .RN(n345), .Q(phitOut1[14]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[13]  ( .D(phitOut0[13]), .CP(na_clk), .RN(n341), .Q(phitOut1[13]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[12]  ( .D(phitOut0[12]), .CP(na_clk), .RN(n351), .Q(phitOut1[12]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[11]  ( .D(phitOut0[11]), .CP(na_clk), .RN(n343), .Q(phitOut1[11]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[10]  ( .D(phitOut0[10]), .CP(na_clk), .RN(n351), .Q(phitOut1[10]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[9]  ( .D(phitOut0[9]), .CP(na_clk), .RN(n346), 
        .Q(phitOut1[9]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[8]  ( .D(phitOut0[8]), .CP(na_clk), .RN(n347), 
        .Q(phitOut1[8]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[7]  ( .D(phitOut0[7]), .CP(na_clk), .RN(n348), 
        .Q(phitOut1[7]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[6]  ( .D(phitOut0[6]), .CP(na_clk), .RN(n338), 
        .Q(phitOut1[6]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[5]  ( .D(phitOut0[5]), .CP(na_clk), .RN(n338), 
        .Q(phitOut1[5]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[4]  ( .D(phitOut0[4]), .CP(na_clk), .RN(n338), 
        .Q(phitOut1[4]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[3]  ( .D(phitOut0[3]), .CP(na_clk), .RN(n338), 
        .Q(phitOut1[3]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[2]  ( .D(phitOut0[2]), .CP(na_clk), .RN(n338), 
        .Q(phitOut1[2]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[1]  ( .D(phitOut0[1]), .CP(na_clk), .RN(n338), 
        .Q(phitOut1[1]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[0]  ( .D(phitOut0[0]), .CP(na_clk), .RN(n338), 
        .Q(phitOut1[0]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[34]  ( .D(phitOut1[34]), .CP(na_clk), .RN(n338), .Q(phitOut2[34]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[33]  ( .D(phitOut1[33]), .CP(na_clk), .RN(n338), .Q(phitOut2[33]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[32]  ( .D(phitOut1[32]), .CP(na_clk), .RN(n338), .Q(phitOut2[32]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[31]  ( .D(phitOut1[31]), .CP(na_clk), .RN(n338), .Q(phitOut2[31]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[30]  ( .D(phitOut1[30]), .CP(na_clk), .RN(n338), .Q(phitOut2[30]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[29]  ( .D(phitOut1[29]), .CP(na_clk), .RN(n338), .Q(phitOut2[29]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[28]  ( .D(phitOut1[28]), .CP(na_clk), .RN(n338), .Q(phitOut2[28]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[27]  ( .D(phitOut1[27]), .CP(na_clk), .RN(n338), .Q(phitOut2[27]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[26]  ( .D(phitOut1[26]), .CP(na_clk), .RN(n339), .Q(phitOut2[26]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[25]  ( .D(phitOut1[25]), .CP(na_clk), .RN(n339), .Q(phitOut2[25]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[24]  ( .D(phitOut1[24]), .CP(na_clk), .RN(n339), .Q(phitOut2[24]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[23]  ( .D(phitOut1[23]), .CP(na_clk), .RN(n339), .Q(phitOut2[23]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[22]  ( .D(phitOut1[22]), .CP(na_clk), .RN(n339), .Q(phitOut2[22]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[21]  ( .D(phitOut1[21]), .CP(na_clk), .RN(n339), .Q(phitOut2[21]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[20]  ( .D(phitOut1[20]), .CP(na_clk), .RN(n339), .Q(phitOut2[20]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[19]  ( .D(phitOut1[19]), .CP(na_clk), .RN(n339), .Q(phitOut2[19]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[18]  ( .D(phitOut1[18]), .CP(na_clk), .RN(n339), .Q(phitOut2[18]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[17]  ( .D(phitOut1[17]), .CP(na_clk), .RN(n339), .Q(phitOut2[17]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[16]  ( .D(phitOut1[16]), .CP(na_clk), .RN(n339), .Q(phitOut2[16]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[15]  ( .D(phitOut1[15]), .CP(na_clk), .RN(n339), .Q(phitOut2[15]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[14]  ( .D(phitOut1[14]), .CP(na_clk), .RN(n339), .Q(phitOut2[14]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[13]  ( .D(phitOut1[13]), .CP(na_clk), .RN(n339), .Q(phitOut2[13]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[12]  ( .D(phitOut1[12]), .CP(na_clk), .RN(n339), .Q(phitOut2[12]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[11]  ( .D(phitOut1[11]), .CP(na_clk), .RN(n340), .Q(phitOut2[11]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[10]  ( .D(phitOut1[10]), .CP(na_clk), .RN(n340), .Q(phitOut2[10]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[9]  ( .D(phitOut1[9]), .CP(na_clk), .RN(n340), 
        .Q(phitOut2[9]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[8]  ( .D(phitOut1[8]), .CP(na_clk), .RN(n340), 
        .Q(phitOut2[8]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[7]  ( .D(phitOut1[7]), .CP(na_clk), .RN(n340), 
        .Q(phitOut2[7]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[6]  ( .D(phitOut1[6]), .CP(na_clk), .RN(n340), 
        .Q(phitOut2[6]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[5]  ( .D(phitOut1[5]), .CP(na_clk), .RN(n340), 
        .Q(phitOut2[5]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[4]  ( .D(phitOut1[4]), .CP(na_clk), .RN(n340), 
        .Q(phitOut2[4]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[3]  ( .D(phitOut1[3]), .CP(na_clk), .RN(n340), 
        .Q(phitOut2[3]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[2]  ( .D(phitOut1[2]), .CP(na_clk), .RN(n340), 
        .Q(phitOut2[2]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[1]  ( .D(phitOut1[1]), .CP(na_clk), .RN(n340), 
        .Q(phitOut2[1]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[0]  ( .D(phitOut1[0]), .CP(na_clk), .RN(n340), 
        .Q(phitOut2[0]) );
  HS65_LS_DFPRQX9 \config_reg_reg[4]  ( .D(\proc_in[MCMD][1] ), .CP(na_clk), 
        .RN(n340), .Q(config_reg[4]) );
  HS65_LS_DFPRQX9 \config_reg_reg[3]  ( .D(n676), .CP(na_clk), .RN(n340), .Q(
        config_reg[3]) );
  HS65_LS_DFPRQX9 \config_reg_reg[2]  ( .D(n653), .CP(na_clk), .RN(n340), .Q(
        config_reg[2]) );
  HS65_LS_DFPRQX9 \config_reg_reg[1]  ( .D(n654), .CP(na_clk), .RN(n341), .Q(
        config_reg[1]) );
  HS65_LS_DFPRQX9 \config_reg_reg[0]  ( .D(n652), .CP(na_clk), .RN(n341), .Q(
        config_reg[0]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[70]  ( .D(n758), .CP(na_clk), .RN(n341), .Q(
        flit_buf[70]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[69]  ( .D(n759), .CP(na_clk), .RN(n341), .Q(
        flit_buf[69]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[68]  ( .D(n760), .CP(na_clk), .RN(n341), .Q(
        flit_buf[68]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[67]  ( .D(n761), .CP(na_clk), .RN(n341), .Q(
        flit_buf[67]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[66]  ( .D(n762), .CP(na_clk), .RN(n341), .Q(
        flit_buf[66]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[65]  ( .D(n763), .CP(na_clk), .RN(n341), .Q(
        flit_buf[65]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[64]  ( .D(n764), .CP(na_clk), .RN(n341), .Q(
        flit_buf[64]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[63]  ( .D(n765), .CP(na_clk), .RN(n341), .Q(
        \spm_out[MDATA][63] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[62]  ( .D(n766), .CP(na_clk), .RN(n341), .Q(
        \spm_out[MDATA][62] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[61]  ( .D(n767), .CP(na_clk), .RN(n341), .Q(
        \spm_out[MDATA][61] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[60]  ( .D(n768), .CP(na_clk), .RN(n341), .Q(
        \spm_out[MDATA][60] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[59]  ( .D(n769), .CP(na_clk), .RN(n341), .Q(
        \spm_out[MDATA][59] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[58]  ( .D(n770), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][58] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[57]  ( .D(n771), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][57] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[56]  ( .D(n772), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][56] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[55]  ( .D(n773), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][55] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[54]  ( .D(n774), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][54] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[53]  ( .D(n775), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][53] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[52]  ( .D(n776), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][52] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[51]  ( .D(n777), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][51] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[50]  ( .D(n778), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][50] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[49]  ( .D(n779), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][49] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[48]  ( .D(n780), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][48] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[47]  ( .D(n781), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][47] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[46]  ( .D(n782), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][46] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[45]  ( .D(n783), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][45] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[44]  ( .D(n784), .CP(na_clk), .RN(n342), .Q(
        \spm_out[MDATA][44] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[43]  ( .D(n785), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][43] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[42]  ( .D(n786), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][42] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[41]  ( .D(n787), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][41] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[40]  ( .D(n788), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][40] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[39]  ( .D(n789), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][39] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[38]  ( .D(n790), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][38] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[37]  ( .D(n791), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][37] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[36]  ( .D(n792), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][36] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[35]  ( .D(n793), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][35] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[34]  ( .D(n794), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][34] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[33]  ( .D(n795), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][33] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[32]  ( .D(n796), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][32] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[31]  ( .D(n797), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][31] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[30]  ( .D(n798), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][30] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[29]  ( .D(n799), .CP(na_clk), .RN(n343), .Q(
        \spm_out[MDATA][29] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[28]  ( .D(n800), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][28] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[27]  ( .D(n801), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][27] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[26]  ( .D(n802), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][26] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[25]  ( .D(n803), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][25] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[24]  ( .D(n804), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][24] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[23]  ( .D(n805), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][23] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[22]  ( .D(n806), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][22] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[21]  ( .D(n807), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][21] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[20]  ( .D(n808), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][20] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[19]  ( .D(n809), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][19] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[18]  ( .D(n810), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][18] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[17]  ( .D(n811), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][17] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[16]  ( .D(n812), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][16] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[15]  ( .D(n813), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][15] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[14]  ( .D(n814), .CP(na_clk), .RN(n344), .Q(
        \spm_out[MDATA][14] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[13]  ( .D(n815), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][13] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[12]  ( .D(n816), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][12] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[11]  ( .D(n817), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][11] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[10]  ( .D(n818), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][10] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[9]  ( .D(n819), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][9] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[8]  ( .D(n820), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][8] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[7]  ( .D(n821), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][7] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[6]  ( .D(n822), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][6] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[5]  ( .D(n823), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][5] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[4]  ( .D(n824), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][4] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[3]  ( .D(n825), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][3] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[2]  ( .D(n826), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][2] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[1]  ( .D(n827), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][1] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[0]  ( .D(n828), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][0] ) );
  HS65_LS_DFPRQX9 \phase_prev_reg[0]  ( .D(n683), .CP(na_clk), .RN(n345), .Q(
        \phase_prev[0] ) );
  counter_WIDTH3_3 slt_cnt ( .clk(na_clk), .reset(n352), .enable(n648), .cnt(
        slt_index) );
  dma_sdp_DATA64_ADDR2_3 dma_table ( .clk(na_clk), .reset(n353), .ren(dma_ren), 
        .wen(dma_wen), .waddr(dma_waddr), .wdata(dma_wdata), .raddr(dma_raddr), 
        .rdata(dma_rdata) );
  bram_DATA5_ADDR3_3 slt_table ( .clk(na_clk), .reset(n352), .rd_addr(
        slt_index), .wr_addr({\proc_in[MADDR][2] , \proc_in[MADDR][1] , 
        \proc_in[MADDR][0] }), .wr_data({\proc_in[MDATA][4] , 
        \proc_in[MDATA][3] , \proc_in[MDATA][2] , \proc_in[MDATA][1] , 
        \proc_in[MDATA][0] }), .wr_ena(n651), .rd_data(slt_entry) );
  HS65_LS_DFPRQNX9 vld_buf_reg ( .D(n681), .CP(na_clk), .RN(n345), .QN(n684)
         );
  HS65_LS_DFPRQNX9 dma_ctrl_reg_reg ( .D(n679), .CP(na_clk), .RN(n349), .QN(
        n685) );
  HS65_LS_DFPRQNX9 \phase_next_reg[0]  ( .D(n678), .CP(na_clk), .RN(n350), 
        .QN(n686) );
  HS65_LS_DFPRQX9 \phase_prev_reg[1]  ( .D(n682), .CP(na_clk), .RN(n337), .Q(
        n21) );
  HS65_LS_IVX35 U3 ( .A(n465), .Z(n567) );
  HS65_LS_IVX27 U4 ( .A(n112), .Z(n114) );
  HS65_LS_IVX18 U5 ( .A(n576), .Z(n113) );
  HS65_LS_IVX44 U6 ( .A(n5), .Z(n526) );
  HS65_LS_IVX31 U7 ( .A(n112), .Z(n116) );
  HS65_LS_AND2X27 U8 ( .A(n445), .B(n449), .Z(n120) );
  HS65_LS_OR2X27 U9 ( .A(n486), .B(n526), .Z(n28) );
  HS65_LS_IVX31 U10 ( .A(n576), .Z(n112) );
  HS65_LS_NAND2X7 U11 ( .A(phitOut2[5]), .B(n74), .Z(n482) );
  HS65_LS_IVX18 U12 ( .A(n113), .Z(n117) );
  HS65_LS_IVX22 U13 ( .A(n465), .Z(n472) );
  HS65_LS_NAND2X21 U14 ( .A(n105), .B(n573), .Z(n465) );
  HS65_LS_NAND2X5 U15 ( .A(phitOut2[11]), .B(n472), .Z(n500) );
  HS65_LS_IVX4 U16 ( .A(n573), .Z(n6) );
  HS65_LS_NAND2X14 U17 ( .A(n20), .B(n462), .Z(n450) );
  HS65_LS_OAI222X2 U18 ( .A(n658), .B(n851), .C(n646), .D(n37), .E(n657), .F(
        n853), .Z(dma_waddr[1]) );
  HS65_LS_OAI222X2 U19 ( .A(n659), .B(n851), .C(n647), .D(n37), .E(n658), .F(
        n853), .Z(dma_waddr[0]) );
  HS65_LS_IVX9 U20 ( .A(n460), .Z(n19) );
  HS65_LS_NAND3X13 U21 ( .A(n27), .B(n28), .C(n485), .Z(pkt_out[6]) );
  HS65_LS_AND2X4 U22 ( .A(\proc_in[MCMD][0] ), .B(n593), .Z(n1) );
  HS65_LS_AND2X4 U23 ( .A(n612), .B(n51), .Z(n2) );
  HS65_LS_AND2X4 U24 ( .A(\add_545/A[14] ), .B(n64), .Z(n3) );
  HS65_LS_AND2X4 U25 ( .A(n133), .B(n412), .Z(n4) );
  HS65_LS_NAND2X5 U26 ( .A(phitOut2[4]), .B(n74), .Z(n479) );
  HS65_LS_NAND2X5 U27 ( .A(phitOut2[12]), .B(n74), .Z(n503) );
  HS65_LS_NAND2X5 U28 ( .A(phitOut2[9]), .B(n74), .Z(n494) );
  HS65_LS_NAND2X5 U29 ( .A(phitOut2[8]), .B(n74), .Z(n491) );
  HS65_LS_NAND2X5 U30 ( .A(phitOut2[7]), .B(n74), .Z(n488) );
  HS65_LS_NAND2X4 U31 ( .A(phitOut2[6]), .B(n567), .Z(n485) );
  HS65_LS_NAND2X5 U32 ( .A(phitOut2[31]), .B(n567), .Z(n561) );
  HS65_LS_NAND2X5 U33 ( .A(phitOut2[30]), .B(n567), .Z(n558) );
  HS65_LS_NAND2X5 U34 ( .A(phitOut2[27]), .B(n567), .Z(n549) );
  HS65_LS_NAND2X5 U35 ( .A(phitOut2[23]), .B(n567), .Z(n537) );
  HS65_LS_NAND2X5 U36 ( .A(phitOut2[21]), .B(n567), .Z(n531) );
  HS65_LS_NAND2X5 U37 ( .A(phitOut2[32]), .B(n567), .Z(n564) );
  HS65_LS_NAND2X5 U38 ( .A(phitOut2[24]), .B(n567), .Z(n540) );
  HS65_LS_NAND2X5 U39 ( .A(phitOut2[22]), .B(n567), .Z(n534) );
  HS65_LS_NAND2X5 U40 ( .A(phitOut2[28]), .B(n567), .Z(n552) );
  HS65_LS_NAND2X5 U41 ( .A(phitOut2[33]), .B(n567), .Z(n568) );
  HS65_LS_NAND2X5 U42 ( .A(phitOut2[25]), .B(n567), .Z(n543) );
  HS65_LS_NAND2X5 U43 ( .A(phitOut2[20]), .B(n567), .Z(n528) );
  HS65_LS_NAND2X5 U44 ( .A(phitOut2[19]), .B(n567), .Z(n524) );
  HS65_LS_NAND2X5 U45 ( .A(phitOut2[17]), .B(n567), .Z(n518) );
  HS65_LS_NAND2X5 U46 ( .A(phitOut2[29]), .B(n567), .Z(n555) );
  HS65_LS_BFX27 U47 ( .A(n570), .Z(n22) );
  HS65_LS_NAND2X5 U48 ( .A(phitOut2[26]), .B(n567), .Z(n546) );
  HS65_LS_NAND2X5 U49 ( .A(phitOut2[16]), .B(n567), .Z(n515) );
  HS65_LS_IVX2 U50 ( .A(n32), .Z(n17) );
  HS65_LS_BFX18 U51 ( .A(n570), .Z(n24) );
  HS65_LS_NAND2X5 U52 ( .A(phitOut2[18]), .B(n567), .Z(n521) );
  HS65_LS_BFX27 U53 ( .A(n570), .Z(n23) );
  HS65_LS_IVX13 U54 ( .A(n113), .Z(n29) );
  HS65_LS_NOR2X13 U55 ( .A(n6), .B(n15), .Z(n74) );
  HS65_LS_IVX18 U56 ( .A(n450), .Z(n31) );
  HS65_LS_IVX9 U57 ( .A(n450), .Z(n457) );
  HS65_LS_NAND2X5 U58 ( .A(phitOut2[2]), .B(n472), .Z(n473) );
  HS65_LS_NAND2X5 U59 ( .A(phitOut2[1]), .B(n472), .Z(n469) );
  HS65_LS_NAND2X4 U60 ( .A(phitOut2[10]), .B(n472), .Z(n497) );
  HS65_LS_NAND2X4 U61 ( .A(phitOut2[3]), .B(n472), .Z(n476) );
  HS65_LS_NAND2X5 U62 ( .A(phitOut2[0]), .B(n472), .Z(n466) );
  HS65_LS_NAND2X5 U63 ( .A(phitOut2[13]), .B(n472), .Z(n506) );
  HS65_LS_NAND2X5 U64 ( .A(phitOut2[14]), .B(n472), .Z(n509) );
  HS65_LS_NAND2X5 U65 ( .A(phitOut2[15]), .B(n472), .Z(n512) );
  HS65_LS_NAND2X7 U66 ( .A(n572), .B(n105), .Z(n570) );
  HS65_LS_OAI21X24 U67 ( .A(n463), .B(n464), .C(n572), .Z(n576) );
  HS65_LS_IVX7 U68 ( .A(state_cnt[1]), .Z(n449) );
  HS65_LS_IVX9 U69 ( .A(n459), .Z(n460) );
  HS65_LS_IVX31 U70 ( .A(n573), .Z(n572) );
  HS65_LS_OAI21X6 U71 ( .A(n117), .B(n575), .C(n574), .Z(pkt_out[34]) );
  HS65_LS_NAND3X13 U72 ( .A(n120), .B(n452), .C(n453), .Z(n454) );
  HS65_LS_NAND2X29 U73 ( .A(n109), .B(n104), .Z(n573) );
  HS65_LS_AOI312X8 U74 ( .A(n122), .B(n120), .C(n462), .D(n461), .E(n26), .F(
        n460), .Z(n109) );
  HS65_LS_NAND2X4 U75 ( .A(state_cnt[0]), .B(state_cnt[1]), .Z(n459) );
  HS65_LS_IVX4 U76 ( .A(n105), .Z(n15) );
  HS65_LS_CB4I1X27 U77 ( .A(n31), .B(n456), .C(n455), .D(n454), .Z(n104) );
  HS65_LS_AND2X18 U78 ( .A(n105), .B(n572), .Z(n5) );
  HS65_LS_NAND2X14 U79 ( .A(n451), .B(n21), .Z(n458) );
  HS65_LS_NAND2X29 U80 ( .A(n458), .B(n35), .Z(n462) );
  HS65_LS_IVX4 U81 ( .A(n17), .Z(n18) );
  HS65_LS_IVX2 U82 ( .A(n445), .Z(n26) );
  HS65_LS_CBI4I1X16 U83 ( .A(n456), .B(n457), .C(n686), .D(n19), .Z(n463) );
  HS65_LS_IVX2 U84 ( .A(n458), .Z(n461) );
  HS65_LS_NAND2X21 U85 ( .A(n34), .B(n32), .Z(n35) );
  HS65_LS_IVX2 U86 ( .A(n32), .Z(n25) );
  HS65_LS_IVX9 U87 ( .A(state_cnt[1]), .Z(n20) );
  HS65_LS_IVX18 U88 ( .A(n21), .Z(n34) );
  HS65_LS_NAND2X5 U89 ( .A(state_cnt[0]), .B(n458), .Z(n456) );
  HS65_LS_IVX18 U90 ( .A(n451), .Z(n32) );
  HS65_LS_NAND2X5 U91 ( .A(n25), .B(n462), .Z(n447) );
  HS65_LS_OR2X18 U92 ( .A(n118), .B(n487), .Z(n27) );
  HS65_LS_OAI212X5 U93 ( .A(n116), .B(n468), .C(n526), .D(n467), .E(n466), .Z(
        pkt_out[0]) );
  HS65_LS_IVX7 U94 ( .A(n34), .Z(n122) );
  HS65_LS_IVX18 U95 ( .A(state_cnt[0]), .Z(n445) );
  HS65_LS_IVX9 U96 ( .A(n462), .Z(n453) );
  HS65_LS_AOI33X2 U97 ( .A(n573), .B(phitOut2[34]), .C(n105), .D(n105), .E(
        n572), .F(phitOut0[34]), .Z(n574) );
  HS65_LS_NOR2X19 U98 ( .A(n463), .B(n464), .Z(n105) );
  HS65_LH_MUX21I1X3 U99 ( .D0(n25), .D1(n452), .S0(n648), .Z(n683) );
  HS65_LS_IVX18 U100 ( .A(n112), .Z(n118) );
  HS65_LS_IVX9 U101 ( .A(n113), .Z(n30) );
  HS65_LS_OAI212X3 U102 ( .A(n117), .B(n475), .C(n526), .D(n474), .E(n473), 
        .Z(pkt_out[2]) );
  HS65_LS_OAI212X3 U103 ( .A(n117), .B(n471), .C(n526), .D(n470), .E(n469), 
        .Z(pkt_out[1]) );
  HS65_LS_BFX9 U104 ( .A(n331), .Z(n327) );
  HS65_LS_BFX9 U105 ( .A(n331), .Z(n326) );
  HS65_LS_BFX9 U106 ( .A(n312), .Z(n303) );
  HS65_LS_BFX9 U107 ( .A(n312), .Z(n304) );
  HS65_LS_BFX9 U108 ( .A(n294), .Z(n297) );
  HS65_LS_BFX9 U109 ( .A(n336), .Z(n354) );
  HS65_LS_BFX9 U110 ( .A(n335), .Z(n353) );
  HS65_LS_BFX9 U111 ( .A(n335), .Z(n352) );
  HS65_LH_MUXI21X2 U112 ( .D0(n455), .D1(n108), .S0(n648), .Z(n677) );
  HS65_LS_NAND2X2 U113 ( .A(state_cnt[1]), .B(n445), .Z(n448) );
  HS65_LH_NAND2X2 U114 ( .A(state_cnt[1]), .B(n445), .Z(n37) );
  HS65_LS_OAI212X3 U115 ( .A(n116), .B(n502), .C(n526), .D(n501), .E(n500), 
        .Z(pkt_out[11]) );
  HS65_LS_OAI212X3 U116 ( .A(n117), .B(n499), .C(n526), .D(n498), .E(n497), 
        .Z(pkt_out[10]) );
  HS65_LS_OAI212X3 U117 ( .A(n116), .B(n478), .C(n526), .D(n477), .E(n476), 
        .Z(pkt_out[3]) );
  HS65_LS_IVX9 U118 ( .A(n327), .Z(n313) );
  HS65_LS_IVX9 U119 ( .A(n327), .Z(n314) );
  HS65_LS_IVX9 U120 ( .A(n326), .Z(n323) );
  HS65_LS_IVX9 U121 ( .A(n326), .Z(n324) );
  HS65_LS_IVX9 U122 ( .A(n326), .Z(n325) );
  HS65_LS_AND2X4 U123 ( .A(n615), .B(n614), .Z(n39) );
  HS65_LS_AND2X4 U124 ( .A(n601), .B(n72), .Z(n41) );
  HS65_LS_AND2X4 U125 ( .A(n602), .B(n41), .Z(n42) );
  HS65_LS_AND2X4 U126 ( .A(n603), .B(n42), .Z(n43) );
  HS65_LS_AND2X4 U127 ( .A(n604), .B(n43), .Z(n44) );
  HS65_LS_AND2X4 U128 ( .A(n605), .B(n44), .Z(n45) );
  HS65_LS_AND2X4 U129 ( .A(n606), .B(n45), .Z(n46) );
  HS65_LS_AND2X4 U130 ( .A(n607), .B(n46), .Z(n47) );
  HS65_LS_AND2X4 U131 ( .A(n608), .B(n47), .Z(n48) );
  HS65_LS_AND2X4 U132 ( .A(n609), .B(n48), .Z(n49) );
  HS65_LS_AND2X4 U133 ( .A(n610), .B(n49), .Z(n50) );
  HS65_LS_AND2X4 U134 ( .A(n611), .B(n50), .Z(n51) );
  HS65_LS_AND2X4 U135 ( .A(n620), .B(n73), .Z(n52) );
  HS65_LS_AND2X4 U136 ( .A(n616), .B(n39), .Z(n53) );
  HS65_LS_AND2X4 U137 ( .A(n617), .B(n53), .Z(n54) );
  HS65_LS_AND2X4 U138 ( .A(n618), .B(n54), .Z(n55) );
  HS65_LS_AND2X4 U139 ( .A(\add_545/A[8] ), .B(n52), .Z(n56) );
  HS65_LS_AND2X4 U140 ( .A(\add_545/A[9] ), .B(n56), .Z(n57) );
  HS65_LS_AND2X4 U141 ( .A(\add_545/A[10] ), .B(n57), .Z(n58) );
  HS65_LS_AND2X4 U142 ( .A(\add_545/A[11] ), .B(n58), .Z(n59) );
  HS65_LS_AND2X4 U143 ( .A(\add_545/A[12] ), .B(n59), .Z(n62) );
  HS65_LS_AND2X4 U144 ( .A(\add_545/A[13] ), .B(n62), .Z(n64) );
  HS65_LS_AND2X4 U145 ( .A(n600), .B(n599), .Z(n72) );
  HS65_LS_AND2X4 U146 ( .A(n619), .B(n55), .Z(n73) );
  HS65_LS_BFX9 U147 ( .A(n330), .Z(n328) );
  HS65_LS_BFX9 U148 ( .A(n330), .Z(n329) );
  HS65_LS_IVX9 U149 ( .A(n303), .Z(n302) );
  HS65_LS_IVX9 U150 ( .A(n304), .Z(n301) );
  HS65_LS_IVX9 U151 ( .A(n304), .Z(n300) );
  HS65_LS_OAI21X3 U152 ( .A(n867), .B(n855), .C(n313), .Z(dma_wen[2]) );
  HS65_LS_NOR2AX3 U153 ( .A(n853), .B(n597), .Z(n867) );
  HS65_LS_IVX9 U154 ( .A(n851), .Z(n597) );
  HS65_LSS_XNOR2X6 U155 ( .A(n93), .B(\sub_544/A[10] ), .Z(dma_cnt_new[10]) );
  HS65_LSS_XNOR2X6 U156 ( .A(n87), .B(\sub_544/A[5] ), .Z(dma_cnt_new[5]) );
  HS65_LSS_XNOR2X6 U157 ( .A(n91), .B(\sub_544/A[9] ), .Z(dma_cnt_new[9]) );
  HS65_LSS_XNOR2X6 U158 ( .A(n84), .B(\sub_544/A[4] ), .Z(dma_cnt_new[4]) );
  HS65_LSS_XNOR2X6 U159 ( .A(n90), .B(\sub_544/A[8] ), .Z(dma_cnt_new[8]) );
  HS65_LS_NOR4ABX2 U160 ( .A(n101), .B(n102), .C(n863), .D(dma_cnt_new[13]), 
        .Z(n845) );
  HS65_LSS_XOR2X6 U161 ( .A(n89), .B(\sub_544/A[7] ), .Z(n75) );
  HS65_LSS_XOR2X6 U162 ( .A(n80), .B(\sub_544/A[3] ), .Z(n77) );
  HS65_LSS_XOR2X6 U163 ( .A(n88), .B(\sub_544/A[6] ), .Z(n78) );
  HS65_LS_IVX9 U164 ( .A(n877), .Z(\add_545/A[8] ) );
  HS65_LS_IVX9 U165 ( .A(n878), .Z(\add_545/A[9] ) );
  HS65_LS_IVX9 U166 ( .A(n879), .Z(\add_545/A[10] ) );
  HS65_LS_IVX9 U167 ( .A(n872), .Z(\add_545/A[11] ) );
  HS65_LS_IVX9 U168 ( .A(n873), .Z(\add_545/A[12] ) );
  HS65_LS_IVX9 U169 ( .A(n874), .Z(\add_545/A[13] ) );
  HS65_LS_IVX9 U170 ( .A(n875), .Z(\add_545/A[14] ) );
  HS65_LS_BFX9 U171 ( .A(n103), .Z(n330) );
  HS65_LS_BFX9 U172 ( .A(n103), .Z(n331) );
  HS65_LSS_XOR2X6 U173 ( .A(\sub_544/A[1] ), .B(\sub_544/A[2] ), .Z(n79) );
  HS65_LS_OR2X9 U174 ( .A(\sub_544/A[2] ), .B(\sub_544/A[1] ), .Z(n80) );
  HS65_LS_OR2X9 U175 ( .A(\sub_544/A[3] ), .B(n80), .Z(n84) );
  HS65_LS_OR2X9 U176 ( .A(\sub_544/A[4] ), .B(n84), .Z(n87) );
  HS65_LS_OR2X9 U177 ( .A(\sub_544/A[5] ), .B(n87), .Z(n88) );
  HS65_LS_OR2X9 U178 ( .A(\sub_544/A[6] ), .B(n88), .Z(n89) );
  HS65_LS_OR2X9 U179 ( .A(\sub_544/A[7] ), .B(n89), .Z(n90) );
  HS65_LS_OR2X9 U180 ( .A(\sub_544/A[8] ), .B(n90), .Z(n91) );
  HS65_LS_OR2X9 U181 ( .A(\sub_544/A[9] ), .B(n91), .Z(n93) );
  HS65_LS_OR2X9 U182 ( .A(\sub_544/A[10] ), .B(n93), .Z(n94) );
  HS65_LS_OR2X9 U183 ( .A(\sub_544/A[11] ), .B(n94), .Z(n95) );
  HS65_LSS_XOR2X6 U184 ( .A(n94), .B(\sub_544/A[11] ), .Z(n101) );
  HS65_LSS_XOR2X6 U185 ( .A(n95), .B(\sub_544/A[12] ), .Z(n102) );
  HS65_LS_BFX9 U186 ( .A(n621), .Z(n138) );
  HS65_LS_BFX9 U187 ( .A(n621), .Z(n139) );
  HS65_LS_BFX9 U188 ( .A(n142), .Z(n149) );
  HS65_LS_BFX9 U189 ( .A(n142), .Z(n144) );
  HS65_LS_BFX9 U190 ( .A(n621), .Z(n140) );
  HS65_LS_BFX9 U191 ( .A(n142), .Z(n293) );
  HS65_LS_IVX9 U192 ( .A(n297), .Z(n295) );
  HS65_LS_IVX9 U193 ( .A(n297), .Z(n296) );
  HS65_LS_BFX9 U194 ( .A(n312), .Z(n305) );
  HS65_LS_BFX9 U195 ( .A(n312), .Z(n310) );
  HS65_LS_BFX9 U196 ( .A(n312), .Z(n306) );
  HS65_LS_BFX9 U197 ( .A(n312), .Z(n311) );
  HS65_LS_BFX9 U198 ( .A(n128), .Z(n129) );
  HS65_LS_BFX9 U199 ( .A(n128), .Z(n130) );
  HS65_LS_BFX9 U200 ( .A(n4), .Z(n124) );
  HS65_LS_BFX9 U201 ( .A(n4), .Z(n125) );
  HS65_LS_BFX9 U202 ( .A(n128), .Z(n132) );
  HS65_LS_BFX9 U203 ( .A(n4), .Z(n127) );
  HS65_LS_IVX9 U204 ( .A(n855), .Z(n653) );
  HS65_LS_IVX9 U205 ( .A(\proc_out[SRESP] ), .Z(n332) );
  HS65_LS_IVX9 U206 ( .A(n354), .Z(n345) );
  HS65_LS_IVX9 U207 ( .A(n354), .Z(n344) );
  HS65_LS_IVX9 U208 ( .A(n354), .Z(n348) );
  HS65_LS_IVX9 U209 ( .A(n354), .Z(n347) );
  HS65_LS_IVX9 U210 ( .A(n354), .Z(n346) );
  HS65_LS_IVX9 U211 ( .A(n353), .Z(n343) );
  HS65_LS_IVX9 U212 ( .A(n353), .Z(n342) );
  HS65_LS_IVX9 U213 ( .A(n353), .Z(n340) );
  HS65_LS_IVX9 U214 ( .A(n353), .Z(n339) );
  HS65_LS_IVX9 U215 ( .A(n353), .Z(n338) );
  HS65_LS_IVX9 U216 ( .A(n353), .Z(n341) );
  HS65_LS_IVX9 U217 ( .A(n355), .Z(n351) );
  HS65_LS_IVX9 U218 ( .A(n355), .Z(n350) );
  HS65_LS_IVX9 U219 ( .A(n355), .Z(n349) );
  HS65_LS_IVX9 U220 ( .A(n352), .Z(n337) );
  HS65_LS_NOR2X6 U221 ( .A(n355), .B(n877), .Z(\spm_out[MADDR][7] ) );
  HS65_LS_NOR2X6 U222 ( .A(n355), .B(n878), .Z(\spm_out[MADDR][8] ) );
  HS65_LS_NOR2X6 U223 ( .A(n355), .B(n879), .Z(\spm_out[MADDR][9] ) );
  HS65_LS_NOR2X6 U224 ( .A(n355), .B(n872), .Z(\spm_out[MADDR][10] ) );
  HS65_LS_NOR2X6 U225 ( .A(n355), .B(n873), .Z(\spm_out[MADDR][11] ) );
  HS65_LS_NOR2X6 U226 ( .A(n355), .B(n874), .Z(\spm_out[MADDR][12] ) );
  HS65_LS_NOR2X6 U227 ( .A(n355), .B(n875), .Z(\spm_out[MADDR][13] ) );
  HS65_LS_NOR2X6 U228 ( .A(n355), .B(n876), .Z(\spm_out[MADDR][14] ) );
  HS65_LS_NOR2X6 U229 ( .A(n332), .B(n643), .Z(\proc_out[SDATA][0] ) );
  HS65_LS_NOR2X6 U230 ( .A(n332), .B(n642), .Z(\proc_out[SDATA][1] ) );
  HS65_LS_NOR2X6 U231 ( .A(n332), .B(n641), .Z(\proc_out[SDATA][2] ) );
  HS65_LS_NOR2X6 U232 ( .A(n871), .B(n640), .Z(\proc_out[SDATA][3] ) );
  HS65_LS_NOR2X6 U233 ( .A(n332), .B(n639), .Z(\proc_out[SDATA][4] ) );
  HS65_LS_NOR2X6 U234 ( .A(n871), .B(n638), .Z(\proc_out[SDATA][5] ) );
  HS65_LS_NOR2X6 U235 ( .A(n871), .B(n637), .Z(\proc_out[SDATA][6] ) );
  HS65_LS_NOR2X6 U236 ( .A(n871), .B(n636), .Z(\proc_out[SDATA][7] ) );
  HS65_LS_NOR2X6 U237 ( .A(n332), .B(n635), .Z(\proc_out[SDATA][8] ) );
  HS65_LS_NOR2X6 U238 ( .A(n332), .B(n634), .Z(\proc_out[SDATA][9] ) );
  HS65_LS_NOR2X6 U239 ( .A(n332), .B(n633), .Z(\proc_out[SDATA][10] ) );
  HS65_LS_NOR2X6 U240 ( .A(n332), .B(n632), .Z(\proc_out[SDATA][11] ) );
  HS65_LS_NOR2X6 U241 ( .A(n332), .B(n631), .Z(\proc_out[SDATA][12] ) );
  HS65_LS_NOR2X6 U242 ( .A(n332), .B(n630), .Z(\proc_out[SDATA][13] ) );
  HS65_LS_NOR2X6 U243 ( .A(n332), .B(n629), .Z(\proc_out[SDATA][14] ) );
  HS65_LS_NOR2X6 U244 ( .A(n332), .B(n628), .Z(\proc_out[SDATA][15] ) );
  HS65_LS_AND3X9 U245 ( .A(dma_rdata[63]), .B(n645), .C(n140), .Z(n103) );
  HS65_LS_OAI222X2 U246 ( .A(n327), .B(n837), .C(n850), .D(n675), .E(n313), 
        .F(n837), .Z(dma_wdata[48]) );
  HS65_LS_NOR2X6 U247 ( .A(n867), .B(n854), .Z(dma_wen[0]) );
  HS65_LS_OAI222X2 U248 ( .A(n327), .B(n838), .C(n850), .D(n672), .E(n313), 
        .F(n77), .Z(dma_wdata[51]) );
  HS65_LS_OAI222X2 U249 ( .A(n327), .B(n839), .C(n850), .D(n671), .E(n313), 
        .F(n627), .Z(dma_wdata[52]) );
  HS65_LS_IVX9 U250 ( .A(dma_cnt_new[4]), .Z(n627) );
  HS65_LS_OAI222X2 U251 ( .A(n327), .B(n840), .C(n668), .D(n850), .E(n313), 
        .F(n75), .Z(dma_wdata[55]) );
  HS65_LS_OAI222X2 U252 ( .A(n327), .B(n841), .C(n667), .D(n850), .E(n313), 
        .F(n625), .Z(dma_wdata[56]) );
  HS65_LS_IVX9 U253 ( .A(dma_cnt_new[8]), .Z(n625) );
  HS65_LS_OAI222X2 U254 ( .A(n327), .B(n842), .C(n850), .D(n665), .E(n314), 
        .F(n623), .Z(dma_wdata[58]) );
  HS65_LS_IVX9 U255 ( .A(dma_cnt_new[10]), .Z(n623) );
  HS65_LS_OAI222X2 U256 ( .A(n326), .B(n843), .C(n850), .D(n663), .E(n314), 
        .F(n102), .Z(dma_wdata[60]) );
  HS65_LS_OAI222X2 U257 ( .A(n327), .B(n844), .C(n850), .D(n662), .E(n313), 
        .F(n622), .Z(dma_wdata[61]) );
  HS65_LS_IVX9 U258 ( .A(dma_cnt_new[13]), .Z(n622) );
  HS65_LS_OAI222X2 U259 ( .A(n327), .B(n863), .C(n850), .D(n674), .E(n313), 
        .F(\sub_544/A[1] ), .Z(dma_wdata[49]) );
  HS65_LS_OAI222X2 U260 ( .A(n327), .B(n862), .C(n850), .D(n673), .E(n313), 
        .F(n79), .Z(dma_wdata[50]) );
  HS65_LS_OAI222X2 U261 ( .A(n327), .B(n861), .C(n850), .D(n670), .E(n313), 
        .F(n626), .Z(dma_wdata[53]) );
  HS65_LS_IVX9 U262 ( .A(dma_cnt_new[5]), .Z(n626) );
  HS65_LS_OAI222X2 U263 ( .A(n327), .B(n860), .C(n669), .D(n850), .E(n313), 
        .F(n78), .Z(dma_wdata[54]) );
  HS65_LS_OAI222X2 U264 ( .A(n327), .B(n859), .C(n666), .D(n850), .E(n313), 
        .F(n624), .Z(dma_wdata[57]) );
  HS65_LS_IVX9 U265 ( .A(dma_cnt_new[9]), .Z(n624) );
  HS65_LS_OAI222X2 U266 ( .A(n327), .B(n858), .C(n850), .D(n664), .E(n313), 
        .F(n101), .Z(dma_wdata[59]) );
  HS65_LS_OAI212X5 U267 ( .A(n850), .B(n661), .C(n852), .D(n645), .E(n849), 
        .Z(dma_wdata[62]) );
  HS65_LS_NAND4ABX3 U268 ( .A(n848), .B(n847), .C(n846), .D(n845), .Z(n849) );
  HS65_LS_NAND4ABX3 U269 ( .A(dma_cnt_new[5]), .B(dma_cnt_new[4]), .C(n79), 
        .D(n77), .Z(n847) );
  HS65_LS_NAND4ABX3 U270 ( .A(dma_cnt_new[9]), .B(dma_cnt_new[8]), .C(n78), 
        .D(n75), .Z(n848) );
  HS65_LS_NAND2X7 U271 ( .A(n652), .B(n1), .Z(n851) );
  HS65_LS_OAI21X3 U272 ( .A(n867), .B(n857), .C(n313), .Z(dma_wen[1]) );
  HS65_LS_NAND2X7 U273 ( .A(n362), .B(n361), .Z(n593) );
  HS65_LSS_XNOR2X6 U274 ( .A(n844), .B(n111), .Z(dma_cnt_new[13]) );
  HS65_LS_NOR2X6 U275 ( .A(\sub_544/A[12] ), .B(n95), .Z(n111) );
  HS65_LS_NOR3X4 U276 ( .A(n313), .B(dma_cnt_new[10]), .C(dma_cnt_new[0]), .Z(
        n846) );
  HS65_LS_IVX9 U277 ( .A(n837), .Z(dma_cnt_new[0]) );
  HS65_LS_IVX9 U278 ( .A(n863), .Z(\sub_544/A[1] ) );
  HS65_LS_NAND2X7 U279 ( .A(dma_rdata[40]), .B(n138), .Z(n877) );
  HS65_LS_NAND2X7 U280 ( .A(dma_rdata[41]), .B(n138), .Z(n878) );
  HS65_LS_NAND2X7 U281 ( .A(dma_rdata[42]), .B(n138), .Z(n879) );
  HS65_LS_NAND2X7 U282 ( .A(dma_rdata[43]), .B(n138), .Z(n872) );
  HS65_LS_NAND2X7 U283 ( .A(dma_rdata[44]), .B(n138), .Z(n873) );
  HS65_LS_NAND2X7 U284 ( .A(dma_rdata[45]), .B(n139), .Z(n874) );
  HS65_LS_NAND2X7 U285 ( .A(dma_rdata[46]), .B(n139), .Z(n875) );
  HS65_LS_IVX9 U286 ( .A(n838), .Z(\sub_544/A[3] ) );
  HS65_LS_IVX9 U287 ( .A(n839), .Z(\sub_544/A[4] ) );
  HS65_LS_IVX9 U288 ( .A(n840), .Z(\sub_544/A[7] ) );
  HS65_LS_IVX9 U289 ( .A(n841), .Z(\sub_544/A[8] ) );
  HS65_LS_IVX9 U290 ( .A(n842), .Z(\sub_544/A[10] ) );
  HS65_LS_IVX9 U291 ( .A(n843), .Z(\sub_544/A[12] ) );
  HS65_LS_IVX9 U292 ( .A(n862), .Z(\sub_544/A[2] ) );
  HS65_LS_IVX9 U293 ( .A(n861), .Z(\sub_544/A[5] ) );
  HS65_LS_IVX9 U294 ( .A(n860), .Z(\sub_544/A[6] ) );
  HS65_LS_IVX9 U295 ( .A(n859), .Z(\sub_544/A[9] ) );
  HS65_LS_IVX9 U296 ( .A(n858), .Z(\sub_544/A[11] ) );
  HS65_LS_BFX9 U297 ( .A(n836), .Z(n142) );
  HS65_LS_NOR2AX3 U298 ( .A(n1), .B(n857), .Z(n836) );
  HS65_LS_OAI22X6 U299 ( .A(n852), .B(n644), .C(n850), .D(n660), .Z(
        dma_wdata[63]) );
  HS65_LS_IVX9 U300 ( .A(dma_rdata[63]), .Z(n644) );
  HS65_LS_OAI22X6 U301 ( .A(n852), .B(n643), .C(n851), .D(n675), .Z(
        dma_wdata[0]) );
  HS65_LS_OAI22X6 U302 ( .A(n852), .B(n642), .C(n851), .D(n674), .Z(
        dma_wdata[1]) );
  HS65_LS_OAI22X6 U303 ( .A(n852), .B(n641), .C(n851), .D(n673), .Z(
        dma_wdata[2]) );
  HS65_LS_OAI22X6 U304 ( .A(n852), .B(n640), .C(n851), .D(n672), .Z(
        dma_wdata[3]) );
  HS65_LS_OAI22X6 U305 ( .A(n852), .B(n639), .C(n851), .D(n671), .Z(
        dma_wdata[4]) );
  HS65_LS_OAI22X6 U306 ( .A(n852), .B(n638), .C(n851), .D(n670), .Z(
        dma_wdata[5]) );
  HS65_LS_OAI22X6 U307 ( .A(n852), .B(n637), .C(n851), .D(n669), .Z(
        dma_wdata[6]) );
  HS65_LS_OAI22X6 U308 ( .A(n852), .B(n636), .C(n851), .D(n668), .Z(
        dma_wdata[7]) );
  HS65_LS_OAI22X6 U309 ( .A(n852), .B(n635), .C(n851), .D(n667), .Z(
        dma_wdata[8]) );
  HS65_LS_OAI22X6 U310 ( .A(n852), .B(n634), .C(n851), .D(n666), .Z(
        dma_wdata[9]) );
  HS65_LS_OAI22X6 U311 ( .A(n852), .B(n633), .C(n851), .D(n665), .Z(
        dma_wdata[10]) );
  HS65_LS_OAI22X6 U312 ( .A(n852), .B(n632), .C(n851), .D(n664), .Z(
        dma_wdata[11]) );
  HS65_LS_OAI22X6 U313 ( .A(n852), .B(n631), .C(n851), .D(n663), .Z(
        dma_wdata[12]) );
  HS65_LS_OAI22X6 U314 ( .A(n852), .B(n630), .C(n851), .D(n662), .Z(
        dma_wdata[13]) );
  HS65_LS_OAI22X6 U315 ( .A(n852), .B(n629), .C(n851), .D(n661), .Z(
        dma_wdata[14]) );
  HS65_LS_OAI22X6 U316 ( .A(n852), .B(n628), .C(n851), .D(n660), .Z(
        dma_wdata[15]) );
  HS65_LS_OAI21X3 U317 ( .A(n652), .B(n835), .C(n357), .Z(n594) );
  HS65_LH_OAI21X2 U318 ( .A(n854), .B(n594), .C(n362), .Z(dma_ren[0]) );
  HS65_LH_OAI21X2 U319 ( .A(n857), .B(n594), .C(n362), .Z(dma_ren[1]) );
  HS65_LH_OAI21X2 U320 ( .A(n855), .B(n594), .C(n362), .Z(dma_ren[2]) );
  HS65_LS_NAND2X7 U321 ( .A(n653), .B(n1), .Z(n850) );
  HS65_LS_IVX9 U322 ( .A(n864), .Z(n649) );
  HS65_LS_NAND2X7 U323 ( .A(dma_rdata[47]), .B(n139), .Z(n876) );
  HS65_LS_IVX9 U324 ( .A(dma_rdata[0]), .Z(n643) );
  HS65_LS_IVX9 U325 ( .A(dma_rdata[1]), .Z(n642) );
  HS65_LS_IVX9 U326 ( .A(dma_rdata[2]), .Z(n641) );
  HS65_LS_IVX9 U327 ( .A(dma_rdata[3]), .Z(n640) );
  HS65_LS_IVX9 U328 ( .A(dma_rdata[4]), .Z(n639) );
  HS65_LS_IVX9 U329 ( .A(dma_rdata[5]), .Z(n638) );
  HS65_LS_IVX9 U330 ( .A(dma_rdata[6]), .Z(n637) );
  HS65_LS_IVX9 U331 ( .A(dma_rdata[7]), .Z(n636) );
  HS65_LS_IVX9 U332 ( .A(dma_rdata[8]), .Z(n635) );
  HS65_LS_IVX9 U333 ( .A(dma_rdata[9]), .Z(n634) );
  HS65_LS_IVX9 U334 ( .A(dma_rdata[10]), .Z(n633) );
  HS65_LS_IVX9 U335 ( .A(dma_rdata[11]), .Z(n632) );
  HS65_LS_IVX9 U336 ( .A(dma_rdata[12]), .Z(n631) );
  HS65_LS_IVX9 U337 ( .A(dma_rdata[13]), .Z(n630) );
  HS65_LS_IVX9 U338 ( .A(dma_rdata[14]), .Z(n629) );
  HS65_LS_IVX9 U339 ( .A(dma_rdata[15]), .Z(n628) );
  HS65_LS_BFX9 U340 ( .A(n411), .Z(n128) );
  HS65_LS_BFX9 U341 ( .A(n294), .Z(n298) );
  HS65_LS_IVX9 U342 ( .A(n866), .Z(n312) );
  HS65_LS_BFX9 U343 ( .A(n294), .Z(n299) );
  HS65_LS_NAND3X5 U344 ( .A(n137), .B(n577), .C(n337), .Z(n592) );
  HS65_LS_IVX9 U345 ( .A(n854), .Z(n652) );
  HS65_LS_NAND2X7 U346 ( .A(n855), .B(n857), .Z(n835) );
  HS65_LS_NAND2X7 U347 ( .A(n832), .B(n659), .Z(n855) );
  HS65_LS_BFX9 U348 ( .A(n334), .Z(\proc_out[SRESP] ) );
  HS65_LS_IVX9 U349 ( .A(n871), .Z(n334) );
  HS65_LS_BFX9 U350 ( .A(n336), .Z(n355) );
  HS65_LS_IVX9 U351 ( .A(n868), .Z(n651) );
  HS65_LS_NOR2AX3 U352 ( .A(dma_rdata[16]), .B(n871), .Z(\proc_out[SDATA][16] ) );
  HS65_LS_NOR2AX3 U353 ( .A(dma_rdata[17]), .B(n871), .Z(\proc_out[SDATA][17] ) );
  HS65_LS_NOR2AX3 U354 ( .A(dma_rdata[18]), .B(n871), .Z(\proc_out[SDATA][18] ) );
  HS65_LS_NOR2AX3 U355 ( .A(dma_rdata[19]), .B(n871), .Z(\proc_out[SDATA][19] ) );
  HS65_LS_NOR2AX3 U356 ( .A(dma_rdata[20]), .B(n871), .Z(\proc_out[SDATA][20] ) );
  HS65_LS_NOR2AX3 U357 ( .A(dma_rdata[21]), .B(n871), .Z(\proc_out[SDATA][21] ) );
  HS65_LS_NOR2AX3 U358 ( .A(dma_rdata[22]), .B(n871), .Z(\proc_out[SDATA][22] ) );
  HS65_LS_NOR2AX3 U359 ( .A(dma_rdata[23]), .B(n871), .Z(\proc_out[SDATA][23] ) );
  HS65_LS_NOR2AX3 U360 ( .A(dma_rdata[24]), .B(n871), .Z(\proc_out[SDATA][24] ) );
  HS65_LS_NOR2AX3 U361 ( .A(dma_rdata[25]), .B(n871), .Z(\proc_out[SDATA][25] ) );
  HS65_LS_NOR2AX3 U362 ( .A(dma_rdata[26]), .B(n332), .Z(\proc_out[SDATA][26] ) );
  HS65_LS_NOR2AX3 U363 ( .A(dma_rdata[27]), .B(n871), .Z(\proc_out[SDATA][27] ) );
  HS65_LS_NOR2AX3 U364 ( .A(dma_rdata[28]), .B(n871), .Z(\proc_out[SDATA][28] ) );
  HS65_LS_NOR2AX3 U365 ( .A(dma_rdata[29]), .B(n332), .Z(\proc_out[SDATA][29] ) );
  HS65_LS_NOR2AX3 U366 ( .A(dma_rdata[30]), .B(n871), .Z(\proc_out[SDATA][30] ) );
  HS65_LS_NOR2AX3 U367 ( .A(dma_rdata[31]), .B(n871), .Z(\proc_out[SDATA][31] ) );
  HS65_LS_IVX9 U368 ( .A(n857), .Z(n654) );
  HS65_LS_AOI22X6 U369 ( .A(\proc_in[MADDR][1] ), .B(n652), .C(
        \proc_in[MADDR][2] ), .D(n835), .Z(n834) );
  HS65_LS_AOI22X6 U370 ( .A(\proc_in[MADDR][0] ), .B(n652), .C(
        \proc_in[MADDR][1] ), .D(n835), .Z(n833) );
  HS65_LS_IVX9 U371 ( .A(\proc_in[MADDR][2] ), .Z(n657) );
  HS65_LS_NAND2X7 U372 ( .A(slt_entry[4]), .B(n648), .Z(n852) );
  HS65_LS_OAI21X3 U373 ( .A(n648), .B(n133), .C(n356), .Z(n358) );
  HS65_LH_MUXI21X2 U374 ( .D0(n686), .D1(n106), .S0(n648), .Z(n678) );
  HS65_LS_NOR2X6 U375 ( .A(slt_entry[0]), .B(n323), .Z(n106) );
  HS65_LS_NOR2X6 U376 ( .A(slt_entry[1]), .B(n323), .Z(n108) );
  HS65_LS_OAI21X3 U377 ( .A(n685), .B(n648), .C(n323), .Z(n679) );
  HS65_LS_MX41X7 U378 ( .D0(n596), .S0(n328), .D1(n596), .S1(n314), .D2(
        \proc_in[MDATA][16] ), .S2(n597), .D3(n144), .S3(\proc_in[MDATA][0] ), 
        .Z(dma_wdata[16]) );
  HS65_LS_MX41X7 U379 ( .D0(n382), .S0(n327), .D1(n599), .S1(n314), .D2(
        \proc_in[MDATA][17] ), .S2(n597), .D3(n144), .S3(\proc_in[MDATA][1] ), 
        .Z(dma_wdata[17]) );
  HS65_LS_MX41X7 U380 ( .D0(dma_wp_new[2]), .S0(n327), .D1(n600), .S1(n314), 
        .D2(\proc_in[MDATA][18] ), .S2(n597), .D3(n144), .S3(
        \proc_in[MDATA][2] ), .Z(dma_wdata[18]) );
  HS65_LSS_XOR2X6 U381 ( .A(n599), .B(n600), .Z(dma_wp_new[2]) );
  HS65_LS_MX41X7 U382 ( .D0(dma_wp_new[3]), .S0(n327), .D1(n601), .S1(n314), 
        .D2(\proc_in[MDATA][19] ), .S2(n597), .D3(n144), .S3(
        \proc_in[MDATA][3] ), .Z(dma_wdata[19]) );
  HS65_LSS_XOR2X6 U383 ( .A(n72), .B(n601), .Z(dma_wp_new[3]) );
  HS65_LS_MX41X7 U384 ( .D0(dma_wp_new[4]), .S0(n327), .D1(n602), .S1(n314), 
        .D2(\proc_in[MDATA][20] ), .S2(n597), .D3(n144), .S3(
        \proc_in[MDATA][4] ), .Z(dma_wdata[20]) );
  HS65_LSS_XOR2X6 U385 ( .A(n41), .B(n602), .Z(dma_wp_new[4]) );
  HS65_LS_MX41X7 U386 ( .D0(dma_wp_new[5]), .S0(n327), .D1(n603), .S1(n314), 
        .D2(\proc_in[MDATA][21] ), .S2(n597), .D3(n144), .S3(
        \proc_in[MDATA][5] ), .Z(dma_wdata[21]) );
  HS65_LSS_XOR2X6 U387 ( .A(n42), .B(n603), .Z(dma_wp_new[5]) );
  HS65_LS_MX41X7 U388 ( .D0(dma_wp_new[6]), .S0(n328), .D1(n604), .S1(n314), 
        .D2(\proc_in[MDATA][22] ), .S2(n597), .D3(n144), .S3(
        \proc_in[MDATA][6] ), .Z(dma_wdata[22]) );
  HS65_LSS_XOR2X6 U389 ( .A(n43), .B(n604), .Z(dma_wp_new[6]) );
  HS65_LS_MX41X7 U390 ( .D0(dma_wp_new[7]), .S0(n328), .D1(n605), .S1(n314), 
        .D2(\proc_in[MDATA][23] ), .S2(n597), .D3(n144), .S3(
        \proc_in[MDATA][7] ), .Z(dma_wdata[23]) );
  HS65_LSS_XOR2X6 U391 ( .A(n44), .B(n605), .Z(dma_wp_new[7]) );
  HS65_LS_MX41X7 U392 ( .D0(dma_wp_new[8]), .S0(n328), .D1(n606), .S1(n314), 
        .D2(\proc_in[MDATA][24] ), .S2(n597), .D3(n144), .S3(
        \proc_in[MDATA][8] ), .Z(dma_wdata[24]) );
  HS65_LSS_XOR2X6 U393 ( .A(n45), .B(n606), .Z(dma_wp_new[8]) );
  HS65_LS_MX41X7 U394 ( .D0(dma_wp_new[9]), .S0(n328), .D1(n607), .S1(n314), 
        .D2(\proc_in[MDATA][25] ), .S2(n597), .D3(n144), .S3(
        \proc_in[MDATA][9] ), .Z(dma_wdata[25]) );
  HS65_LSS_XOR2X6 U395 ( .A(n46), .B(n607), .Z(dma_wp_new[9]) );
  HS65_LS_MX41X7 U396 ( .D0(dma_wp_new[10]), .S0(n328), .D1(n608), .S1(n314), 
        .D2(\proc_in[MDATA][26] ), .S2(n597), .D3(n144), .S3(
        \proc_in[MDATA][10] ), .Z(dma_wdata[26]) );
  HS65_LSS_XOR2X6 U397 ( .A(n47), .B(n608), .Z(dma_wp_new[10]) );
  HS65_LS_MX41X7 U398 ( .D0(dma_wp_new[11]), .S0(n328), .D1(n609), .S1(n314), 
        .D2(\proc_in[MDATA][27] ), .S2(n597), .D3(n144), .S3(
        \proc_in[MDATA][11] ), .Z(dma_wdata[27]) );
  HS65_LSS_XOR2X6 U399 ( .A(n48), .B(n609), .Z(dma_wp_new[11]) );
  HS65_LS_MX41X7 U400 ( .D0(dma_wp_new[12]), .S0(n328), .D1(n610), .S1(n314), 
        .D2(\proc_in[MDATA][28] ), .S2(n597), .D3(n149), .S3(
        \proc_in[MDATA][12] ), .Z(dma_wdata[28]) );
  HS65_LSS_XOR2X6 U401 ( .A(n49), .B(n610), .Z(dma_wp_new[12]) );
  HS65_LS_MX41X7 U402 ( .D0(dma_wp_new[13]), .S0(n328), .D1(n611), .S1(n314), 
        .D2(\proc_in[MDATA][29] ), .S2(n597), .D3(n149), .S3(
        \proc_in[MDATA][13] ), .Z(dma_wdata[29]) );
  HS65_LSS_XOR2X6 U403 ( .A(n50), .B(n611), .Z(dma_wp_new[13]) );
  HS65_LS_MX41X7 U404 ( .D0(dma_wp_new[14]), .S0(n328), .D1(n612), .S1(n314), 
        .D2(\proc_in[MDATA][30] ), .S2(n597), .D3(n149), .S3(
        \proc_in[MDATA][14] ), .Z(dma_wdata[30]) );
  HS65_LSS_XOR2X6 U405 ( .A(n51), .B(n612), .Z(dma_wp_new[14]) );
  HS65_LS_MX41X7 U406 ( .D0(dma_wp_new[15]), .S0(n328), .D1(n613), .S1(n314), 
        .D2(\proc_in[MDATA][31] ), .S2(n597), .D3(n149), .S3(
        \proc_in[MDATA][15] ), .Z(dma_wdata[31]) );
  HS65_LSS_XOR2X6 U407 ( .A(n613), .B(n2), .Z(dma_wp_new[15]) );
  HS65_LS_AO222X4 U408 ( .A(n614), .B(n323), .C(\proc_in[MDATA][17] ), .D(n149), .E(n579), .F(n328), .Z(dma_wdata[33]) );
  HS65_LS_AO222X4 U409 ( .A(n615), .B(n323), .C(\proc_in[MDATA][18] ), .D(n149), .E(dma_rp_new[2]), .F(n328), .Z(dma_wdata[34]) );
  HS65_LSS_XOR2X6 U410 ( .A(n614), .B(n615), .Z(dma_rp_new[2]) );
  HS65_LS_AO222X4 U411 ( .A(n616), .B(n323), .C(\proc_in[MDATA][19] ), .D(n149), .E(dma_rp_new[3]), .F(n328), .Z(dma_wdata[35]) );
  HS65_LSS_XOR2X6 U412 ( .A(n39), .B(n616), .Z(dma_rp_new[3]) );
  HS65_LS_AO222X4 U413 ( .A(n617), .B(n314), .C(\proc_in[MDATA][20] ), .D(n149), .E(dma_rp_new[4]), .F(n328), .Z(dma_wdata[36]) );
  HS65_LSS_XOR2X6 U414 ( .A(n53), .B(n617), .Z(dma_rp_new[4]) );
  HS65_LS_AO222X4 U415 ( .A(n618), .B(n323), .C(\proc_in[MDATA][21] ), .D(n149), .E(dma_rp_new[5]), .F(n328), .Z(dma_wdata[37]) );
  HS65_LSS_XOR2X6 U416 ( .A(n54), .B(n618), .Z(dma_rp_new[5]) );
  HS65_LS_AO222X4 U417 ( .A(n619), .B(n323), .C(\proc_in[MDATA][22] ), .D(n149), .E(dma_rp_new[6]), .F(n328), .Z(dma_wdata[38]) );
  HS65_LSS_XOR2X6 U418 ( .A(n55), .B(n619), .Z(dma_rp_new[6]) );
  HS65_LS_AO222X4 U419 ( .A(n620), .B(n323), .C(\proc_in[MDATA][23] ), .D(n149), .E(dma_rp_new[7]), .F(n328), .Z(dma_wdata[39]) );
  HS65_LSS_XOR2X6 U420 ( .A(n73), .B(n620), .Z(dma_rp_new[7]) );
  HS65_LS_AO222X4 U421 ( .A(\add_545/A[8] ), .B(n323), .C(\proc_in[MDATA][24] ), .D(n149), .E(dma_rp_new[8]), .F(n328), .Z(dma_wdata[40]) );
  HS65_LSS_XOR2X6 U422 ( .A(n52), .B(\add_545/A[8] ), .Z(dma_rp_new[8]) );
  HS65_LS_AO222X4 U423 ( .A(\add_545/A[9] ), .B(n323), .C(\proc_in[MDATA][25] ), .D(n293), .E(dma_rp_new[9]), .F(n329), .Z(dma_wdata[41]) );
  HS65_LSS_XOR2X6 U424 ( .A(n56), .B(\add_545/A[9] ), .Z(dma_rp_new[9]) );
  HS65_LS_AO222X4 U425 ( .A(\add_545/A[10] ), .B(n323), .C(
        \proc_in[MDATA][26] ), .D(n293), .E(dma_rp_new[10]), .F(n329), .Z(
        dma_wdata[42]) );
  HS65_LSS_XOR2X6 U426 ( .A(n57), .B(\add_545/A[10] ), .Z(dma_rp_new[10]) );
  HS65_LS_AO222X4 U427 ( .A(\add_545/A[11] ), .B(n323), .C(
        \proc_in[MDATA][27] ), .D(n293), .E(dma_rp_new[11]), .F(n329), .Z(
        dma_wdata[43]) );
  HS65_LSS_XOR2X6 U428 ( .A(n58), .B(\add_545/A[11] ), .Z(dma_rp_new[11]) );
  HS65_LS_AO222X4 U429 ( .A(\add_545/A[12] ), .B(n323), .C(
        \proc_in[MDATA][28] ), .D(n293), .E(dma_rp_new[12]), .F(n329), .Z(
        dma_wdata[44]) );
  HS65_LSS_XOR2X6 U430 ( .A(n59), .B(\add_545/A[12] ), .Z(dma_rp_new[12]) );
  HS65_LS_AO222X4 U431 ( .A(\add_545/A[13] ), .B(n323), .C(
        \proc_in[MDATA][29] ), .D(n293), .E(dma_rp_new[13]), .F(n329), .Z(
        dma_wdata[45]) );
  HS65_LSS_XOR2X6 U432 ( .A(n62), .B(\add_545/A[13] ), .Z(dma_rp_new[13]) );
  HS65_LS_AO222X4 U433 ( .A(\add_545/A[14] ), .B(n314), .C(
        \proc_in[MDATA][30] ), .D(n293), .E(dma_rp_new[14]), .F(n329), .Z(
        dma_wdata[46]) );
  HS65_LSS_XOR2X6 U434 ( .A(n64), .B(\add_545/A[14] ), .Z(dma_rp_new[14]) );
  HS65_LS_AO222X4 U435 ( .A(dma_rp_new[0]), .B(n323), .C(\proc_in[MDATA][16] ), 
        .D(n149), .E(dma_rp_new[0]), .F(n328), .Z(dma_wdata[32]) );
  HS65_LS_NOR2AX3 U436 ( .A(dma_rdata[32]), .B(n852), .Z(dma_rp_new[0]) );
  HS65_LS_AO222X4 U437 ( .A(\add_545/A[15] ), .B(n323), .C(
        \proc_in[MDATA][31] ), .D(n293), .E(dma_rp_new[15]), .F(n329), .Z(
        dma_wdata[47]) );
  HS65_LSS_XOR2X6 U438 ( .A(\add_545/A[15] ), .B(n3), .Z(dma_rp_new[15]) );
  HS65_LS_IVX9 U439 ( .A(n876), .Z(\add_545/A[15] ) );
  HS65_LS_OAI212X5 U440 ( .A(n118), .B(n539), .C(n23), .D(n538), .E(n537), .Z(
        pkt_out[23]) );
  HS65_LS_OAI212X5 U441 ( .A(n30), .B(n542), .C(n22), .D(n541), .E(n540), .Z(
        pkt_out[24]) );
  HS65_LH_OAI12X2 U442 ( .A(state_cnt[1]), .B(n685), .C(n313), .Z(
        phit_togo[34]) );
  HS65_LS_NAND2X7 U443 ( .A(dma_rdata[51]), .B(n138), .Z(n838) );
  HS65_LS_NAND2X7 U444 ( .A(dma_rdata[52]), .B(n138), .Z(n839) );
  HS65_LS_NAND2X7 U445 ( .A(dma_rdata[55]), .B(n138), .Z(n840) );
  HS65_LS_NAND2X7 U446 ( .A(dma_rdata[56]), .B(n138), .Z(n841) );
  HS65_LS_NAND2X7 U447 ( .A(dma_rdata[58]), .B(n138), .Z(n842) );
  HS65_LS_NAND2X7 U448 ( .A(dma_rdata[60]), .B(n138), .Z(n843) );
  HS65_LS_NAND2X7 U449 ( .A(dma_rdata[49]), .B(n139), .Z(n863) );
  HS65_LS_NAND2X7 U450 ( .A(dma_rdata[50]), .B(n139), .Z(n862) );
  HS65_LS_NAND2X7 U451 ( .A(dma_rdata[53]), .B(n139), .Z(n861) );
  HS65_LS_NAND2X7 U452 ( .A(dma_rdata[54]), .B(n139), .Z(n860) );
  HS65_LS_NAND2X7 U453 ( .A(dma_rdata[57]), .B(n139), .Z(n859) );
  HS65_LS_NAND2X7 U454 ( .A(dma_rdata[59]), .B(n139), .Z(n858) );
  HS65_LS_IVX9 U455 ( .A(dma_rdata[62]), .Z(n645) );
  HS65_LH_MUX21X4 U456 ( .D0(n122), .D1(\phase_next[1] ), .S0(n648), .Z(n682)
         );
  HS65_LS_NAND3AX6 U457 ( .A(phitIn[33]), .B(phitIn[32]), .C(phitIn[34]), .Z(
        n866) );
  HS65_LS_NAND2X7 U458 ( .A(phitIn[33]), .B(phitIn[34]), .Z(n864) );
  HS65_LS_NAND3X5 U459 ( .A(n446), .B(n577), .C(n302), .Z(n359) );
  HS65_LS_NAND2X7 U460 ( .A(dma_rdata[48]), .B(n138), .Z(n837) );
  HS65_LS_NAND2X7 U461 ( .A(dma_rdata[61]), .B(n138), .Z(n844) );
  HS65_LS_BFX9 U462 ( .A(n865), .Z(n294) );
  HS65_LS_NOR3AX2 U463 ( .A(phitIn[34]), .B(phitIn[32]), .C(phitIn[33]), .Z(
        n865) );
  HS65_LS_AO22X9 U464 ( .A(n864), .B(address[0]), .C(phitIn[17]), .D(n649), 
        .Z(n739) );
  HS65_LS_AO22X9 U465 ( .A(n864), .B(address[1]), .C(phitIn[18]), .D(n649), 
        .Z(n737) );
  HS65_LS_AO22X9 U466 ( .A(n864), .B(address[2]), .C(phitIn[19]), .D(n649), 
        .Z(n735) );
  HS65_LS_AO22X9 U467 ( .A(n864), .B(address[3]), .C(phitIn[20]), .D(n649), 
        .Z(n733) );
  HS65_LS_AO22X9 U468 ( .A(n864), .B(address[4]), .C(phitIn[21]), .D(n649), 
        .Z(n731) );
  HS65_LS_AO22X9 U469 ( .A(n864), .B(address[5]), .C(phitIn[22]), .D(n649), 
        .Z(n729) );
  HS65_LS_AO22X9 U470 ( .A(n864), .B(address[6]), .C(phitIn[23]), .D(n649), 
        .Z(n727) );
  HS65_LS_IVX9 U471 ( .A(slt_entry[3]), .Z(n646) );
  HS65_LS_IVX9 U472 ( .A(slt_entry[2]), .Z(n647) );
  HS65_LS_AO22X9 U473 ( .A(phitIn[0]), .B(n305), .C(\spm_out[MDATA][0] ), .D(
        n302), .Z(n828) );
  HS65_LS_AO22X9 U474 ( .A(phitIn[1]), .B(n311), .C(\spm_out[MDATA][1] ), .D(
        n302), .Z(n827) );
  HS65_LS_AO22X9 U475 ( .A(phitIn[2]), .B(n311), .C(\spm_out[MDATA][2] ), .D(
        n302), .Z(n826) );
  HS65_LS_AO22X9 U476 ( .A(phitIn[3]), .B(n311), .C(\spm_out[MDATA][3] ), .D(
        n302), .Z(n825) );
  HS65_LS_AO22X9 U477 ( .A(phitIn[4]), .B(n311), .C(\spm_out[MDATA][4] ), .D(
        n301), .Z(n824) );
  HS65_LS_AO22X9 U478 ( .A(phitIn[5]), .B(n311), .C(\spm_out[MDATA][5] ), .D(
        n866), .Z(n823) );
  HS65_LS_AO22X9 U479 ( .A(phitIn[6]), .B(n311), .C(\spm_out[MDATA][6] ), .D(
        n300), .Z(n822) );
  HS65_LS_AO22X9 U480 ( .A(phitIn[7]), .B(n311), .C(\spm_out[MDATA][7] ), .D(
        n866), .Z(n821) );
  HS65_LS_AO22X9 U481 ( .A(phitIn[8]), .B(n311), .C(\spm_out[MDATA][8] ), .D(
        n866), .Z(n820) );
  HS65_LS_AO22X9 U482 ( .A(phitIn[9]), .B(n311), .C(\spm_out[MDATA][9] ), .D(
        n866), .Z(n819) );
  HS65_LS_AO22X9 U483 ( .A(phitIn[10]), .B(n310), .C(\spm_out[MDATA][10] ), 
        .D(n866), .Z(n818) );
  HS65_LS_AO22X9 U484 ( .A(phitIn[11]), .B(n310), .C(\spm_out[MDATA][11] ), 
        .D(n866), .Z(n817) );
  HS65_LS_AO22X9 U485 ( .A(phitIn[12]), .B(n310), .C(\spm_out[MDATA][12] ), 
        .D(n866), .Z(n816) );
  HS65_LS_AO22X9 U486 ( .A(phitIn[13]), .B(n310), .C(\spm_out[MDATA][13] ), 
        .D(n866), .Z(n815) );
  HS65_LS_AO22X9 U487 ( .A(phitIn[14]), .B(n310), .C(\spm_out[MDATA][14] ), 
        .D(n866), .Z(n814) );
  HS65_LS_AO22X9 U488 ( .A(phitIn[15]), .B(n310), .C(\spm_out[MDATA][15] ), 
        .D(n866), .Z(n813) );
  HS65_LS_AO22X9 U489 ( .A(phitIn[16]), .B(n310), .C(\spm_out[MDATA][16] ), 
        .D(n866), .Z(n812) );
  HS65_LS_AO22X9 U490 ( .A(phitIn[17]), .B(n310), .C(\spm_out[MDATA][17] ), 
        .D(n866), .Z(n811) );
  HS65_LS_AO22X9 U491 ( .A(phitIn[18]), .B(n310), .C(\spm_out[MDATA][18] ), 
        .D(n866), .Z(n810) );
  HS65_LS_AO22X9 U492 ( .A(phitIn[19]), .B(n310), .C(\spm_out[MDATA][19] ), 
        .D(n302), .Z(n809) );
  HS65_LS_AO22X9 U493 ( .A(phitIn[20]), .B(n310), .C(\spm_out[MDATA][20] ), 
        .D(n302), .Z(n808) );
  HS65_LS_AO22X9 U494 ( .A(phitIn[21]), .B(n310), .C(\spm_out[MDATA][21] ), 
        .D(n302), .Z(n807) );
  HS65_LS_AO22X9 U495 ( .A(phitIn[22]), .B(n310), .C(\spm_out[MDATA][22] ), 
        .D(n302), .Z(n806) );
  HS65_LS_AO22X9 U496 ( .A(phitIn[23]), .B(n310), .C(\spm_out[MDATA][23] ), 
        .D(n302), .Z(n805) );
  HS65_LS_AO22X9 U497 ( .A(phitIn[24]), .B(n310), .C(\spm_out[MDATA][24] ), 
        .D(n302), .Z(n804) );
  HS65_LS_AO22X9 U498 ( .A(phitIn[25]), .B(n310), .C(\spm_out[MDATA][25] ), 
        .D(n302), .Z(n803) );
  HS65_LS_AO22X9 U499 ( .A(phitIn[26]), .B(n310), .C(\spm_out[MDATA][26] ), 
        .D(n302), .Z(n802) );
  HS65_LS_AO22X9 U500 ( .A(phitIn[27]), .B(n310), .C(\spm_out[MDATA][27] ), 
        .D(n302), .Z(n801) );
  HS65_LS_AO22X9 U501 ( .A(phitIn[28]), .B(n310), .C(\spm_out[MDATA][28] ), 
        .D(n302), .Z(n800) );
  HS65_LS_AO22X9 U502 ( .A(phitIn[29]), .B(n310), .C(\spm_out[MDATA][29] ), 
        .D(n302), .Z(n799) );
  HS65_LS_AO22X9 U503 ( .A(phitIn[30]), .B(n306), .C(\spm_out[MDATA][30] ), 
        .D(n302), .Z(n798) );
  HS65_LS_AO22X9 U504 ( .A(phitIn[31]), .B(n306), .C(\spm_out[MDATA][31] ), 
        .D(n302), .Z(n797) );
  HS65_LS_AO22X9 U505 ( .A(dIn_h[0]), .B(n306), .C(\spm_out[MDATA][32] ), .D(
        n301), .Z(n796) );
  HS65_LS_AO22X9 U506 ( .A(dIn_h[1]), .B(n306), .C(\spm_out[MDATA][33] ), .D(
        n301), .Z(n795) );
  HS65_LS_AO22X9 U507 ( .A(dIn_h[2]), .B(n306), .C(\spm_out[MDATA][34] ), .D(
        n301), .Z(n794) );
  HS65_LS_AO22X9 U508 ( .A(dIn_h[3]), .B(n306), .C(\spm_out[MDATA][35] ), .D(
        n301), .Z(n793) );
  HS65_LS_AO22X9 U509 ( .A(dIn_h[4]), .B(n306), .C(\spm_out[MDATA][36] ), .D(
        n301), .Z(n792) );
  HS65_LS_AO22X9 U510 ( .A(dIn_h[5]), .B(n306), .C(\spm_out[MDATA][37] ), .D(
        n301), .Z(n791) );
  HS65_LS_AO22X9 U511 ( .A(dIn_h[6]), .B(n306), .C(\spm_out[MDATA][38] ), .D(
        n301), .Z(n790) );
  HS65_LS_AO22X9 U512 ( .A(dIn_h[7]), .B(n306), .C(\spm_out[MDATA][39] ), .D(
        n301), .Z(n789) );
  HS65_LS_AO22X9 U513 ( .A(dIn_h[8]), .B(n306), .C(\spm_out[MDATA][40] ), .D(
        n301), .Z(n788) );
  HS65_LS_AO22X9 U514 ( .A(dIn_h[9]), .B(n306), .C(\spm_out[MDATA][41] ), .D(
        n301), .Z(n787) );
  HS65_LS_AO22X9 U515 ( .A(dIn_h[10]), .B(n306), .C(\spm_out[MDATA][42] ), .D(
        n301), .Z(n786) );
  HS65_LS_AO22X9 U516 ( .A(dIn_h[11]), .B(n306), .C(\spm_out[MDATA][43] ), .D(
        n301), .Z(n785) );
  HS65_LS_AO22X9 U517 ( .A(dIn_h[12]), .B(n306), .C(\spm_out[MDATA][44] ), .D(
        n300), .Z(n784) );
  HS65_LS_AO22X9 U518 ( .A(dIn_h[13]), .B(n306), .C(\spm_out[MDATA][45] ), .D(
        n300), .Z(n783) );
  HS65_LS_AO22X9 U519 ( .A(dIn_h[14]), .B(n306), .C(\spm_out[MDATA][46] ), .D(
        n300), .Z(n782) );
  HS65_LS_AO22X9 U520 ( .A(dIn_h[15]), .B(n306), .C(\spm_out[MDATA][47] ), .D(
        n300), .Z(n781) );
  HS65_LS_AO22X9 U521 ( .A(dIn_h[16]), .B(n306), .C(\spm_out[MDATA][48] ), .D(
        n300), .Z(n780) );
  HS65_LS_AO22X9 U522 ( .A(dIn_h[17]), .B(n305), .C(\spm_out[MDATA][49] ), .D(
        n300), .Z(n779) );
  HS65_LS_AO22X9 U523 ( .A(dIn_h[18]), .B(n305), .C(\spm_out[MDATA][50] ), .D(
        n300), .Z(n778) );
  HS65_LS_AO22X9 U524 ( .A(dIn_h[19]), .B(n305), .C(\spm_out[MDATA][51] ), .D(
        n300), .Z(n777) );
  HS65_LS_AO22X9 U525 ( .A(dIn_h[20]), .B(n306), .C(\spm_out[MDATA][52] ), .D(
        n300), .Z(n776) );
  HS65_LS_AO22X9 U526 ( .A(dIn_h[21]), .B(n305), .C(\spm_out[MDATA][53] ), .D(
        n301), .Z(n775) );
  HS65_LS_AO22X9 U527 ( .A(dIn_h[22]), .B(n305), .C(\spm_out[MDATA][54] ), .D(
        n300), .Z(n774) );
  HS65_LS_AO22X9 U528 ( .A(dIn_h[23]), .B(n305), .C(\spm_out[MDATA][55] ), .D(
        n300), .Z(n773) );
  HS65_LS_AO22X9 U529 ( .A(dIn_h[24]), .B(n305), .C(\spm_out[MDATA][56] ), .D(
        n300), .Z(n772) );
  HS65_LS_AO22X9 U530 ( .A(dIn_h[25]), .B(n305), .C(\spm_out[MDATA][57] ), .D(
        n300), .Z(n771) );
  HS65_LS_AO22X9 U531 ( .A(dIn_h[26]), .B(n305), .C(\spm_out[MDATA][58] ), .D(
        n300), .Z(n770) );
  HS65_LS_AO22X9 U532 ( .A(dIn_h[27]), .B(n305), .C(\spm_out[MDATA][59] ), .D(
        n301), .Z(n769) );
  HS65_LS_AO22X9 U533 ( .A(dIn_h[28]), .B(n305), .C(\spm_out[MDATA][60] ), .D(
        n300), .Z(n768) );
  HS65_LS_AO22X9 U534 ( .A(dIn_h[29]), .B(n305), .C(\spm_out[MDATA][61] ), .D(
        n301), .Z(n767) );
  HS65_LS_AO22X9 U535 ( .A(dIn_h[30]), .B(n305), .C(\spm_out[MDATA][62] ), .D(
        n300), .Z(n766) );
  HS65_LS_AO22X9 U536 ( .A(dIn_h[31]), .B(n305), .C(\spm_out[MDATA][63] ), .D(
        n302), .Z(n765) );
  HS65_LS_AO22X9 U537 ( .A(phitIn[17]), .B(n298), .C(n296), .D(dIn_h[17]), .Z(
        n740) );
  HS65_LS_AO22X9 U538 ( .A(phitIn[18]), .B(n298), .C(n296), .D(dIn_h[18]), .Z(
        n738) );
  HS65_LS_AO22X9 U539 ( .A(phitIn[19]), .B(n298), .C(n296), .D(dIn_h[19]), .Z(
        n736) );
  HS65_LS_AO22X9 U540 ( .A(phitIn[20]), .B(n298), .C(n296), .D(dIn_h[20]), .Z(
        n734) );
  HS65_LS_AO22X9 U541 ( .A(phitIn[21]), .B(n299), .C(n296), .D(dIn_h[21]), .Z(
        n732) );
  HS65_LS_AO22X9 U542 ( .A(phitIn[22]), .B(n299), .C(n296), .D(dIn_h[22]), .Z(
        n730) );
  HS65_LS_AO22X9 U543 ( .A(phitIn[23]), .B(n299), .C(n296), .D(dIn_h[23]), .Z(
        n728) );
  HS65_LS_AO22X9 U544 ( .A(phitIn[0]), .B(n297), .C(n295), .D(dIn_h[0]), .Z(
        n757) );
  HS65_LS_AO22X9 U545 ( .A(phitIn[1]), .B(n298), .C(n295), .D(dIn_h[1]), .Z(
        n756) );
  HS65_LS_AO22X9 U546 ( .A(phitIn[2]), .B(n298), .C(n295), .D(dIn_h[2]), .Z(
        n755) );
  HS65_LS_AO22X9 U547 ( .A(phitIn[3]), .B(n298), .C(n295), .D(dIn_h[3]), .Z(
        n754) );
  HS65_LS_AO22X9 U548 ( .A(phitIn[4]), .B(n298), .C(n295), .D(dIn_h[4]), .Z(
        n753) );
  HS65_LS_AO22X9 U549 ( .A(phitIn[5]), .B(n298), .C(n295), .D(dIn_h[5]), .Z(
        n752) );
  HS65_LS_AO22X9 U550 ( .A(phitIn[6]), .B(n298), .C(n295), .D(dIn_h[6]), .Z(
        n751) );
  HS65_LS_AO22X9 U551 ( .A(phitIn[7]), .B(n298), .C(n295), .D(dIn_h[7]), .Z(
        n750) );
  HS65_LS_AO22X9 U552 ( .A(phitIn[8]), .B(n298), .C(n295), .D(dIn_h[8]), .Z(
        n749) );
  HS65_LS_AO22X9 U553 ( .A(phitIn[9]), .B(n298), .C(n295), .D(dIn_h[9]), .Z(
        n748) );
  HS65_LS_AO22X9 U554 ( .A(phitIn[10]), .B(n298), .C(n295), .D(dIn_h[10]), .Z(
        n747) );
  HS65_LS_AO22X9 U555 ( .A(phitIn[11]), .B(n298), .C(n295), .D(dIn_h[11]), .Z(
        n746) );
  HS65_LS_AO22X9 U556 ( .A(phitIn[12]), .B(n298), .C(n295), .D(dIn_h[12]), .Z(
        n745) );
  HS65_LS_AO22X9 U557 ( .A(phitIn[13]), .B(n298), .C(n296), .D(dIn_h[13]), .Z(
        n744) );
  HS65_LS_AO22X9 U558 ( .A(phitIn[14]), .B(n298), .C(n296), .D(dIn_h[14]), .Z(
        n743) );
  HS65_LS_AO22X9 U559 ( .A(phitIn[15]), .B(n298), .C(n296), .D(dIn_h[15]), .Z(
        n742) );
  HS65_LS_AO22X9 U560 ( .A(phitIn[16]), .B(n298), .C(n296), .D(dIn_h[16]), .Z(
        n741) );
  HS65_LS_AO22X9 U561 ( .A(phitIn[24]), .B(n299), .C(n296), .D(dIn_h[24]), .Z(
        n726) );
  HS65_LS_AO22X9 U562 ( .A(phitIn[25]), .B(n299), .C(n296), .D(dIn_h[25]), .Z(
        n725) );
  HS65_LS_AO22X9 U563 ( .A(phitIn[26]), .B(n299), .C(n295), .D(dIn_h[26]), .Z(
        n724) );
  HS65_LS_AO22X9 U564 ( .A(phitIn[27]), .B(n299), .C(n296), .D(dIn_h[27]), .Z(
        n723) );
  HS65_LS_AO22X9 U565 ( .A(phitIn[28]), .B(n299), .C(n295), .D(dIn_h[28]), .Z(
        n722) );
  HS65_LS_AO22X9 U566 ( .A(phitIn[29]), .B(n299), .C(n296), .D(dIn_h[29]), .Z(
        n721) );
  HS65_LS_AO22X9 U567 ( .A(phitIn[30]), .B(n299), .C(n295), .D(dIn_h[30]), .Z(
        n720) );
  HS65_LS_AO22X9 U568 ( .A(phitIn[31]), .B(n299), .C(n296), .D(dIn_h[31]), .Z(
        n719) );
  HS65_LS_AO22X9 U569 ( .A(n305), .B(address[0]), .C(n301), .D(flit_buf[64]), 
        .Z(n764) );
  HS65_LS_AO22X9 U570 ( .A(n305), .B(address[1]), .C(n300), .D(flit_buf[65]), 
        .Z(n763) );
  HS65_LS_AO22X9 U571 ( .A(n305), .B(address[2]), .C(n301), .D(flit_buf[66]), 
        .Z(n762) );
  HS65_LS_AO22X9 U572 ( .A(n305), .B(address[3]), .C(n300), .D(flit_buf[67]), 
        .Z(n761) );
  HS65_LS_AO22X9 U573 ( .A(n304), .B(address[4]), .C(n301), .D(flit_buf[68]), 
        .Z(n760) );
  HS65_LS_AO22X9 U574 ( .A(n303), .B(address[5]), .C(n300), .D(flit_buf[69]), 
        .Z(n759) );
  HS65_LS_AO22X9 U575 ( .A(n305), .B(address[6]), .C(n301), .D(flit_buf[70]), 
        .Z(n758) );
  HS65_LS_OR2X9 U576 ( .A(vld_pkt), .B(n649), .Z(n680) );
  HS65_LS_NAND2X7 U577 ( .A(\proc_in[MADDR][0] ), .B(n832), .Z(n857) );
  HS65_LS_NOR4ABX2 U578 ( .A(n656), .B(n829), .C(\proc_in[MADDR][26] ), .D(
        \proc_in[MADDR][24] ), .Z(n856) );
  HS65_LS_IVX9 U579 ( .A(\proc_in[MADDR][25] ), .Z(n656) );
  HS65_LS_NOR3X4 U580 ( .A(\proc_in[MADDR][27] ), .B(\proc_in[MADDR][31] ), 
        .C(\proc_in[MADDR][30] ), .Z(n829) );
  HS65_LS_NAND4ABX3 U581 ( .A(\proc_in[MADDR][29] ), .B(\proc_in[MADDR][26] ), 
        .C(n831), .D(n830), .Z(n854) );
  HS65_LS_NOR2X6 U582 ( .A(\proc_in[MADDR][31] ), .B(\proc_in[MADDR][30] ), 
        .Z(n831) );
  HS65_LS_NOR4ABX2 U583 ( .A(\proc_in[MADDR][28] ), .B(\proc_in[MADDR][27] ), 
        .C(\proc_in[MADDR][25] ), .D(\proc_in[MADDR][24] ), .Z(n830) );
  HS65_LS_NOR3AX2 U584 ( .A(n856), .B(n655), .C(\proc_in[MADDR][29] ), .Z(n676) );
  HS65_LS_NAND4ABX3 U585 ( .A(config_reg[3]), .B(n870), .C(config_reg[4]), .D(
        n593), .Z(n871) );
  HS65_LS_OA32X4 U586 ( .A(config_reg[0]), .B(config_reg[1]), .C(n650), .D(
        n869), .E(config_reg[2]), .Z(n870) );
  HS65_LS_IVX9 U587 ( .A(config_reg[2]), .Z(n650) );
  HS65_LSS_XNOR2X6 U588 ( .A(config_reg[1]), .B(config_reg[0]), .Z(n869) );
  HS65_LS_BFX9 U589 ( .A(na_reset), .Z(n336) );
  HS65_LS_BFX9 U590 ( .A(na_reset), .Z(n335) );
  HS65_LS_NAND2X7 U591 ( .A(n676), .B(\proc_in[MCMD][0] ), .Z(n868) );
  HS65_LS_IVX9 U592 ( .A(\proc_in[MDATA][15] ), .Z(n660) );
  HS65_LS_IVX9 U593 ( .A(\proc_in[MDATA][6] ), .Z(n669) );
  HS65_LS_IVX9 U594 ( .A(\proc_in[MDATA][7] ), .Z(n668) );
  HS65_LS_IVX9 U595 ( .A(\proc_in[MDATA][8] ), .Z(n667) );
  HS65_LS_IVX9 U596 ( .A(\proc_in[MDATA][9] ), .Z(n666) );
  HS65_LS_IVX9 U597 ( .A(\proc_in[MADDR][28] ), .Z(n655) );
  HS65_LS_AND3X9 U598 ( .A(n856), .B(n655), .C(\proc_in[MADDR][29] ), .Z(n832)
         );
  HS65_LS_IVX9 U599 ( .A(\proc_in[MDATA][14] ), .Z(n661) );
  HS65_LS_IVX9 U600 ( .A(\proc_in[MDATA][0] ), .Z(n675) );
  HS65_LS_IVX9 U601 ( .A(\proc_in[MDATA][1] ), .Z(n674) );
  HS65_LS_IVX9 U602 ( .A(\proc_in[MDATA][2] ), .Z(n673) );
  HS65_LS_IVX9 U603 ( .A(\proc_in[MDATA][3] ), .Z(n672) );
  HS65_LS_IVX9 U604 ( .A(\proc_in[MDATA][4] ), .Z(n671) );
  HS65_LS_IVX9 U605 ( .A(\proc_in[MDATA][5] ), .Z(n670) );
  HS65_LS_IVX9 U606 ( .A(\proc_in[MDATA][10] ), .Z(n665) );
  HS65_LS_IVX9 U607 ( .A(\proc_in[MDATA][11] ), .Z(n664) );
  HS65_LS_IVX9 U608 ( .A(\proc_in[MDATA][12] ), .Z(n663) );
  HS65_LS_IVX9 U609 ( .A(\proc_in[MDATA][13] ), .Z(n662) );
  HS65_LS_IVX9 U610 ( .A(\proc_in[MADDR][0] ), .Z(n659) );
  HS65_LS_IVX9 U611 ( .A(\proc_in[MADDR][1] ), .Z(n658) );
  HS65_LH_NAND2X2 U612 ( .A(n26), .B(n20), .Z(n362) );
  HS65_LH_AND2X4 U613 ( .A(n26), .B(n412), .Z(phit_togo[32]) );
  HS65_LH_BFX2 U614 ( .A(n120), .Z(n133) );
  HS65_LS_BFX9 U615 ( .A(n133), .Z(n136) );
  HS65_LS_BFX9 U616 ( .A(n133), .Z(n134) );
  HS65_LS_BFX9 U617 ( .A(n133), .Z(n137) );
  HS65_LS_NAND2X5 U618 ( .A(n445), .B(n20), .Z(n361) );
  HS65_LH_NAND2X2 U619 ( .A(n445), .B(n20), .Z(n446) );
  HS65_LH_CBI4I1X5 U620 ( .A(n446), .B(n360), .C(n302), .D(n359), .Z(n681) );
  HS65_LS_IVX18 U621 ( .A(\phase_prev[0] ), .Z(n451) );
  HS65_LS_IVX9 U622 ( .A(n37), .Z(n648) );
  HS65_LS_IVX9 U623 ( .A(n852), .Z(n621) );
  HS65_LS_NAND2X7 U624 ( .A(dma_rdata[39]), .B(n139), .Z(n591) );
  HS65_LS_IVX9 U625 ( .A(n591), .Z(n620) );
  HS65_LS_NAND2X7 U626 ( .A(dma_rdata[38]), .B(n139), .Z(n589) );
  HS65_LS_IVX9 U627 ( .A(n589), .Z(n619) );
  HS65_LS_NAND2X7 U628 ( .A(dma_rdata[37]), .B(n140), .Z(n587) );
  HS65_LS_IVX9 U629 ( .A(n587), .Z(n618) );
  HS65_LS_NAND2X7 U630 ( .A(dma_rdata[36]), .B(n140), .Z(n585) );
  HS65_LS_IVX9 U631 ( .A(n585), .Z(n617) );
  HS65_LS_NAND2X7 U632 ( .A(dma_rdata[35]), .B(n140), .Z(n583) );
  HS65_LS_IVX9 U633 ( .A(n583), .Z(n616) );
  HS65_LS_NAND2X7 U634 ( .A(dma_rdata[34]), .B(n140), .Z(n581) );
  HS65_LS_IVX9 U635 ( .A(n581), .Z(n615) );
  HS65_LS_NAND2X7 U636 ( .A(dma_rdata[33]), .B(n140), .Z(n579) );
  HS65_LS_IVX9 U637 ( .A(n579), .Z(n614) );
  HS65_LS_NAND2X7 U638 ( .A(dma_rdata[31]), .B(n140), .Z(n410) );
  HS65_LS_IVX9 U639 ( .A(n410), .Z(n613) );
  HS65_LS_NAND2X7 U640 ( .A(dma_rdata[30]), .B(n140), .Z(n408) );
  HS65_LS_IVX9 U641 ( .A(n408), .Z(n612) );
  HS65_LS_NAND2X7 U642 ( .A(dma_rdata[29]), .B(n140), .Z(n406) );
  HS65_LS_IVX9 U643 ( .A(n406), .Z(n611) );
  HS65_LS_NAND2X7 U644 ( .A(dma_rdata[28]), .B(n140), .Z(n404) );
  HS65_LS_IVX9 U645 ( .A(n404), .Z(n610) );
  HS65_LS_NAND2X7 U646 ( .A(dma_rdata[27]), .B(n140), .Z(n402) );
  HS65_LS_IVX9 U647 ( .A(n402), .Z(n609) );
  HS65_LS_NAND2X7 U648 ( .A(dma_rdata[26]), .B(n140), .Z(n400) );
  HS65_LS_IVX9 U649 ( .A(n400), .Z(n608) );
  HS65_LS_NAND2X7 U650 ( .A(dma_rdata[25]), .B(n140), .Z(n398) );
  HS65_LS_IVX9 U651 ( .A(n398), .Z(n607) );
  HS65_LS_NAND2X7 U652 ( .A(dma_rdata[24]), .B(n140), .Z(n396) );
  HS65_LS_IVX9 U653 ( .A(n396), .Z(n606) );
  HS65_LS_NAND2X7 U654 ( .A(dma_rdata[23]), .B(n140), .Z(n394) );
  HS65_LS_IVX9 U655 ( .A(n394), .Z(n605) );
  HS65_LS_NAND2X7 U656 ( .A(dma_rdata[22]), .B(n140), .Z(n392) );
  HS65_LS_IVX9 U657 ( .A(n392), .Z(n604) );
  HS65_LS_NAND2X7 U658 ( .A(dma_rdata[21]), .B(n140), .Z(n390) );
  HS65_LS_IVX9 U659 ( .A(n390), .Z(n603) );
  HS65_LS_NAND2X7 U660 ( .A(dma_rdata[20]), .B(n140), .Z(n388) );
  HS65_LS_IVX9 U661 ( .A(n388), .Z(n602) );
  HS65_LS_NAND2X7 U662 ( .A(dma_rdata[19]), .B(n139), .Z(n386) );
  HS65_LS_IVX9 U663 ( .A(n386), .Z(n601) );
  HS65_LS_NAND2X7 U664 ( .A(dma_rdata[18]), .B(n139), .Z(n384) );
  HS65_LS_IVX9 U665 ( .A(n384), .Z(n600) );
  HS65_LS_NAND2X7 U666 ( .A(dma_rdata[17]), .B(n139), .Z(n382) );
  HS65_LS_IVX9 U667 ( .A(n382), .Z(n599) );
  HS65_LS_IVX9 U668 ( .A(\proc_in[MCMD][0] ), .Z(n356) );
  HS65_LS_IVX9 U669 ( .A(n358), .Z(n357) );
  HS65_LS_NAND2X7 U670 ( .A(n835), .B(n1), .Z(n853) );
  HS65_LS_OAI22X6 U671 ( .A(n646), .B(n362), .C(n834), .D(n358), .Z(
        dma_raddr[1]) );
  HS65_LS_OAI22X6 U672 ( .A(n647), .B(n362), .C(n833), .D(n358), .Z(
        dma_raddr[0]) );
  HS65_LS_NAND2X7 U673 ( .A(dma_rdata[16]), .B(n139), .Z(n380) );
  HS65_LS_IVX9 U674 ( .A(n380), .Z(n596) );
  HS65_LS_IVX9 U675 ( .A(n686), .Z(n452) );
  HS65_LS_IVX9 U676 ( .A(vld_pkt), .Z(n360) );
  HS65_LS_IVX9 U677 ( .A(n684), .Z(n577) );
  HS65_LS_IVX9 U678 ( .A(n362), .Z(n598) );
  HS65_LS_IVX9 U679 ( .A(n685), .Z(n412) );
  HS65_LS_NAND2X7 U680 ( .A(n598), .B(n412), .Z(n411) );
  HS65_LS_IVX9 U681 ( .A(dOut_l[0]), .Z(n413) );
  HS65_LS_NAND2X7 U682 ( .A(\spm_in[SDATA][32] ), .B(n124), .Z(n363) );
  HS65_LS_OAI212X5 U683 ( .A(n129), .B(n413), .C(n325), .D(n643), .E(n363), 
        .Z(mux_out[0]) );
  HS65_LS_IVX9 U684 ( .A(dOut_l[1]), .Z(n414) );
  HS65_LS_NAND2X7 U685 ( .A(\spm_in[SDATA][33] ), .B(n124), .Z(n364) );
  HS65_LS_OAI212X5 U686 ( .A(n129), .B(n414), .C(n325), .D(n642), .E(n364), 
        .Z(mux_out[1]) );
  HS65_LS_IVX9 U687 ( .A(dOut_l[2]), .Z(n415) );
  HS65_LS_NAND2X7 U688 ( .A(\spm_in[SDATA][34] ), .B(n124), .Z(n365) );
  HS65_LS_OAI212X5 U689 ( .A(n129), .B(n415), .C(n325), .D(n641), .E(n365), 
        .Z(mux_out[2]) );
  HS65_LS_IVX9 U690 ( .A(dOut_l[3]), .Z(n416) );
  HS65_LS_NAND2X7 U691 ( .A(\spm_in[SDATA][35] ), .B(n124), .Z(n366) );
  HS65_LS_OAI212X5 U692 ( .A(n129), .B(n416), .C(n325), .D(n640), .E(n366), 
        .Z(mux_out[3]) );
  HS65_LS_IVX9 U693 ( .A(dOut_l[4]), .Z(n417) );
  HS65_LS_NAND2X7 U694 ( .A(\spm_in[SDATA][36] ), .B(n124), .Z(n367) );
  HS65_LS_OAI212X5 U695 ( .A(n129), .B(n417), .C(n325), .D(n639), .E(n367), 
        .Z(mux_out[4]) );
  HS65_LS_IVX9 U696 ( .A(dOut_l[5]), .Z(n418) );
  HS65_LS_NAND2X7 U697 ( .A(\spm_in[SDATA][37] ), .B(n124), .Z(n368) );
  HS65_LS_OAI212X5 U698 ( .A(n129), .B(n418), .C(n325), .D(n638), .E(n368), 
        .Z(mux_out[5]) );
  HS65_LS_IVX9 U699 ( .A(dOut_l[6]), .Z(n419) );
  HS65_LS_NAND2X7 U700 ( .A(\spm_in[SDATA][38] ), .B(n124), .Z(n369) );
  HS65_LS_OAI212X5 U701 ( .A(n129), .B(n419), .C(n325), .D(n637), .E(n369), 
        .Z(mux_out[6]) );
  HS65_LS_IVX9 U702 ( .A(dOut_l[7]), .Z(n420) );
  HS65_LS_NAND2X7 U703 ( .A(\spm_in[SDATA][39] ), .B(n124), .Z(n370) );
  HS65_LS_OAI212X5 U704 ( .A(n129), .B(n420), .C(n325), .D(n636), .E(n370), 
        .Z(mux_out[7]) );
  HS65_LS_IVX9 U705 ( .A(dOut_l[8]), .Z(n421) );
  HS65_LS_NAND2X7 U706 ( .A(\spm_in[SDATA][40] ), .B(n124), .Z(n371) );
  HS65_LS_OAI212X5 U707 ( .A(n129), .B(n421), .C(n325), .D(n635), .E(n371), 
        .Z(mux_out[8]) );
  HS65_LS_IVX9 U708 ( .A(dOut_l[9]), .Z(n422) );
  HS65_LS_NAND2X7 U709 ( .A(\spm_in[SDATA][41] ), .B(n124), .Z(n372) );
  HS65_LS_OAI212X5 U710 ( .A(n129), .B(n422), .C(n324), .D(n634), .E(n372), 
        .Z(mux_out[9]) );
  HS65_LS_IVX9 U711 ( .A(dOut_l[10]), .Z(n423) );
  HS65_LS_NAND2X7 U712 ( .A(\spm_in[SDATA][42] ), .B(n124), .Z(n373) );
  HS65_LS_OAI212X5 U713 ( .A(n129), .B(n423), .C(n324), .D(n633), .E(n373), 
        .Z(mux_out[10]) );
  HS65_LS_IVX9 U714 ( .A(dOut_l[11]), .Z(n424) );
  HS65_LS_NAND2X7 U715 ( .A(\spm_in[SDATA][43] ), .B(n124), .Z(n374) );
  HS65_LS_OAI212X5 U716 ( .A(n129), .B(n424), .C(n324), .D(n632), .E(n374), 
        .Z(mux_out[11]) );
  HS65_LS_IVX9 U717 ( .A(dOut_l[12]), .Z(n425) );
  HS65_LS_NAND2X7 U718 ( .A(\spm_in[SDATA][44] ), .B(n125), .Z(n375) );
  HS65_LS_OAI212X5 U719 ( .A(n130), .B(n425), .C(n324), .D(n631), .E(n375), 
        .Z(mux_out[12]) );
  HS65_LS_IVX9 U720 ( .A(dOut_l[13]), .Z(n426) );
  HS65_LS_NAND2X7 U721 ( .A(\spm_in[SDATA][45] ), .B(n125), .Z(n376) );
  HS65_LS_OAI212X5 U722 ( .A(n130), .B(n426), .C(n324), .D(n630), .E(n376), 
        .Z(mux_out[13]) );
  HS65_LS_IVX9 U723 ( .A(dOut_l[14]), .Z(n427) );
  HS65_LS_NAND2X7 U724 ( .A(\spm_in[SDATA][46] ), .B(n125), .Z(n377) );
  HS65_LS_OAI212X5 U725 ( .A(n130), .B(n427), .C(n324), .D(n629), .E(n377), 
        .Z(mux_out[14]) );
  HS65_LS_IVX9 U726 ( .A(dOut_l[15]), .Z(n428) );
  HS65_LS_NAND2X7 U727 ( .A(\spm_in[SDATA][47] ), .B(n125), .Z(n378) );
  HS65_LS_OAI212X5 U728 ( .A(n130), .B(n428), .C(n324), .D(n628), .E(n378), 
        .Z(mux_out[15]) );
  HS65_LS_IVX9 U729 ( .A(dOut_l[16]), .Z(n429) );
  HS65_LS_NAND2X7 U730 ( .A(\spm_in[SDATA][48] ), .B(n125), .Z(n379) );
  HS65_LS_OAI212X5 U731 ( .A(n130), .B(n429), .C(n324), .D(n380), .E(n379), 
        .Z(mux_out[16]) );
  HS65_LS_IVX9 U732 ( .A(dOut_l[17]), .Z(n430) );
  HS65_LS_NAND2X7 U733 ( .A(\spm_in[SDATA][49] ), .B(n125), .Z(n381) );
  HS65_LS_OAI212X5 U734 ( .A(n130), .B(n430), .C(n324), .D(n382), .E(n381), 
        .Z(mux_out[17]) );
  HS65_LS_IVX9 U735 ( .A(dOut_l[18]), .Z(n431) );
  HS65_LS_NAND2X7 U736 ( .A(\spm_in[SDATA][50] ), .B(n125), .Z(n383) );
  HS65_LS_OAI212X5 U737 ( .A(n130), .B(n431), .C(n324), .D(n384), .E(n383), 
        .Z(mux_out[18]) );
  HS65_LS_IVX9 U738 ( .A(dOut_l[19]), .Z(n432) );
  HS65_LS_NAND2X7 U739 ( .A(\spm_in[SDATA][51] ), .B(n125), .Z(n385) );
  HS65_LS_OAI212X5 U740 ( .A(n130), .B(n432), .C(n324), .D(n386), .E(n385), 
        .Z(mux_out[19]) );
  HS65_LS_IVX9 U741 ( .A(dOut_l[20]), .Z(n433) );
  HS65_LS_NAND2X7 U742 ( .A(\spm_in[SDATA][52] ), .B(n125), .Z(n387) );
  HS65_LS_OAI212X5 U743 ( .A(n130), .B(n433), .C(n324), .D(n388), .E(n387), 
        .Z(mux_out[20]) );
  HS65_LS_IVX9 U744 ( .A(dOut_l[21]), .Z(n434) );
  HS65_LS_NAND2X7 U745 ( .A(\spm_in[SDATA][53] ), .B(n125), .Z(n389) );
  HS65_LS_OAI212X5 U746 ( .A(n130), .B(n434), .C(n324), .D(n390), .E(n389), 
        .Z(mux_out[21]) );
  HS65_LS_IVX9 U747 ( .A(dOut_l[22]), .Z(n435) );
  HS65_LS_NAND2X7 U748 ( .A(\spm_in[SDATA][54] ), .B(n125), .Z(n391) );
  HS65_LS_OAI212X5 U749 ( .A(n130), .B(n435), .C(n324), .D(n392), .E(n391), 
        .Z(mux_out[22]) );
  HS65_LS_IVX9 U750 ( .A(dOut_l[23]), .Z(n436) );
  HS65_LS_NAND2X7 U751 ( .A(\spm_in[SDATA][55] ), .B(n125), .Z(n393) );
  HS65_LS_OAI212X5 U752 ( .A(n130), .B(n436), .C(n324), .D(n394), .E(n393), 
        .Z(mux_out[23]) );
  HS65_LS_IVX9 U753 ( .A(dOut_l[24]), .Z(n437) );
  HS65_LS_NAND2X7 U754 ( .A(\spm_in[SDATA][56] ), .B(n127), .Z(n395) );
  HS65_LS_OAI212X5 U755 ( .A(n132), .B(n437), .C(n324), .D(n396), .E(n395), 
        .Z(mux_out[24]) );
  HS65_LS_IVX9 U756 ( .A(dOut_l[25]), .Z(n438) );
  HS65_LS_NAND2X7 U757 ( .A(\spm_in[SDATA][57] ), .B(n127), .Z(n397) );
  HS65_LS_OAI212X5 U758 ( .A(n132), .B(n438), .C(n324), .D(n398), .E(n397), 
        .Z(mux_out[25]) );
  HS65_LS_IVX9 U759 ( .A(dOut_l[26]), .Z(n439) );
  HS65_LS_NAND2X7 U760 ( .A(\spm_in[SDATA][58] ), .B(n127), .Z(n399) );
  HS65_LS_OAI212X5 U761 ( .A(n132), .B(n439), .C(n324), .D(n400), .E(n399), 
        .Z(mux_out[26]) );
  HS65_LS_IVX9 U762 ( .A(dOut_l[27]), .Z(n440) );
  HS65_LS_NAND2X7 U763 ( .A(\spm_in[SDATA][59] ), .B(n127), .Z(n401) );
  HS65_LS_OAI212X5 U764 ( .A(n132), .B(n440), .C(n323), .D(n402), .E(n401), 
        .Z(mux_out[27]) );
  HS65_LS_IVX9 U765 ( .A(dOut_l[28]), .Z(n441) );
  HS65_LS_NAND2X7 U766 ( .A(\spm_in[SDATA][60] ), .B(n127), .Z(n403) );
  HS65_LS_OAI212X5 U767 ( .A(n132), .B(n441), .C(n324), .D(n404), .E(n403), 
        .Z(mux_out[28]) );
  HS65_LS_IVX9 U768 ( .A(dOut_l[29]), .Z(n442) );
  HS65_LS_NAND2X7 U769 ( .A(\spm_in[SDATA][61] ), .B(n127), .Z(n405) );
  HS65_LS_OAI212X5 U770 ( .A(n132), .B(n442), .C(n323), .D(n406), .E(n405), 
        .Z(mux_out[29]) );
  HS65_LS_IVX9 U771 ( .A(dOut_l[30]), .Z(n443) );
  HS65_LS_NAND2X7 U772 ( .A(\spm_in[SDATA][62] ), .B(n127), .Z(n407) );
  HS65_LS_OAI212X5 U773 ( .A(n132), .B(n443), .C(n324), .D(n408), .E(n407), 
        .Z(mux_out[30]) );
  HS65_LS_IVX9 U774 ( .A(dOut_l[31]), .Z(n444) );
  HS65_LS_NAND2X7 U775 ( .A(\spm_in[SDATA][63] ), .B(n127), .Z(n409) );
  HS65_LS_OAI212X5 U776 ( .A(n132), .B(n444), .C(n323), .D(n410), .E(n409), 
        .Z(mux_out[31]) );
  HS65_LS_MUX21I1X6 U777 ( .D0(n413), .D1(\spm_in[SDATA][0] ), .S0(n136), .Z(
        n718) );
  HS65_LS_MUX21I1X6 U778 ( .D0(n414), .D1(\spm_in[SDATA][1] ), .S0(n136), .Z(
        n717) );
  HS65_LS_MUX21I1X6 U779 ( .D0(n415), .D1(\spm_in[SDATA][2] ), .S0(n134), .Z(
        n716) );
  HS65_LS_MUX21I1X6 U780 ( .D0(n416), .D1(\spm_in[SDATA][3] ), .S0(n137), .Z(
        n715) );
  HS65_LS_MUX21I1X6 U781 ( .D0(n417), .D1(\spm_in[SDATA][4] ), .S0(n134), .Z(
        n714) );
  HS65_LS_MUX21I1X6 U782 ( .D0(n418), .D1(\spm_in[SDATA][5] ), .S0(n137), .Z(
        n713) );
  HS65_LS_MUX21I1X6 U783 ( .D0(n419), .D1(\spm_in[SDATA][6] ), .S0(n136), .Z(
        n712) );
  HS65_LS_MUX21I1X6 U784 ( .D0(n420), .D1(\spm_in[SDATA][7] ), .S0(n134), .Z(
        n711) );
  HS65_LS_MUX21I1X6 U785 ( .D0(n421), .D1(\spm_in[SDATA][8] ), .S0(n137), .Z(
        n710) );
  HS65_LS_MUX21I1X6 U786 ( .D0(n422), .D1(\spm_in[SDATA][9] ), .S0(n136), .Z(
        n709) );
  HS65_LS_MUX21I1X6 U787 ( .D0(n423), .D1(\spm_in[SDATA][10] ), .S0(n134), .Z(
        n708) );
  HS65_LS_MUX21I1X6 U788 ( .D0(n424), .D1(\spm_in[SDATA][11] ), .S0(n137), .Z(
        n707) );
  HS65_LS_MUX21I1X6 U789 ( .D0(n425), .D1(\spm_in[SDATA][12] ), .S0(n136), .Z(
        n706) );
  HS65_LS_MUX21I1X6 U790 ( .D0(n426), .D1(\spm_in[SDATA][13] ), .S0(n134), .Z(
        n705) );
  HS65_LS_MUX21I1X6 U791 ( .D0(n427), .D1(\spm_in[SDATA][14] ), .S0(n137), .Z(
        n704) );
  HS65_LS_MUX21I1X6 U792 ( .D0(n428), .D1(\spm_in[SDATA][15] ), .S0(n134), .Z(
        n703) );
  HS65_LS_MUX21I1X6 U793 ( .D0(n429), .D1(\spm_in[SDATA][16] ), .S0(n137), .Z(
        n702) );
  HS65_LS_MUX21I1X6 U794 ( .D0(n430), .D1(\spm_in[SDATA][17] ), .S0(n136), .Z(
        n701) );
  HS65_LS_MUX21I1X6 U795 ( .D0(n431), .D1(\spm_in[SDATA][18] ), .S0(n134), .Z(
        n700) );
  HS65_LS_MUX21I1X6 U796 ( .D0(n432), .D1(\spm_in[SDATA][19] ), .S0(n137), .Z(
        n699) );
  HS65_LS_MUX21I1X6 U797 ( .D0(n433), .D1(\spm_in[SDATA][20] ), .S0(n136), .Z(
        n698) );
  HS65_LS_MUX21I1X6 U798 ( .D0(n434), .D1(\spm_in[SDATA][21] ), .S0(n134), .Z(
        n697) );
  HS65_LS_MUX21I1X6 U799 ( .D0(n435), .D1(\spm_in[SDATA][22] ), .S0(n137), .Z(
        n696) );
  HS65_LS_MUX21I1X6 U800 ( .D0(n436), .D1(\spm_in[SDATA][23] ), .S0(n136), .Z(
        n695) );
  HS65_LS_MUX21I1X6 U801 ( .D0(n437), .D1(\spm_in[SDATA][24] ), .S0(n134), .Z(
        n694) );
  HS65_LS_MUX21I1X6 U802 ( .D0(n438), .D1(\spm_in[SDATA][25] ), .S0(n137), .Z(
        n693) );
  HS65_LS_MUX21I1X6 U803 ( .D0(n439), .D1(\spm_in[SDATA][26] ), .S0(n136), .Z(
        n692) );
  HS65_LS_MUX21I1X6 U804 ( .D0(n440), .D1(\spm_in[SDATA][27] ), .S0(n136), .Z(
        n691) );
  HS65_LS_MUX21I1X6 U805 ( .D0(n441), .D1(\spm_in[SDATA][28] ), .S0(n134), .Z(
        n690) );
  HS65_LS_MUX21I1X6 U806 ( .D0(n442), .D1(\spm_in[SDATA][29] ), .S0(n137), .Z(
        n689) );
  HS65_LS_MUX21I1X6 U807 ( .D0(n443), .D1(\spm_in[SDATA][30] ), .S0(n136), .Z(
        n688) );
  HS65_LS_MUX21I1X6 U808 ( .D0(n444), .D1(\spm_in[SDATA][31] ), .S0(n134), .Z(
        n687) );
  HS65_LS_IVX9 U809 ( .A(\phase_next[1] ), .Z(n455) );
  HS65_LS_AO33X18 U810 ( .A(n462), .B(n18), .C(n120), .D(\phase_next[1] ), .E(
        n448), .F(n447), .Z(n464) );
  HS65_LS_IVX9 U811 ( .A(phitOut1[0]), .Z(n468) );
  HS65_LS_IVX9 U812 ( .A(phitOut0[0]), .Z(n467) );
  HS65_LS_IVX9 U813 ( .A(phitOut1[1]), .Z(n471) );
  HS65_LS_IVX9 U814 ( .A(phitOut0[1]), .Z(n470) );
  HS65_LS_IVX9 U815 ( .A(phitOut1[2]), .Z(n475) );
  HS65_LS_IVX9 U816 ( .A(phitOut0[2]), .Z(n474) );
  HS65_LS_IVX9 U817 ( .A(phitOut1[3]), .Z(n478) );
  HS65_LS_IVX9 U818 ( .A(phitOut0[3]), .Z(n477) );
  HS65_LS_IVX9 U819 ( .A(phitOut1[4]), .Z(n481) );
  HS65_LS_IVX9 U820 ( .A(phitOut0[4]), .Z(n480) );
  HS65_LS_OAI212X5 U821 ( .A(n116), .B(n481), .C(n570), .D(n480), .E(n479), 
        .Z(pkt_out[4]) );
  HS65_LS_IVX9 U822 ( .A(phitOut1[5]), .Z(n484) );
  HS65_LS_IVX9 U823 ( .A(phitOut0[5]), .Z(n483) );
  HS65_LS_OAI212X5 U824 ( .A(n114), .B(n484), .C(n526), .D(n483), .E(n482), 
        .Z(pkt_out[5]) );
  HS65_LS_IVX9 U825 ( .A(phitOut1[6]), .Z(n487) );
  HS65_LS_IVX9 U826 ( .A(phitOut0[6]), .Z(n486) );
  HS65_LS_IVX9 U827 ( .A(phitOut1[7]), .Z(n490) );
  HS65_LS_IVX9 U828 ( .A(phitOut0[7]), .Z(n489) );
  HS65_LS_OAI212X5 U829 ( .A(n114), .B(n490), .C(n526), .D(n489), .E(n488), 
        .Z(pkt_out[7]) );
  HS65_LS_IVX9 U830 ( .A(phitOut1[8]), .Z(n493) );
  HS65_LS_IVX9 U831 ( .A(phitOut0[8]), .Z(n492) );
  HS65_LS_OAI212X5 U832 ( .A(n114), .B(n493), .C(n526), .D(n492), .E(n491), 
        .Z(pkt_out[8]) );
  HS65_LS_IVX9 U833 ( .A(phitOut1[9]), .Z(n496) );
  HS65_LS_IVX9 U834 ( .A(phitOut0[9]), .Z(n495) );
  HS65_LS_OAI212X5 U835 ( .A(n29), .B(n496), .C(n526), .D(n495), .E(n494), .Z(
        pkt_out[9]) );
  HS65_LS_IVX9 U836 ( .A(phitOut1[10]), .Z(n499) );
  HS65_LS_IVX9 U837 ( .A(phitOut0[10]), .Z(n498) );
  HS65_LS_IVX9 U838 ( .A(phitOut1[11]), .Z(n502) );
  HS65_LS_IVX9 U839 ( .A(phitOut0[11]), .Z(n501) );
  HS65_LS_IVX9 U840 ( .A(phitOut1[12]), .Z(n505) );
  HS65_LS_IVX9 U841 ( .A(phitOut0[12]), .Z(n504) );
  HS65_LS_OAI212X5 U842 ( .A(n30), .B(n505), .C(n526), .D(n504), .E(n503), .Z(
        pkt_out[12]) );
  HS65_LS_IVX9 U843 ( .A(phitOut1[13]), .Z(n508) );
  HS65_LS_IVX9 U844 ( .A(phitOut0[13]), .Z(n507) );
  HS65_LS_OAI212X5 U845 ( .A(n508), .B(n114), .C(n526), .D(n507), .E(n506), 
        .Z(pkt_out[13]) );
  HS65_LS_IVX9 U846 ( .A(phitOut1[14]), .Z(n511) );
  HS65_LS_IVX9 U847 ( .A(phitOut0[14]), .Z(n510) );
  HS65_LS_OAI212X5 U848 ( .A(n511), .B(n114), .C(n526), .D(n510), .E(n509), 
        .Z(pkt_out[14]) );
  HS65_LS_IVX9 U849 ( .A(phitOut1[15]), .Z(n514) );
  HS65_LS_IVX9 U850 ( .A(phitOut0[15]), .Z(n513) );
  HS65_LS_OAI212X5 U851 ( .A(n116), .B(n514), .C(n526), .D(n513), .E(n512), 
        .Z(pkt_out[15]) );
  HS65_LS_IVX9 U852 ( .A(phitOut1[16]), .Z(n517) );
  HS65_LS_IVX9 U853 ( .A(phitOut0[16]), .Z(n516) );
  HS65_LS_OAI212X5 U854 ( .A(n114), .B(n517), .C(n526), .D(n516), .E(n515), 
        .Z(pkt_out[16]) );
  HS65_LS_IVX9 U855 ( .A(phitOut1[17]), .Z(n520) );
  HS65_LS_IVX9 U856 ( .A(phitOut0[17]), .Z(n519) );
  HS65_LS_OAI212X5 U857 ( .A(n29), .B(n520), .C(n526), .D(n519), .E(n518), .Z(
        pkt_out[17]) );
  HS65_LS_IVX9 U858 ( .A(phitOut1[18]), .Z(n523) );
  HS65_LS_IVX9 U859 ( .A(phitOut0[18]), .Z(n522) );
  HS65_LS_OAI212X5 U860 ( .A(n30), .B(n523), .C(n526), .D(n522), .E(n521), .Z(
        pkt_out[18]) );
  HS65_LS_IVX9 U861 ( .A(phitOut1[19]), .Z(n527) );
  HS65_LS_IVX9 U862 ( .A(phitOut0[19]), .Z(n525) );
  HS65_LS_OAI212X5 U863 ( .A(n116), .B(n527), .C(n526), .D(n525), .E(n524), 
        .Z(pkt_out[19]) );
  HS65_LS_IVX9 U864 ( .A(phitOut1[20]), .Z(n530) );
  HS65_LS_IVX9 U865 ( .A(phitOut0[20]), .Z(n529) );
  HS65_LS_OAI212X5 U866 ( .A(n114), .B(n530), .C(n24), .D(n529), .E(n528), .Z(
        pkt_out[20]) );
  HS65_LS_IVX9 U867 ( .A(phitOut1[21]), .Z(n533) );
  HS65_LS_IVX9 U868 ( .A(phitOut0[21]), .Z(n532) );
  HS65_LS_OAI212X5 U869 ( .A(n116), .B(n533), .C(n23), .D(n532), .E(n531), .Z(
        pkt_out[21]) );
  HS65_LS_IVX9 U870 ( .A(phitOut1[22]), .Z(n536) );
  HS65_LS_IVX9 U871 ( .A(phitOut0[22]), .Z(n535) );
  HS65_LS_OAI212X5 U872 ( .A(n114), .B(n536), .C(n22), .D(n535), .E(n534), .Z(
        pkt_out[22]) );
  HS65_LS_IVX9 U873 ( .A(phitOut1[23]), .Z(n539) );
  HS65_LS_IVX9 U874 ( .A(phitOut0[23]), .Z(n538) );
  HS65_LS_IVX9 U875 ( .A(phitOut1[24]), .Z(n542) );
  HS65_LS_IVX9 U876 ( .A(phitOut0[24]), .Z(n541) );
  HS65_LS_IVX9 U877 ( .A(phitOut1[25]), .Z(n545) );
  HS65_LS_IVX9 U878 ( .A(phitOut0[25]), .Z(n544) );
  HS65_LS_OAI212X5 U879 ( .A(n116), .B(n545), .C(n24), .D(n544), .E(n543), .Z(
        pkt_out[25]) );
  HS65_LS_IVX9 U880 ( .A(phitOut1[26]), .Z(n548) );
  HS65_LS_IVX9 U881 ( .A(phitOut0[26]), .Z(n547) );
  HS65_LS_OAI212X5 U882 ( .A(n114), .B(n548), .C(n22), .D(n547), .E(n546), .Z(
        pkt_out[26]) );
  HS65_LS_IVX9 U883 ( .A(phitOut1[27]), .Z(n551) );
  HS65_LS_IVX9 U884 ( .A(phitOut0[27]), .Z(n550) );
  HS65_LS_OAI212X5 U885 ( .A(n118), .B(n551), .C(n23), .D(n550), .E(n549), .Z(
        pkt_out[27]) );
  HS65_LS_IVX9 U886 ( .A(phitOut1[28]), .Z(n554) );
  HS65_LS_IVX9 U887 ( .A(phitOut0[28]), .Z(n553) );
  HS65_LS_OAI212X5 U888 ( .A(n29), .B(n554), .C(n22), .D(n553), .E(n552), .Z(
        pkt_out[28]) );
  HS65_LS_IVX9 U889 ( .A(phitOut1[29]), .Z(n557) );
  HS65_LS_IVX9 U890 ( .A(phitOut0[29]), .Z(n556) );
  HS65_LS_OAI212X5 U891 ( .A(n29), .B(n557), .C(n24), .D(n556), .E(n555), .Z(
        pkt_out[29]) );
  HS65_LS_IVX9 U892 ( .A(phitOut1[30]), .Z(n560) );
  HS65_LS_IVX9 U893 ( .A(phitOut0[30]), .Z(n559) );
  HS65_LS_OAI212X5 U894 ( .A(n29), .B(n560), .C(n23), .D(n559), .E(n558), .Z(
        pkt_out[30]) );
  HS65_LS_IVX9 U895 ( .A(phitOut1[31]), .Z(n563) );
  HS65_LS_IVX9 U896 ( .A(phitOut0[31]), .Z(n562) );
  HS65_LS_OAI212X5 U897 ( .A(n118), .B(n563), .C(n23), .D(n562), .E(n561), .Z(
        pkt_out[31]) );
  HS65_LS_IVX9 U898 ( .A(phitOut1[32]), .Z(n566) );
  HS65_LS_IVX9 U899 ( .A(phitOut0[32]), .Z(n565) );
  HS65_LS_OAI212X5 U900 ( .A(n118), .B(n566), .C(n22), .D(n565), .E(n564), .Z(
        pkt_out[32]) );
  HS65_LS_IVX9 U901 ( .A(phitOut1[33]), .Z(n571) );
  HS65_LS_IVX9 U902 ( .A(phitOut0[33]), .Z(n569) );
  HS65_LS_OAI212X5 U903 ( .A(n114), .B(n571), .C(n24), .D(n569), .E(n568), .Z(
        pkt_out[33]) );
  HS65_LS_IVX9 U904 ( .A(phitOut1[34]), .Z(n575) );
  HS65_LS_IVX9 U905 ( .A(flit_buf[64]), .Z(n578) );
  HS65_LS_OAI22X6 U906 ( .A(n355), .B(n579), .C(n592), .D(n578), .Z(
        \spm_out[MADDR][0] ) );
  HS65_LS_IVX9 U907 ( .A(flit_buf[65]), .Z(n580) );
  HS65_LS_OAI22X6 U908 ( .A(n355), .B(n581), .C(n592), .D(n580), .Z(
        \spm_out[MADDR][1] ) );
  HS65_LS_IVX9 U909 ( .A(flit_buf[66]), .Z(n582) );
  HS65_LS_OAI22X6 U910 ( .A(n355), .B(n583), .C(n592), .D(n582), .Z(
        \spm_out[MADDR][2] ) );
  HS65_LS_IVX9 U911 ( .A(flit_buf[67]), .Z(n584) );
  HS65_LS_OAI22X6 U912 ( .A(n355), .B(n585), .C(n592), .D(n584), .Z(
        \spm_out[MADDR][3] ) );
  HS65_LS_IVX9 U913 ( .A(flit_buf[68]), .Z(n586) );
  HS65_LS_OAI22X6 U914 ( .A(n355), .B(n587), .C(n592), .D(n586), .Z(
        \spm_out[MADDR][4] ) );
  HS65_LS_IVX9 U915 ( .A(flit_buf[69]), .Z(n588) );
  HS65_LS_OAI22X6 U916 ( .A(n355), .B(n589), .C(n592), .D(n588), .Z(
        \spm_out[MADDR][5] ) );
  HS65_LS_IVX9 U917 ( .A(flit_buf[70]), .Z(n590) );
  HS65_LS_OAI22X6 U918 ( .A(n591), .B(n355), .C(n592), .D(n590), .Z(
        \spm_out[MADDR][6] ) );
  HS65_LS_IVX9 U919 ( .A(n592), .Z(\spm_out[MCMD][0] ) );
  HS65_LS_IVX9 U920 ( .A(n593), .Z(n595) );
  HS65_LS_OAI112X5 U921 ( .A(n868), .B(n595), .C(n867), .D(n594), .Z(
        \proc_out[SCMDACCEPT] ) );
endmodule


module latch_controller_1_35 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_35 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n3, n4, n5, n6;
  assign N0 = preset;

  latch_controller_1_35 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n4), .RN(n3), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n3), .Z(n5) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n6), .B(n5), .Z(N5) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_IVX9 U3 ( .A(lt_enable), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(N0), .Z(n3) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n4), .Z(lt_gated) );
endmodule


module latch_controller_1_34 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_34 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n3, n4, n5, n6;
  assign N0 = preset;

  latch_controller_1_34 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n4), .RN(n3), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n3), .Z(n5) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n6), .B(n5), .Z(N5) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_IVX9 U3 ( .A(lt_enable), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(N0), .Z(n3) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n4), .Z(lt_gated) );
endmodule


module latch_controller_1_33 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_33 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n3, n4, n5, n6;
  assign N0 = preset;

  latch_controller_1_33 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n4), .RN(n3), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n3), .Z(n5) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n6), .B(n5), .Z(N5) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_IVX9 U3 ( .A(lt_enable), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(N0), .Z(n3) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n4), .Z(lt_gated) );
endmodule


module latch_controller_1_32 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_32 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n3, n4, n5, n6;
  assign N0 = preset;

  latch_controller_1_32 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n4), .RN(n3), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n3), .Z(n5) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n6), .B(n5), .Z(N5) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_IVX9 U3 ( .A(lt_enable), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(N0), .Z(n3) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n4), .Z(lt_gated) );
endmodule


module latch_controller_1_31 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_NOR2AX3 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_31 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n3, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_31 controller ( .preset(n3), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLRQX18 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(n3), .Z(n7) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_LDHQX18 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX18 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX18 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX18 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX18 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX18 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX18 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX18 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX18 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX18 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX18 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX18 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX18 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX18 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX18 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX4 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX4 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX18 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX18 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX18 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX18 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX18 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX18 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX4 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX4 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX4 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX18 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX18 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX18 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX18 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX18 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX18 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX18 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX18 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_NAND2X5 U3 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
  HS65_LS_IVX9 U4 ( .A(n4), .Z(n3) );
  HS65_LS_IVX9 U5 ( .A(lt_enable), .Z(n5) );
  HS65_LS_IVX9 U9 ( .A(N0), .Z(n4) );
endmodule


module hpu_comb_0_0_3 ( data_valid, data_in, preset, data_out, sel );
  input [34:0] data_in;
  output [34:0] data_out;
  output [4:0] sel;
  input data_valid, preset;
  wire   data_in_34, data_in_33, data_in_32, \data_in[31] , \data_in[30] ,
         \data_in[29] , \data_in[28] , \data_in[27] , \data_in[26] ,
         \data_in[25] , \data_in[24] , \data_in[23] , \data_in[22] ,
         \data_in[21] , \data_in[20] , \data_in[19] , \data_in[18] ,
         \data_in[17] , \data_in[16] , N23, N25, N26, N27, N28, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n22,
         n23, n24;
  assign data_out[34] = data_in_34;
  assign data_in_34 = data_in[34];
  assign data_out[33] = data_in_33;
  assign data_in_33 = data_in[33];
  assign data_out[32] = data_in_32;
  assign data_in_32 = data_in[32];
  assign data_out[31] = \data_in[31] ;
  assign \data_in[31]  = data_in[31];
  assign data_out[30] = \data_in[30] ;
  assign \data_in[30]  = data_in[30];
  assign data_out[29] = \data_in[29] ;
  assign \data_in[29]  = data_in[29];
  assign data_out[28] = \data_in[28] ;
  assign \data_in[28]  = data_in[28];
  assign data_out[27] = \data_in[27] ;
  assign \data_in[27]  = data_in[27];
  assign data_out[26] = \data_in[26] ;
  assign \data_in[26]  = data_in[26];
  assign data_out[25] = \data_in[25] ;
  assign \data_in[25]  = data_in[25];
  assign data_out[24] = \data_in[24] ;
  assign \data_in[24]  = data_in[24];
  assign data_out[23] = \data_in[23] ;
  assign \data_in[23]  = data_in[23];
  assign data_out[22] = \data_in[22] ;
  assign \data_in[22]  = data_in[22];
  assign data_out[21] = \data_in[21] ;
  assign \data_in[21]  = data_in[21];
  assign data_out[20] = \data_in[20] ;
  assign \data_in[20]  = data_in[20];
  assign data_out[19] = \data_in[19] ;
  assign \data_in[19]  = data_in[19];
  assign data_out[18] = \data_in[18] ;
  assign \data_in[18]  = data_in[18];
  assign data_out[17] = \data_in[17] ;
  assign \data_in[17]  = data_in[17];
  assign data_out[16] = \data_in[16] ;
  assign \data_in[16]  = data_in[16];
  assign sel[0] = 1'b0;

  HS65_LS_LDHQX9 \sel_reg[4]  ( .G(N23), .D(N28), .Q(sel[4]) );
  HS65_LS_LDHQX9 \sel_reg[3]  ( .G(N23), .D(N27), .Q(sel[3]) );
  HS65_LS_LDHQX9 \sel_reg[2]  ( .G(N23), .D(N26), .Q(sel[2]) );
  HS65_LS_LDHQX9 \sel_reg[1]  ( .G(N23), .D(N25), .Q(sel[1]) );
  HS65_LS_NAND3AX6 U4 ( .A(preset), .B(n23), .C(n2), .Z(n22) );
  HS65_LS_OAI22X6 U5 ( .A(n9), .B(n24), .C(n2), .D(n11), .Z(data_out[7]) );
  HS65_LS_OAI22X6 U6 ( .A(n24), .B(n16), .C(n2), .D(n18), .Z(data_out[0]) );
  HS65_LS_OAI22X6 U7 ( .A(n24), .B(n15), .C(n2), .D(n17), .Z(data_out[1]) );
  HS65_LS_OAI22X6 U8 ( .A(n24), .B(n14), .C(n2), .D(n16), .Z(data_out[2]) );
  HS65_LS_OAI22X6 U9 ( .A(n24), .B(n13), .C(n2), .D(n15), .Z(data_out[3]) );
  HS65_LS_OAI22X6 U10 ( .A(n24), .B(n12), .C(n2), .D(n14), .Z(data_out[4]) );
  HS65_LS_OAI22X6 U11 ( .A(n24), .B(n11), .C(n2), .D(n13), .Z(data_out[5]) );
  HS65_LS_OAI22X6 U12 ( .A(n24), .B(n10), .C(n2), .D(n12), .Z(data_out[6]) );
  HS65_LS_OAI22X6 U13 ( .A(n24), .B(n8), .C(n2), .D(n10), .Z(data_out[8]) );
  HS65_LS_OAI22X6 U14 ( .A(n24), .B(n7), .C(n2), .D(n9), .Z(data_out[9]) );
  HS65_LS_OAI22X6 U15 ( .A(n24), .B(n6), .C(n2), .D(n8), .Z(data_out[10]) );
  HS65_LS_OAI22X6 U16 ( .A(n24), .B(n5), .C(n2), .D(n7), .Z(data_out[11]) );
  HS65_LS_OAI22X6 U17 ( .A(n24), .B(n4), .C(n2), .D(n6), .Z(data_out[12]) );
  HS65_LS_OAI22X6 U18 ( .A(n24), .B(n3), .C(n2), .D(n5), .Z(data_out[13]) );
  HS65_LS_IVX9 U19 ( .A(n24), .Z(n2) );
  HS65_LS_NOR3X4 U20 ( .A(n23), .B(preset), .C(n24), .Z(N28) );
  HS65_LS_NOR3X4 U21 ( .A(n22), .B(n17), .C(n18), .Z(N27) );
  HS65_LS_NAND2X7 U22 ( .A(n17), .B(n18), .Z(n23) );
  HS65_LS_NOR2X6 U23 ( .A(n2), .B(n4), .Z(data_out[14]) );
  HS65_LS_NOR2X6 U24 ( .A(n2), .B(n3), .Z(data_out[15]) );
  HS65_LS_NAND2X14 U25 ( .A(data_in_34), .B(data_in_33), .Z(n24) );
  HS65_LS_IVX9 U26 ( .A(data_in[1]), .Z(n17) );
  HS65_LS_IVX9 U27 ( .A(data_in[0]), .Z(n18) );
  HS65_LS_NOR2X6 U28 ( .A(data_in[1]), .B(n22), .Z(N25) );
  HS65_LS_NOR2X6 U29 ( .A(data_in[0]), .B(n22), .Z(N26) );
  HS65_LS_IVX9 U30 ( .A(data_in[9]), .Z(n9) );
  HS65_LS_IVX9 U31 ( .A(data_in[2]), .Z(n16) );
  HS65_LS_IVX9 U32 ( .A(data_in[3]), .Z(n15) );
  HS65_LS_IVX9 U33 ( .A(data_in[4]), .Z(n14) );
  HS65_LS_IVX9 U34 ( .A(data_in[5]), .Z(n13) );
  HS65_LS_IVX9 U35 ( .A(data_in[6]), .Z(n12) );
  HS65_LS_IVX9 U36 ( .A(data_in[7]), .Z(n11) );
  HS65_LS_IVX9 U37 ( .A(data_in[8]), .Z(n10) );
  HS65_LS_IVX9 U38 ( .A(data_in[10]), .Z(n8) );
  HS65_LS_IVX9 U39 ( .A(data_in[11]), .Z(n7) );
  HS65_LS_IVX9 U40 ( .A(data_in[12]), .Z(n6) );
  HS65_LS_IVX9 U41 ( .A(data_in[13]), .Z(n5) );
  HS65_LS_IVX9 U42 ( .A(data_in[14]), .Z(n4) );
  HS65_LS_IVX9 U43 ( .A(data_in[15]), .Z(n3) );
  HS65_LS_CB4I6X9 U44 ( .A(n2), .B(n1), .C(data_valid), .D(preset), .Z(N23) );
  HS65_LS_IVX9 U45 ( .A(data_in_34), .Z(n1) );
endmodule


module latch_controller_1_15 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_15 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_15 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n7) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_IVX9 U3 ( .A(N0), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_0_0_3 ( preset, .chan_in_f({\chan_in_f[REQ] , \chan_in_f[DATA][34] , 
        \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , 
        \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , 
        \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , 
        \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , 
        \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , 
        \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , 
        \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , 
        \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , 
        \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , 
        \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , 
        \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , 
        \chan_in_f[DATA][0] }), .chan_in_b(\chan_in_b[ACK] ), .chan_out_f({
        \chan_out_f[REQ] , \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , 
        \chan_out_f[DATA][32] , \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , 
        \chan_out_f[DATA][29] , \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , 
        \chan_out_f[DATA][26] , \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , 
        \chan_out_f[DATA][23] , \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , 
        \chan_out_f[DATA][20] , \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , 
        \chan_out_f[DATA][17] , \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , 
        \chan_out_f[DATA][14] , \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , 
        \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , 
        \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , 
        \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , 
        \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), 
    .chan_out_b(\chan_out_b[ACK] ), sel );
  output [4:0] sel;
  input preset, \chan_in_f[REQ] , \chan_in_f[DATA][34] , \chan_in_f[DATA][33] ,
         \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , \chan_in_f[DATA][30] ,
         \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , \chan_in_f[DATA][27] ,
         \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , \chan_in_f[DATA][24] ,
         \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , \chan_in_f[DATA][21] ,
         \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , \chan_in_f[DATA][18] ,
         \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , \chan_in_f[DATA][15] ,
         \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , \chan_in_f[DATA][12] ,
         \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , \chan_in_f[DATA][9] ,
         \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , \chan_in_f[DATA][6] ,
         \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , \chan_in_f[DATA][3] ,
         \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , \chan_in_f[DATA][0] ,
         \chan_out_b[ACK] ;
  output \chan_in_b[ACK] , \chan_out_f[REQ] , \chan_out_f[DATA][34] ,
         \chan_out_f[DATA][33] , \chan_out_f[DATA][32] ,
         \chan_out_f[DATA][31] , \chan_out_f[DATA][30] ,
         \chan_out_f[DATA][29] , \chan_out_f[DATA][28] ,
         \chan_out_f[DATA][27] , \chan_out_f[DATA][26] ,
         \chan_out_f[DATA][25] , \chan_out_f[DATA][24] ,
         \chan_out_f[DATA][23] , \chan_out_f[DATA][22] ,
         \chan_out_f[DATA][21] , \chan_out_f[DATA][20] ,
         \chan_out_f[DATA][19] , \chan_out_f[DATA][18] ,
         \chan_out_f[DATA][17] , \chan_out_f[DATA][16] ,
         \chan_out_f[DATA][15] , \chan_out_f[DATA][14] ,
         \chan_out_f[DATA][13] , \chan_out_f[DATA][12] ,
         \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] ,
         \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] ,
         \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] ,
         \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] ;
  wire   \chan_internal_f[REQ] , \chan_internal_f[DATA][34] ,
         \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] ,
         \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] ,
         \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] ,
         \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] ,
         \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] ,
         \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] ,
         \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] ,
         \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] ,
         \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] ,
         \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] ,
         \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] ,
         \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] ,
         \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] ,
         \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] ,
         \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] ,
         \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] ,
         \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] , req_n, lt_en,
         n1, n2, n3, n4, n5, n6, n7;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign sel[0] = 1'b0;

  hpu_comb_0_0_3 hpu_combinatorial ( .data_valid(lt_en), .data_in({
        \chan_in_f[DATA][34] , \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , 
        \chan_in_f[DATA][31] , \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , 
        \chan_in_f[DATA][28] , \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , 
        \chan_in_f[DATA][25] , \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , 
        \chan_in_f[DATA][22] , \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , 
        \chan_in_f[DATA][19] , \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , 
        \chan_in_f[DATA][16] , \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , 
        \chan_in_f[DATA][13] , \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , 
        \chan_in_f[DATA][10] , \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , 
        \chan_in_f[DATA][7] , \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , 
        \chan_in_f[DATA][4] , \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , 
        \chan_in_f[DATA][1] , \chan_in_f[DATA][0] }), .preset(n7), .data_out({
        \chan_internal_f[DATA][34] , \chan_internal_f[DATA][33] , 
        \chan_internal_f[DATA][32] , \chan_internal_f[DATA][31] , 
        \chan_internal_f[DATA][30] , \chan_internal_f[DATA][29] , 
        \chan_internal_f[DATA][28] , \chan_internal_f[DATA][27] , 
        \chan_internal_f[DATA][26] , \chan_internal_f[DATA][25] , 
        \chan_internal_f[DATA][24] , \chan_internal_f[DATA][23] , 
        \chan_internal_f[DATA][22] , \chan_internal_f[DATA][21] , 
        \chan_internal_f[DATA][20] , \chan_internal_f[DATA][19] , 
        \chan_internal_f[DATA][18] , \chan_internal_f[DATA][17] , 
        \chan_internal_f[DATA][16] , \chan_internal_f[DATA][15] , 
        \chan_internal_f[DATA][14] , \chan_internal_f[DATA][13] , 
        \chan_internal_f[DATA][12] , \chan_internal_f[DATA][11] , 
        \chan_internal_f[DATA][10] , \chan_internal_f[DATA][9] , 
        \chan_internal_f[DATA][8] , \chan_internal_f[DATA][7] , 
        \chan_internal_f[DATA][6] , \chan_internal_f[DATA][5] , 
        \chan_internal_f[DATA][4] , \chan_internal_f[DATA][3] , 
        \chan_internal_f[DATA][2] , \chan_internal_f[DATA][1] , 
        \chan_internal_f[DATA][0] }), .sel({sel[4:1], SYNOPSYS_UNCONNECTED__0}) );
  channel_latch_1_xxxxxxxxx_15 token_latch ( .preset(n7), .left_in({
        \chan_internal_f[REQ] , \chan_internal_f[DATA][34] , 
        \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] , 
        \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] , 
        \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] , 
        \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] , 
        \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] , 
        \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] , 
        \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] , 
        \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] , 
        \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] , 
        \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] , 
        \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] , 
        \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] , 
        \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] , 
        \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] , 
        \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] , 
        \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] , 
        \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] }), .left_out(
        \chan_in_b[ACK] ), .right_out({\chan_out_f[REQ] , 
        \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , \chan_out_f[DATA][32] , 
        \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , \chan_out_f[DATA][29] , 
        \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , \chan_out_f[DATA][26] , 
        \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , \chan_out_f[DATA][23] , 
        \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , \chan_out_f[DATA][20] , 
        \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , \chan_out_f[DATA][17] , 
        \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , \chan_out_f[DATA][14] , 
        \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , \chan_out_f[DATA][11] , 
        \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , \chan_out_f[DATA][8] , 
        \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , \chan_out_f[DATA][5] , 
        \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , \chan_out_f[DATA][2] , 
        \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), .right_in(
        \chan_out_b[ACK] ), .lt_enable(lt_en) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chan_internal_f[REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(\chan_in_f[REQ] ), .Z(req_n) );
  HS65_LS_BFX9 U1 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U2 ( .A(n3), .Z(n2) );
  HS65_LS_BFX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_BFX9 U4 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U6 ( .A(req_n), .Z(n6) );
  HS65_LS_BFX9 U7 ( .A(preset), .Z(n7) );
endmodule


module hpu_comb_0_2_3 ( data_valid, data_in, preset, data_out, sel );
  input [34:0] data_in;
  output [34:0] data_out;
  output [4:0] sel;
  input data_valid, preset;
  wire   data_in_34, data_in_33, data_in_32, \data_in[31] , \data_in[30] ,
         \data_in[29] , \data_in[28] , \data_in[27] , \data_in[26] ,
         \data_in[25] , \data_in[24] , \data_in[23] , \data_in[22] ,
         \data_in[21] , \data_in[20] , \data_in[19] , \data_in[18] ,
         \data_in[17] , \data_in[16] , N26, N27, N28, N30, N31, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n15, n16, n17, n18;
  assign data_out[34] = data_in_34;
  assign data_in_34 = data_in[34];
  assign data_out[33] = data_in_33;
  assign data_in_33 = data_in[33];
  assign data_out[32] = data_in_32;
  assign data_in_32 = data_in[32];
  assign data_out[31] = \data_in[31] ;
  assign \data_in[31]  = data_in[31];
  assign data_out[30] = \data_in[30] ;
  assign \data_in[30]  = data_in[30];
  assign data_out[29] = \data_in[29] ;
  assign \data_in[29]  = data_in[29];
  assign data_out[28] = \data_in[28] ;
  assign \data_in[28]  = data_in[28];
  assign data_out[27] = \data_in[27] ;
  assign \data_in[27]  = data_in[27];
  assign data_out[26] = \data_in[26] ;
  assign \data_in[26]  = data_in[26];
  assign data_out[25] = \data_in[25] ;
  assign \data_in[25]  = data_in[25];
  assign data_out[24] = \data_in[24] ;
  assign \data_in[24]  = data_in[24];
  assign data_out[23] = \data_in[23] ;
  assign \data_in[23]  = data_in[23];
  assign data_out[22] = \data_in[22] ;
  assign \data_in[22]  = data_in[22];
  assign data_out[21] = \data_in[21] ;
  assign \data_in[21]  = data_in[21];
  assign data_out[20] = \data_in[20] ;
  assign \data_in[20]  = data_in[20];
  assign data_out[19] = \data_in[19] ;
  assign \data_in[19]  = data_in[19];
  assign data_out[18] = \data_in[18] ;
  assign \data_in[18]  = data_in[18];
  assign data_out[17] = \data_in[17] ;
  assign \data_in[17]  = data_in[17];
  assign data_out[16] = \data_in[16] ;
  assign \data_in[16]  = data_in[16];
  assign sel[2] = 1'b0;

  HS65_LS_LDHQX9 \sel_reg[4]  ( .G(N26), .D(N31), .Q(sel[4]) );
  HS65_LS_LDHQX9 \sel_reg[3]  ( .G(N26), .D(N30), .Q(sel[3]) );
  HS65_LS_LDHQX9 \sel_reg[1]  ( .G(N26), .D(N28), .Q(sel[1]) );
  HS65_LS_LDHQX9 \sel_reg[0]  ( .G(N26), .D(N27), .Q(sel[0]) );
  HS65_LS_OAI22X6 U4 ( .A(n18), .B(n9), .C(n2), .D(n10), .Z(data_out[0]) );
  HS65_LS_OAI22X6 U5 ( .A(n18), .B(n8), .C(n2), .D(n9), .Z(data_out[2]) );
  HS65_LS_OAI22X6 U6 ( .A(n18), .B(n7), .C(n2), .D(n8), .Z(data_out[4]) );
  HS65_LS_OAI22X6 U7 ( .A(n18), .B(n6), .C(n2), .D(n7), .Z(data_out[6]) );
  HS65_LS_OAI22X6 U8 ( .A(n18), .B(n5), .C(n2), .D(n6), .Z(data_out[8]) );
  HS65_LS_OAI22X6 U9 ( .A(n18), .B(n4), .C(n2), .D(n5), .Z(data_out[10]) );
  HS65_LS_OAI22X6 U10 ( .A(n18), .B(n3), .C(n2), .D(n4), .Z(data_out[12]) );
  HS65_LS_NAND3AX6 U11 ( .A(preset), .B(n17), .C(n2), .Z(n16) );
  HS65_LS_NOR3X4 U12 ( .A(n17), .B(preset), .C(n18), .Z(N31) );
  HS65_LS_IVX9 U13 ( .A(n18), .Z(n2) );
  HS65_LS_NOR3X4 U14 ( .A(n16), .B(n10), .C(n15), .Z(N30) );
  HS65_LS_NOR2AX3 U15 ( .A(n15), .B(n16), .Z(N28) );
  HS65_LS_NOR2X6 U16 ( .A(n2), .B(n3), .Z(data_out[14]) );
  HS65_LS_NAND2X14 U17 ( .A(data_in_34), .B(data_in_33), .Z(n18) );
  HS65_LS_IVX9 U18 ( .A(data_in[0]), .Z(n10) );
  HS65_LS_NAND2X7 U19 ( .A(data_in[1]), .B(n10), .Z(n17) );
  HS65_LS_NOR2X6 U20 ( .A(n10), .B(data_in[1]), .Z(n15) );
  HS65_LS_NOR2X6 U21 ( .A(data_in[0]), .B(n16), .Z(N27) );
  HS65_LS_IVX9 U22 ( .A(data_in[2]), .Z(n9) );
  HS65_LS_IVX9 U23 ( .A(data_in[4]), .Z(n8) );
  HS65_LS_IVX9 U24 ( .A(data_in[6]), .Z(n7) );
  HS65_LS_IVX9 U25 ( .A(data_in[8]), .Z(n6) );
  HS65_LS_IVX9 U26 ( .A(data_in[10]), .Z(n5) );
  HS65_LS_IVX9 U27 ( .A(data_in[12]), .Z(n4) );
  HS65_LS_IVX9 U28 ( .A(data_in[14]), .Z(n3) );
  HS65_LS_AO22X9 U29 ( .A(n2), .B(data_in[3]), .C(n18), .D(data_in[1]), .Z(
        data_out[1]) );
  HS65_LS_AO22X9 U30 ( .A(n2), .B(data_in[5]), .C(n18), .D(data_in[3]), .Z(
        data_out[3]) );
  HS65_LS_AO22X9 U31 ( .A(n2), .B(data_in[7]), .C(n18), .D(data_in[5]), .Z(
        data_out[5]) );
  HS65_LS_AO22X9 U32 ( .A(data_in[9]), .B(n2), .C(n18), .D(data_in[7]), .Z(
        data_out[7]) );
  HS65_LS_AO22X9 U33 ( .A(n2), .B(data_in[11]), .C(n18), .D(data_in[9]), .Z(
        data_out[9]) );
  HS65_LS_AO22X9 U34 ( .A(n2), .B(data_in[13]), .C(n18), .D(data_in[11]), .Z(
        data_out[11]) );
  HS65_LS_AO22X9 U35 ( .A(n2), .B(data_in[15]), .C(n18), .D(data_in[13]), .Z(
        data_out[13]) );
  HS65_LS_AND2X4 U36 ( .A(data_in[15]), .B(n18), .Z(data_out[15]) );
  HS65_LS_CB4I6X9 U37 ( .A(n2), .B(n1), .C(data_valid), .D(preset), .Z(N26) );
  HS65_LS_IVX9 U38 ( .A(data_in_34), .Z(n1) );
endmodule


module latch_controller_1_14 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_14 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_14 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n7) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_IVX9 U3 ( .A(N0), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_0_2_3 ( preset, .chan_in_f({\chan_in_f[REQ] , \chan_in_f[DATA][34] , 
        \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , 
        \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , 
        \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , 
        \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , 
        \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , 
        \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , 
        \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , 
        \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , 
        \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , 
        \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , 
        \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , 
        \chan_in_f[DATA][0] }), .chan_in_b(\chan_in_b[ACK] ), .chan_out_f({
        \chan_out_f[REQ] , \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , 
        \chan_out_f[DATA][32] , \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , 
        \chan_out_f[DATA][29] , \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , 
        \chan_out_f[DATA][26] , \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , 
        \chan_out_f[DATA][23] , \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , 
        \chan_out_f[DATA][20] , \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , 
        \chan_out_f[DATA][17] , \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , 
        \chan_out_f[DATA][14] , \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , 
        \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , 
        \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , 
        \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , 
        \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), 
    .chan_out_b(\chan_out_b[ACK] ), sel );
  output [4:0] sel;
  input preset, \chan_in_f[REQ] , \chan_in_f[DATA][34] , \chan_in_f[DATA][33] ,
         \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , \chan_in_f[DATA][30] ,
         \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , \chan_in_f[DATA][27] ,
         \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , \chan_in_f[DATA][24] ,
         \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , \chan_in_f[DATA][21] ,
         \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , \chan_in_f[DATA][18] ,
         \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , \chan_in_f[DATA][15] ,
         \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , \chan_in_f[DATA][12] ,
         \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , \chan_in_f[DATA][9] ,
         \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , \chan_in_f[DATA][6] ,
         \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , \chan_in_f[DATA][3] ,
         \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , \chan_in_f[DATA][0] ,
         \chan_out_b[ACK] ;
  output \chan_in_b[ACK] , \chan_out_f[REQ] , \chan_out_f[DATA][34] ,
         \chan_out_f[DATA][33] , \chan_out_f[DATA][32] ,
         \chan_out_f[DATA][31] , \chan_out_f[DATA][30] ,
         \chan_out_f[DATA][29] , \chan_out_f[DATA][28] ,
         \chan_out_f[DATA][27] , \chan_out_f[DATA][26] ,
         \chan_out_f[DATA][25] , \chan_out_f[DATA][24] ,
         \chan_out_f[DATA][23] , \chan_out_f[DATA][22] ,
         \chan_out_f[DATA][21] , \chan_out_f[DATA][20] ,
         \chan_out_f[DATA][19] , \chan_out_f[DATA][18] ,
         \chan_out_f[DATA][17] , \chan_out_f[DATA][16] ,
         \chan_out_f[DATA][15] , \chan_out_f[DATA][14] ,
         \chan_out_f[DATA][13] , \chan_out_f[DATA][12] ,
         \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] ,
         \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] ,
         \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] ,
         \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] ;
  wire   \chan_internal_f[REQ] , \chan_internal_f[DATA][34] ,
         \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] ,
         \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] ,
         \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] ,
         \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] ,
         \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] ,
         \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] ,
         \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] ,
         \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] ,
         \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] ,
         \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] ,
         \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] ,
         \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] ,
         \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] ,
         \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] ,
         \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] ,
         \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] ,
         \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] , req_n, lt_en,
         n1, n2, n3, n4, n5, n6, n7;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign sel[2] = 1'b0;

  hpu_comb_0_2_3 hpu_combinatorial ( .data_valid(lt_en), .data_in({
        \chan_in_f[DATA][34] , \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , 
        \chan_in_f[DATA][31] , \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , 
        \chan_in_f[DATA][28] , \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , 
        \chan_in_f[DATA][25] , \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , 
        \chan_in_f[DATA][22] , \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , 
        \chan_in_f[DATA][19] , \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , 
        \chan_in_f[DATA][16] , \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , 
        \chan_in_f[DATA][13] , \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , 
        \chan_in_f[DATA][10] , \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , 
        \chan_in_f[DATA][7] , \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , 
        \chan_in_f[DATA][4] , \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , 
        \chan_in_f[DATA][1] , \chan_in_f[DATA][0] }), .preset(n7), .data_out({
        \chan_internal_f[DATA][34] , \chan_internal_f[DATA][33] , 
        \chan_internal_f[DATA][32] , \chan_internal_f[DATA][31] , 
        \chan_internal_f[DATA][30] , \chan_internal_f[DATA][29] , 
        \chan_internal_f[DATA][28] , \chan_internal_f[DATA][27] , 
        \chan_internal_f[DATA][26] , \chan_internal_f[DATA][25] , 
        \chan_internal_f[DATA][24] , \chan_internal_f[DATA][23] , 
        \chan_internal_f[DATA][22] , \chan_internal_f[DATA][21] , 
        \chan_internal_f[DATA][20] , \chan_internal_f[DATA][19] , 
        \chan_internal_f[DATA][18] , \chan_internal_f[DATA][17] , 
        \chan_internal_f[DATA][16] , \chan_internal_f[DATA][15] , 
        \chan_internal_f[DATA][14] , \chan_internal_f[DATA][13] , 
        \chan_internal_f[DATA][12] , \chan_internal_f[DATA][11] , 
        \chan_internal_f[DATA][10] , \chan_internal_f[DATA][9] , 
        \chan_internal_f[DATA][8] , \chan_internal_f[DATA][7] , 
        \chan_internal_f[DATA][6] , \chan_internal_f[DATA][5] , 
        \chan_internal_f[DATA][4] , \chan_internal_f[DATA][3] , 
        \chan_internal_f[DATA][2] , \chan_internal_f[DATA][1] , 
        \chan_internal_f[DATA][0] }), .sel({sel[4:3], SYNOPSYS_UNCONNECTED__0, 
        sel[1:0]}) );
  channel_latch_1_xxxxxxxxx_14 token_latch ( .preset(n7), .left_in({
        \chan_internal_f[REQ] , \chan_internal_f[DATA][34] , 
        \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] , 
        \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] , 
        \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] , 
        \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] , 
        \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] , 
        \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] , 
        \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] , 
        \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] , 
        \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] , 
        \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] , 
        \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] , 
        \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] , 
        \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] , 
        \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] , 
        \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] , 
        \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] , 
        \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] }), .left_out(
        \chan_in_b[ACK] ), .right_out({\chan_out_f[REQ] , 
        \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , \chan_out_f[DATA][32] , 
        \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , \chan_out_f[DATA][29] , 
        \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , \chan_out_f[DATA][26] , 
        \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , \chan_out_f[DATA][23] , 
        \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , \chan_out_f[DATA][20] , 
        \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , \chan_out_f[DATA][17] , 
        \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , \chan_out_f[DATA][14] , 
        \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , \chan_out_f[DATA][11] , 
        \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , \chan_out_f[DATA][8] , 
        \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , \chan_out_f[DATA][5] , 
        \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , \chan_out_f[DATA][2] , 
        \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), .right_in(
        \chan_out_b[ACK] ), .lt_enable(lt_en) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chan_internal_f[REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(\chan_in_f[REQ] ), .Z(req_n) );
  HS65_LS_BFX9 U1 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U2 ( .A(n3), .Z(n2) );
  HS65_LS_BFX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_BFX9 U4 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U6 ( .A(req_n), .Z(n6) );
  HS65_LS_BFX9 U7 ( .A(preset), .Z(n7) );
endmodule


module hpu_comb_0_1_3 ( data_valid, data_in, preset, data_out, sel );
  input [34:0] data_in;
  output [34:0] data_out;
  output [4:0] sel;
  input data_valid, preset;
  wire   data_in_34, data_in_33, data_in_32, \data_in[31] , \data_in[30] ,
         \data_in[29] , \data_in[28] , \data_in[27] , \data_in[26] ,
         \data_in[25] , \data_in[24] , \data_in[23] , \data_in[22] ,
         \data_in[21] , \data_in[20] , \data_in[19] , \data_in[18] ,
         \data_in[17] , \data_in[16] , N23, N24, N26, N27, N28, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n15, n16, n17, n18;
  assign data_out[34] = data_in_34;
  assign data_in_34 = data_in[34];
  assign data_out[33] = data_in_33;
  assign data_in_33 = data_in[33];
  assign data_out[32] = data_in_32;
  assign data_in_32 = data_in[32];
  assign data_out[31] = \data_in[31] ;
  assign \data_in[31]  = data_in[31];
  assign data_out[30] = \data_in[30] ;
  assign \data_in[30]  = data_in[30];
  assign data_out[29] = \data_in[29] ;
  assign \data_in[29]  = data_in[29];
  assign data_out[28] = \data_in[28] ;
  assign \data_in[28]  = data_in[28];
  assign data_out[27] = \data_in[27] ;
  assign \data_in[27]  = data_in[27];
  assign data_out[26] = \data_in[26] ;
  assign \data_in[26]  = data_in[26];
  assign data_out[25] = \data_in[25] ;
  assign \data_in[25]  = data_in[25];
  assign data_out[24] = \data_in[24] ;
  assign \data_in[24]  = data_in[24];
  assign data_out[23] = \data_in[23] ;
  assign \data_in[23]  = data_in[23];
  assign data_out[22] = \data_in[22] ;
  assign \data_in[22]  = data_in[22];
  assign data_out[21] = \data_in[21] ;
  assign \data_in[21]  = data_in[21];
  assign data_out[20] = \data_in[20] ;
  assign \data_in[20]  = data_in[20];
  assign data_out[19] = \data_in[19] ;
  assign \data_in[19]  = data_in[19];
  assign data_out[18] = \data_in[18] ;
  assign \data_in[18]  = data_in[18];
  assign data_out[17] = \data_in[17] ;
  assign \data_in[17]  = data_in[17];
  assign data_out[16] = \data_in[16] ;
  assign \data_in[16]  = data_in[16];
  assign sel[1] = 1'b0;

  HS65_LS_LDHQX9 \sel_reg[4]  ( .G(N23), .D(N28), .Q(sel[4]) );
  HS65_LS_LDHQX9 \sel_reg[3]  ( .G(N23), .D(N27), .Q(sel[3]) );
  HS65_LS_LDHQX9 \sel_reg[2]  ( .G(N23), .D(N26), .Q(sel[2]) );
  HS65_LS_LDHQX9 \sel_reg[0]  ( .G(N23), .D(N24), .Q(sel[0]) );
  HS65_LS_OAI22X6 U4 ( .A(n6), .B(n18), .C(n2), .D(n7), .Z(data_out[7]) );
  HS65_LS_OAI22X6 U5 ( .A(n18), .B(n9), .C(n2), .D(n10), .Z(data_out[1]) );
  HS65_LS_OAI22X6 U6 ( .A(n18), .B(n8), .C(n2), .D(n9), .Z(data_out[3]) );
  HS65_LS_OAI22X6 U7 ( .A(n18), .B(n7), .C(n2), .D(n8), .Z(data_out[5]) );
  HS65_LS_OAI22X6 U8 ( .A(n18), .B(n5), .C(n2), .D(n6), .Z(data_out[9]) );
  HS65_LS_OAI22X6 U9 ( .A(n18), .B(n4), .C(n2), .D(n5), .Z(data_out[11]) );
  HS65_LS_OAI22X6 U10 ( .A(n18), .B(n3), .C(n2), .D(n4), .Z(data_out[13]) );
  HS65_LS_NAND3AX6 U11 ( .A(preset), .B(n17), .C(n2), .Z(n16) );
  HS65_LS_NOR3X4 U12 ( .A(n17), .B(preset), .C(n18), .Z(N28) );
  HS65_LS_IVX9 U13 ( .A(n18), .Z(n2) );
  HS65_LS_NOR3X4 U14 ( .A(n16), .B(n10), .C(n15), .Z(N27) );
  HS65_LS_NOR2AX3 U15 ( .A(n15), .B(n16), .Z(N26) );
  HS65_LS_NOR2X6 U16 ( .A(n2), .B(n3), .Z(data_out[15]) );
  HS65_LS_NAND2X14 U17 ( .A(data_in_34), .B(data_in_33), .Z(n18) );
  HS65_LS_IVX9 U18 ( .A(data_in[1]), .Z(n10) );
  HS65_LS_NAND2X7 U19 ( .A(data_in[0]), .B(n10), .Z(n17) );
  HS65_LS_NOR2X6 U20 ( .A(n10), .B(data_in[0]), .Z(n15) );
  HS65_LS_NOR2X6 U21 ( .A(data_in[1]), .B(n16), .Z(N24) );
  HS65_LS_IVX9 U22 ( .A(data_in[9]), .Z(n6) );
  HS65_LS_IVX9 U23 ( .A(data_in[3]), .Z(n9) );
  HS65_LS_IVX9 U24 ( .A(data_in[5]), .Z(n8) );
  HS65_LS_IVX9 U25 ( .A(data_in[7]), .Z(n7) );
  HS65_LS_IVX9 U26 ( .A(data_in[11]), .Z(n5) );
  HS65_LS_IVX9 U27 ( .A(data_in[13]), .Z(n4) );
  HS65_LS_IVX9 U28 ( .A(data_in[15]), .Z(n3) );
  HS65_LS_AO22X9 U29 ( .A(n2), .B(data_in[2]), .C(n18), .D(data_in[0]), .Z(
        data_out[0]) );
  HS65_LS_AO22X9 U30 ( .A(n2), .B(data_in[4]), .C(n18), .D(data_in[2]), .Z(
        data_out[2]) );
  HS65_LS_AO22X9 U31 ( .A(n2), .B(data_in[6]), .C(n18), .D(data_in[4]), .Z(
        data_out[4]) );
  HS65_LS_AO22X9 U32 ( .A(n2), .B(data_in[8]), .C(n18), .D(data_in[6]), .Z(
        data_out[6]) );
  HS65_LS_AO22X9 U33 ( .A(n2), .B(data_in[10]), .C(n18), .D(data_in[8]), .Z(
        data_out[8]) );
  HS65_LS_AO22X9 U34 ( .A(n2), .B(data_in[12]), .C(n18), .D(data_in[10]), .Z(
        data_out[10]) );
  HS65_LS_AO22X9 U35 ( .A(n2), .B(data_in[14]), .C(n18), .D(data_in[12]), .Z(
        data_out[12]) );
  HS65_LS_AND2X4 U36 ( .A(data_in[14]), .B(n18), .Z(data_out[14]) );
  HS65_LS_CB4I6X9 U37 ( .A(n2), .B(n1), .C(data_valid), .D(preset), .Z(N23) );
  HS65_LS_IVX9 U38 ( .A(data_in_34), .Z(n1) );
endmodule


module latch_controller_1_13 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_13 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_13 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n7) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_IVX9 U3 ( .A(N0), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_0_1_3 ( preset, .chan_in_f({\chan_in_f[REQ] , \chan_in_f[DATA][34] , 
        \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , 
        \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , 
        \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , 
        \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , 
        \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , 
        \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , 
        \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , 
        \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , 
        \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , 
        \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , 
        \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , 
        \chan_in_f[DATA][0] }), .chan_in_b(\chan_in_b[ACK] ), .chan_out_f({
        \chan_out_f[REQ] , \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , 
        \chan_out_f[DATA][32] , \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , 
        \chan_out_f[DATA][29] , \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , 
        \chan_out_f[DATA][26] , \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , 
        \chan_out_f[DATA][23] , \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , 
        \chan_out_f[DATA][20] , \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , 
        \chan_out_f[DATA][17] , \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , 
        \chan_out_f[DATA][14] , \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , 
        \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , 
        \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , 
        \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , 
        \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), 
    .chan_out_b(\chan_out_b[ACK] ), sel );
  output [4:0] sel;
  input preset, \chan_in_f[REQ] , \chan_in_f[DATA][34] , \chan_in_f[DATA][33] ,
         \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , \chan_in_f[DATA][30] ,
         \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , \chan_in_f[DATA][27] ,
         \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , \chan_in_f[DATA][24] ,
         \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , \chan_in_f[DATA][21] ,
         \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , \chan_in_f[DATA][18] ,
         \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , \chan_in_f[DATA][15] ,
         \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , \chan_in_f[DATA][12] ,
         \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , \chan_in_f[DATA][9] ,
         \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , \chan_in_f[DATA][6] ,
         \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , \chan_in_f[DATA][3] ,
         \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , \chan_in_f[DATA][0] ,
         \chan_out_b[ACK] ;
  output \chan_in_b[ACK] , \chan_out_f[REQ] , \chan_out_f[DATA][34] ,
         \chan_out_f[DATA][33] , \chan_out_f[DATA][32] ,
         \chan_out_f[DATA][31] , \chan_out_f[DATA][30] ,
         \chan_out_f[DATA][29] , \chan_out_f[DATA][28] ,
         \chan_out_f[DATA][27] , \chan_out_f[DATA][26] ,
         \chan_out_f[DATA][25] , \chan_out_f[DATA][24] ,
         \chan_out_f[DATA][23] , \chan_out_f[DATA][22] ,
         \chan_out_f[DATA][21] , \chan_out_f[DATA][20] ,
         \chan_out_f[DATA][19] , \chan_out_f[DATA][18] ,
         \chan_out_f[DATA][17] , \chan_out_f[DATA][16] ,
         \chan_out_f[DATA][15] , \chan_out_f[DATA][14] ,
         \chan_out_f[DATA][13] , \chan_out_f[DATA][12] ,
         \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] ,
         \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] ,
         \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] ,
         \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] ;
  wire   \chan_internal_f[REQ] , \chan_internal_f[DATA][34] ,
         \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] ,
         \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] ,
         \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] ,
         \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] ,
         \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] ,
         \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] ,
         \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] ,
         \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] ,
         \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] ,
         \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] ,
         \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] ,
         \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] ,
         \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] ,
         \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] ,
         \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] ,
         \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] ,
         \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] , req_n, lt_en,
         n1, n2, n3, n4, n5, n6, n7;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign sel[1] = 1'b0;

  hpu_comb_0_1_3 hpu_combinatorial ( .data_valid(lt_en), .data_in({
        \chan_in_f[DATA][34] , \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , 
        \chan_in_f[DATA][31] , \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , 
        \chan_in_f[DATA][28] , \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , 
        \chan_in_f[DATA][25] , \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , 
        \chan_in_f[DATA][22] , \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , 
        \chan_in_f[DATA][19] , \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , 
        \chan_in_f[DATA][16] , \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , 
        \chan_in_f[DATA][13] , \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , 
        \chan_in_f[DATA][10] , \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , 
        \chan_in_f[DATA][7] , \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , 
        \chan_in_f[DATA][4] , \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , 
        \chan_in_f[DATA][1] , \chan_in_f[DATA][0] }), .preset(n7), .data_out({
        \chan_internal_f[DATA][34] , \chan_internal_f[DATA][33] , 
        \chan_internal_f[DATA][32] , \chan_internal_f[DATA][31] , 
        \chan_internal_f[DATA][30] , \chan_internal_f[DATA][29] , 
        \chan_internal_f[DATA][28] , \chan_internal_f[DATA][27] , 
        \chan_internal_f[DATA][26] , \chan_internal_f[DATA][25] , 
        \chan_internal_f[DATA][24] , \chan_internal_f[DATA][23] , 
        \chan_internal_f[DATA][22] , \chan_internal_f[DATA][21] , 
        \chan_internal_f[DATA][20] , \chan_internal_f[DATA][19] , 
        \chan_internal_f[DATA][18] , \chan_internal_f[DATA][17] , 
        \chan_internal_f[DATA][16] , \chan_internal_f[DATA][15] , 
        \chan_internal_f[DATA][14] , \chan_internal_f[DATA][13] , 
        \chan_internal_f[DATA][12] , \chan_internal_f[DATA][11] , 
        \chan_internal_f[DATA][10] , \chan_internal_f[DATA][9] , 
        \chan_internal_f[DATA][8] , \chan_internal_f[DATA][7] , 
        \chan_internal_f[DATA][6] , \chan_internal_f[DATA][5] , 
        \chan_internal_f[DATA][4] , \chan_internal_f[DATA][3] , 
        \chan_internal_f[DATA][2] , \chan_internal_f[DATA][1] , 
        \chan_internal_f[DATA][0] }), .sel({sel[4:2], SYNOPSYS_UNCONNECTED__0, 
        sel[0]}) );
  channel_latch_1_xxxxxxxxx_13 token_latch ( .preset(n7), .left_in({
        \chan_internal_f[REQ] , \chan_internal_f[DATA][34] , 
        \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] , 
        \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] , 
        \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] , 
        \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] , 
        \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] , 
        \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] , 
        \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] , 
        \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] , 
        \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] , 
        \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] , 
        \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] , 
        \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] , 
        \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] , 
        \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] , 
        \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] , 
        \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] , 
        \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] }), .left_out(
        \chan_in_b[ACK] ), .right_out({\chan_out_f[REQ] , 
        \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , \chan_out_f[DATA][32] , 
        \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , \chan_out_f[DATA][29] , 
        \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , \chan_out_f[DATA][26] , 
        \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , \chan_out_f[DATA][23] , 
        \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , \chan_out_f[DATA][20] , 
        \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , \chan_out_f[DATA][17] , 
        \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , \chan_out_f[DATA][14] , 
        \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , \chan_out_f[DATA][11] , 
        \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , \chan_out_f[DATA][8] , 
        \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , \chan_out_f[DATA][5] , 
        \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , \chan_out_f[DATA][2] , 
        \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), .right_in(
        \chan_out_b[ACK] ), .lt_enable(lt_en) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chan_internal_f[REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(\chan_in_f[REQ] ), .Z(req_n) );
  HS65_LS_BFX9 U1 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U2 ( .A(n3), .Z(n2) );
  HS65_LS_BFX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_BFX9 U4 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U6 ( .A(req_n), .Z(n6) );
  HS65_LS_BFX9 U7 ( .A(preset), .Z(n7) );
endmodule


module hpu_comb_0_3_3 ( data_valid, data_in, preset, data_out, sel );
  input [34:0] data_in;
  output [34:0] data_out;
  output [4:0] sel;
  input data_valid, preset;
  wire   data_in_34, data_in_33, data_in_32, \data_in[31] , \data_in[30] ,
         \data_in[29] , \data_in[28] , \data_in[27] , \data_in[26] ,
         \data_in[25] , \data_in[24] , \data_in[23] , \data_in[22] ,
         \data_in[21] , \data_in[20] , \data_in[19] , \data_in[18] ,
         \data_in[17] , \data_in[16] , N25, N26, N27, N28, N30, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n15, n16, n17, n18;
  assign data_out[34] = data_in_34;
  assign data_in_34 = data_in[34];
  assign data_out[33] = data_in_33;
  assign data_in_33 = data_in[33];
  assign data_out[32] = data_in_32;
  assign data_in_32 = data_in[32];
  assign data_out[31] = \data_in[31] ;
  assign \data_in[31]  = data_in[31];
  assign data_out[30] = \data_in[30] ;
  assign \data_in[30]  = data_in[30];
  assign data_out[29] = \data_in[29] ;
  assign \data_in[29]  = data_in[29];
  assign data_out[28] = \data_in[28] ;
  assign \data_in[28]  = data_in[28];
  assign data_out[27] = \data_in[27] ;
  assign \data_in[27]  = data_in[27];
  assign data_out[26] = \data_in[26] ;
  assign \data_in[26]  = data_in[26];
  assign data_out[25] = \data_in[25] ;
  assign \data_in[25]  = data_in[25];
  assign data_out[24] = \data_in[24] ;
  assign \data_in[24]  = data_in[24];
  assign data_out[23] = \data_in[23] ;
  assign \data_in[23]  = data_in[23];
  assign data_out[22] = \data_in[22] ;
  assign \data_in[22]  = data_in[22];
  assign data_out[21] = \data_in[21] ;
  assign \data_in[21]  = data_in[21];
  assign data_out[20] = \data_in[20] ;
  assign \data_in[20]  = data_in[20];
  assign data_out[19] = \data_in[19] ;
  assign \data_in[19]  = data_in[19];
  assign data_out[18] = \data_in[18] ;
  assign \data_in[18]  = data_in[18];
  assign data_out[17] = \data_in[17] ;
  assign \data_in[17]  = data_in[17];
  assign data_out[16] = \data_in[16] ;
  assign \data_in[16]  = data_in[16];
  assign sel[3] = 1'b0;

  HS65_LS_LDHQX9 \sel_reg[4]  ( .G(N25), .D(N30), .Q(sel[4]) );
  HS65_LS_LDHQX9 \sel_reg[2]  ( .G(N25), .D(N28), .Q(sel[2]) );
  HS65_LS_LDHQX9 \sel_reg[1]  ( .G(N25), .D(N27), .Q(sel[1]) );
  HS65_LS_LDHQX9 \sel_reg[0]  ( .G(N25), .D(N26), .Q(sel[0]) );
  HS65_LS_OAI22X6 U4 ( .A(n18), .B(n9), .C(n2), .D(n10), .Z(data_out[0]) );
  HS65_LS_OAI22X6 U5 ( .A(n18), .B(n8), .C(n2), .D(n9), .Z(data_out[2]) );
  HS65_LS_OAI22X6 U6 ( .A(n18), .B(n7), .C(n2), .D(n8), .Z(data_out[4]) );
  HS65_LS_OAI22X6 U7 ( .A(n18), .B(n6), .C(n2), .D(n7), .Z(data_out[6]) );
  HS65_LS_OAI22X6 U8 ( .A(n18), .B(n5), .C(n2), .D(n6), .Z(data_out[8]) );
  HS65_LS_OAI22X6 U9 ( .A(n18), .B(n4), .C(n2), .D(n5), .Z(data_out[10]) );
  HS65_LS_OAI22X6 U10 ( .A(n18), .B(n3), .C(n2), .D(n4), .Z(data_out[12]) );
  HS65_LS_NAND3AX6 U11 ( .A(preset), .B(n17), .C(n2), .Z(n16) );
  HS65_LS_NOR3X4 U12 ( .A(n17), .B(preset), .C(n18), .Z(N30) );
  HS65_LS_IVX9 U13 ( .A(n18), .Z(n2) );
  HS65_LS_NOR2X6 U14 ( .A(n10), .B(n16), .Z(N27) );
  HS65_LS_NOR2AX3 U15 ( .A(n15), .B(n16), .Z(N26) );
  HS65_LS_NOR2X6 U16 ( .A(n2), .B(n3), .Z(data_out[14]) );
  HS65_LS_NAND2X14 U17 ( .A(data_in_34), .B(data_in_33), .Z(n18) );
  HS65_LS_NOR3X4 U18 ( .A(n16), .B(data_in[0]), .C(n15), .Z(N28) );
  HS65_LS_NAND2X7 U19 ( .A(data_in[0]), .B(data_in[1]), .Z(n17) );
  HS65_LS_NOR2X6 U20 ( .A(data_in[1]), .B(data_in[0]), .Z(n15) );
  HS65_LS_IVX9 U21 ( .A(data_in[0]), .Z(n10) );
  HS65_LS_IVX9 U22 ( .A(data_in[2]), .Z(n9) );
  HS65_LS_IVX9 U23 ( .A(data_in[4]), .Z(n8) );
  HS65_LS_IVX9 U24 ( .A(data_in[6]), .Z(n7) );
  HS65_LS_IVX9 U25 ( .A(data_in[8]), .Z(n6) );
  HS65_LS_IVX9 U26 ( .A(data_in[10]), .Z(n5) );
  HS65_LS_IVX9 U27 ( .A(data_in[12]), .Z(n4) );
  HS65_LS_IVX9 U28 ( .A(data_in[14]), .Z(n3) );
  HS65_LS_AO22X9 U29 ( .A(n2), .B(data_in[3]), .C(n18), .D(data_in[1]), .Z(
        data_out[1]) );
  HS65_LS_AO22X9 U30 ( .A(n2), .B(data_in[5]), .C(n18), .D(data_in[3]), .Z(
        data_out[3]) );
  HS65_LS_AO22X9 U31 ( .A(n2), .B(data_in[7]), .C(n18), .D(data_in[5]), .Z(
        data_out[5]) );
  HS65_LS_AO22X9 U32 ( .A(data_in[9]), .B(n2), .C(n18), .D(data_in[7]), .Z(
        data_out[7]) );
  HS65_LS_AO22X9 U33 ( .A(n2), .B(data_in[11]), .C(n18), .D(data_in[9]), .Z(
        data_out[9]) );
  HS65_LS_AO22X9 U34 ( .A(n2), .B(data_in[13]), .C(n18), .D(data_in[11]), .Z(
        data_out[11]) );
  HS65_LS_AO22X9 U35 ( .A(n2), .B(data_in[15]), .C(n18), .D(data_in[13]), .Z(
        data_out[13]) );
  HS65_LS_AND2X4 U36 ( .A(data_in[15]), .B(n18), .Z(data_out[15]) );
  HS65_LS_CB4I6X9 U37 ( .A(n2), .B(n1), .C(data_valid), .D(preset), .Z(N25) );
  HS65_LS_IVX9 U38 ( .A(data_in_34), .Z(n1) );
endmodule


module latch_controller_1_12 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_12 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_12 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n7) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_IVX9 U3 ( .A(N0), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_0_3_3 ( preset, .chan_in_f({\chan_in_f[REQ] , \chan_in_f[DATA][34] , 
        \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , 
        \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , 
        \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , 
        \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , 
        \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , 
        \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , 
        \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , 
        \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , 
        \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , 
        \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , 
        \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , 
        \chan_in_f[DATA][0] }), .chan_in_b(\chan_in_b[ACK] ), .chan_out_f({
        \chan_out_f[REQ] , \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , 
        \chan_out_f[DATA][32] , \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , 
        \chan_out_f[DATA][29] , \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , 
        \chan_out_f[DATA][26] , \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , 
        \chan_out_f[DATA][23] , \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , 
        \chan_out_f[DATA][20] , \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , 
        \chan_out_f[DATA][17] , \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , 
        \chan_out_f[DATA][14] , \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , 
        \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , 
        \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , 
        \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , 
        \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), 
    .chan_out_b(\chan_out_b[ACK] ), sel );
  output [4:0] sel;
  input preset, \chan_in_f[REQ] , \chan_in_f[DATA][34] , \chan_in_f[DATA][33] ,
         \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , \chan_in_f[DATA][30] ,
         \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , \chan_in_f[DATA][27] ,
         \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , \chan_in_f[DATA][24] ,
         \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , \chan_in_f[DATA][21] ,
         \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , \chan_in_f[DATA][18] ,
         \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , \chan_in_f[DATA][15] ,
         \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , \chan_in_f[DATA][12] ,
         \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , \chan_in_f[DATA][9] ,
         \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , \chan_in_f[DATA][6] ,
         \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , \chan_in_f[DATA][3] ,
         \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , \chan_in_f[DATA][0] ,
         \chan_out_b[ACK] ;
  output \chan_in_b[ACK] , \chan_out_f[REQ] , \chan_out_f[DATA][34] ,
         \chan_out_f[DATA][33] , \chan_out_f[DATA][32] ,
         \chan_out_f[DATA][31] , \chan_out_f[DATA][30] ,
         \chan_out_f[DATA][29] , \chan_out_f[DATA][28] ,
         \chan_out_f[DATA][27] , \chan_out_f[DATA][26] ,
         \chan_out_f[DATA][25] , \chan_out_f[DATA][24] ,
         \chan_out_f[DATA][23] , \chan_out_f[DATA][22] ,
         \chan_out_f[DATA][21] , \chan_out_f[DATA][20] ,
         \chan_out_f[DATA][19] , \chan_out_f[DATA][18] ,
         \chan_out_f[DATA][17] , \chan_out_f[DATA][16] ,
         \chan_out_f[DATA][15] , \chan_out_f[DATA][14] ,
         \chan_out_f[DATA][13] , \chan_out_f[DATA][12] ,
         \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] ,
         \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] ,
         \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] ,
         \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] ;
  wire   \chan_internal_f[REQ] , \chan_internal_f[DATA][34] ,
         \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] ,
         \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] ,
         \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] ,
         \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] ,
         \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] ,
         \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] ,
         \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] ,
         \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] ,
         \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] ,
         \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] ,
         \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] ,
         \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] ,
         \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] ,
         \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] ,
         \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] ,
         \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] ,
         \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] , req_n, lt_en,
         n1, n2, n3, n4, n5, n6, n7;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign sel[3] = 1'b0;

  hpu_comb_0_3_3 hpu_combinatorial ( .data_valid(lt_en), .data_in({
        \chan_in_f[DATA][34] , \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , 
        \chan_in_f[DATA][31] , \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , 
        \chan_in_f[DATA][28] , \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , 
        \chan_in_f[DATA][25] , \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , 
        \chan_in_f[DATA][22] , \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , 
        \chan_in_f[DATA][19] , \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , 
        \chan_in_f[DATA][16] , \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , 
        \chan_in_f[DATA][13] , \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , 
        \chan_in_f[DATA][10] , \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , 
        \chan_in_f[DATA][7] , \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , 
        \chan_in_f[DATA][4] , \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , 
        \chan_in_f[DATA][1] , \chan_in_f[DATA][0] }), .preset(n7), .data_out({
        \chan_internal_f[DATA][34] , \chan_internal_f[DATA][33] , 
        \chan_internal_f[DATA][32] , \chan_internal_f[DATA][31] , 
        \chan_internal_f[DATA][30] , \chan_internal_f[DATA][29] , 
        \chan_internal_f[DATA][28] , \chan_internal_f[DATA][27] , 
        \chan_internal_f[DATA][26] , \chan_internal_f[DATA][25] , 
        \chan_internal_f[DATA][24] , \chan_internal_f[DATA][23] , 
        \chan_internal_f[DATA][22] , \chan_internal_f[DATA][21] , 
        \chan_internal_f[DATA][20] , \chan_internal_f[DATA][19] , 
        \chan_internal_f[DATA][18] , \chan_internal_f[DATA][17] , 
        \chan_internal_f[DATA][16] , \chan_internal_f[DATA][15] , 
        \chan_internal_f[DATA][14] , \chan_internal_f[DATA][13] , 
        \chan_internal_f[DATA][12] , \chan_internal_f[DATA][11] , 
        \chan_internal_f[DATA][10] , \chan_internal_f[DATA][9] , 
        \chan_internal_f[DATA][8] , \chan_internal_f[DATA][7] , 
        \chan_internal_f[DATA][6] , \chan_internal_f[DATA][5] , 
        \chan_internal_f[DATA][4] , \chan_internal_f[DATA][3] , 
        \chan_internal_f[DATA][2] , \chan_internal_f[DATA][1] , 
        \chan_internal_f[DATA][0] }), .sel({sel[4], SYNOPSYS_UNCONNECTED__0, 
        sel[2:0]}) );
  channel_latch_1_xxxxxxxxx_12 token_latch ( .preset(n7), .left_in({
        \chan_internal_f[REQ] , \chan_internal_f[DATA][34] , 
        \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] , 
        \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] , 
        \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] , 
        \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] , 
        \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] , 
        \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] , 
        \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] , 
        \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] , 
        \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] , 
        \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] , 
        \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] , 
        \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] , 
        \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] , 
        \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] , 
        \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] , 
        \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] , 
        \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] }), .left_out(
        \chan_in_b[ACK] ), .right_out({\chan_out_f[REQ] , 
        \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , \chan_out_f[DATA][32] , 
        \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , \chan_out_f[DATA][29] , 
        \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , \chan_out_f[DATA][26] , 
        \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , \chan_out_f[DATA][23] , 
        \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , \chan_out_f[DATA][20] , 
        \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , \chan_out_f[DATA][17] , 
        \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , \chan_out_f[DATA][14] , 
        \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , \chan_out_f[DATA][11] , 
        \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , \chan_out_f[DATA][8] , 
        \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , \chan_out_f[DATA][5] , 
        \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , \chan_out_f[DATA][2] , 
        \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), .right_in(
        \chan_out_b[ACK] ), .lt_enable(lt_en) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chan_internal_f[REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(\chan_in_f[REQ] ), .Z(req_n) );
  HS65_LS_BFX9 U1 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U2 ( .A(n3), .Z(n2) );
  HS65_LS_BFX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_BFX9 U4 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U6 ( .A(req_n), .Z(n6) );
  HS65_LS_BFX9 U7 ( .A(preset), .Z(n7) );
endmodule


module hpu_comb_1_x_3 ( data_valid, data_in, preset, data_out, sel );
  input [34:0] data_in;
  output [34:0] data_out;
  output [4:0] sel;
  input data_valid, preset;
  wire   data_in_34, data_in_33, data_in_32, \data_in[31] , \data_in[30] ,
         \data_in[29] , \data_in[28] , \data_in[27] , \data_in[26] ,
         \data_in[25] , \data_in[24] , \data_in[23] , \data_in[22] ,
         \data_in[21] , \data_in[20] , \data_in[19] , \data_in[18] ,
         \data_in[17] , \data_in[16] , N19, N20, N21, N22, N23, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n22,
         n23, n24;
  assign data_out[34] = data_in_34;
  assign data_in_34 = data_in[34];
  assign data_out[33] = data_in_33;
  assign data_in_33 = data_in[33];
  assign data_out[32] = data_in_32;
  assign data_in_32 = data_in[32];
  assign data_out[31] = \data_in[31] ;
  assign \data_in[31]  = data_in[31];
  assign data_out[30] = \data_in[30] ;
  assign \data_in[30]  = data_in[30];
  assign data_out[29] = \data_in[29] ;
  assign \data_in[29]  = data_in[29];
  assign data_out[28] = \data_in[28] ;
  assign \data_in[28]  = data_in[28];
  assign data_out[27] = \data_in[27] ;
  assign \data_in[27]  = data_in[27];
  assign data_out[26] = \data_in[26] ;
  assign \data_in[26]  = data_in[26];
  assign data_out[25] = \data_in[25] ;
  assign \data_in[25]  = data_in[25];
  assign data_out[24] = \data_in[24] ;
  assign \data_in[24]  = data_in[24];
  assign data_out[23] = \data_in[23] ;
  assign \data_in[23]  = data_in[23];
  assign data_out[22] = \data_in[22] ;
  assign \data_in[22]  = data_in[22];
  assign data_out[21] = \data_in[21] ;
  assign \data_in[21]  = data_in[21];
  assign data_out[20] = \data_in[20] ;
  assign \data_in[20]  = data_in[20];
  assign data_out[19] = \data_in[19] ;
  assign \data_in[19]  = data_in[19];
  assign data_out[18] = \data_in[18] ;
  assign \data_in[18]  = data_in[18];
  assign data_out[17] = \data_in[17] ;
  assign \data_in[17]  = data_in[17];
  assign data_out[16] = \data_in[16] ;
  assign \data_in[16]  = data_in[16];
  assign sel[4] = 1'b0;

  HS65_LS_LDHQX9 \sel_reg[3]  ( .G(N19), .D(N23), .Q(sel[3]) );
  HS65_LS_LDHQX9 \sel_reg[2]  ( .G(N19), .D(N22), .Q(sel[2]) );
  HS65_LS_LDHQX9 \sel_reg[1]  ( .G(N19), .D(N21), .Q(sel[1]) );
  HS65_LS_LDHQX9 \sel_reg[0]  ( .G(N19), .D(N20), .Q(sel[0]) );
  HS65_LS_NAND3AX3 U4 ( .A(preset), .B(n22), .C(n2), .Z(n23) );
  HS65_LS_NOR3X3 U5 ( .A(n23), .B(n17), .C(n18), .Z(N23) );
  HS65_LS_NAND2X21 U6 ( .A(data_in_34), .B(data_in_33), .Z(n24) );
  HS65_LS_NOR2X5 U7 ( .A(data_in[1]), .B(n23), .Z(N21) );
  HS65_LS_IVX7 U8 ( .A(data_in_34), .Z(n1) );
  HS65_LS_OAI22X6 U9 ( .A(n9), .B(n24), .C(n2), .D(n11), .Z(data_out[7]) );
  HS65_LS_OAI22X6 U10 ( .A(n24), .B(n16), .C(n2), .D(n18), .Z(data_out[0]) );
  HS65_LS_OAI22X6 U11 ( .A(n24), .B(n15), .C(n2), .D(n17), .Z(data_out[1]) );
  HS65_LS_OAI22X6 U12 ( .A(n24), .B(n14), .C(n2), .D(n16), .Z(data_out[2]) );
  HS65_LS_OAI22X6 U13 ( .A(n24), .B(n13), .C(n2), .D(n15), .Z(data_out[3]) );
  HS65_LS_OAI22X6 U14 ( .A(n24), .B(n12), .C(n2), .D(n14), .Z(data_out[4]) );
  HS65_LS_OAI22X6 U15 ( .A(n24), .B(n11), .C(n2), .D(n13), .Z(data_out[5]) );
  HS65_LS_OAI22X6 U16 ( .A(n24), .B(n10), .C(n2), .D(n12), .Z(data_out[6]) );
  HS65_LS_OAI22X6 U17 ( .A(n24), .B(n8), .C(n2), .D(n10), .Z(data_out[8]) );
  HS65_LS_OAI22X6 U18 ( .A(n24), .B(n7), .C(n2), .D(n9), .Z(data_out[9]) );
  HS65_LS_OAI22X6 U19 ( .A(n24), .B(n6), .C(n2), .D(n8), .Z(data_out[10]) );
  HS65_LS_OAI22X6 U20 ( .A(n24), .B(n5), .C(n2), .D(n7), .Z(data_out[11]) );
  HS65_LS_OAI22X6 U21 ( .A(n24), .B(n4), .C(n2), .D(n6), .Z(data_out[12]) );
  HS65_LS_OAI22X6 U22 ( .A(n24), .B(n3), .C(n2), .D(n5), .Z(data_out[13]) );
  HS65_LS_IVX9 U23 ( .A(n24), .Z(n2) );
  HS65_LS_NOR3X4 U24 ( .A(n22), .B(preset), .C(n24), .Z(N20) );
  HS65_LS_NAND2X7 U25 ( .A(n17), .B(n18), .Z(n22) );
  HS65_LS_NOR2X6 U26 ( .A(n2), .B(n4), .Z(data_out[14]) );
  HS65_LS_NOR2X6 U27 ( .A(n2), .B(n3), .Z(data_out[15]) );
  HS65_LS_IVX9 U28 ( .A(data_in[1]), .Z(n17) );
  HS65_LS_IVX9 U29 ( .A(data_in[0]), .Z(n18) );
  HS65_LS_NOR2X6 U30 ( .A(data_in[0]), .B(n23), .Z(N22) );
  HS65_LS_IVX9 U31 ( .A(data_in[9]), .Z(n9) );
  HS65_LS_IVX9 U32 ( .A(data_in[2]), .Z(n16) );
  HS65_LS_IVX9 U33 ( .A(data_in[3]), .Z(n15) );
  HS65_LS_IVX9 U34 ( .A(data_in[4]), .Z(n14) );
  HS65_LS_IVX9 U35 ( .A(data_in[5]), .Z(n13) );
  HS65_LS_IVX9 U36 ( .A(data_in[7]), .Z(n11) );
  HS65_LS_IVX9 U37 ( .A(data_in[10]), .Z(n8) );
  HS65_LS_IVX9 U38 ( .A(data_in[12]), .Z(n6) );
  HS65_LS_IVX9 U39 ( .A(data_in[13]), .Z(n5) );
  HS65_LS_IVX9 U40 ( .A(data_in[14]), .Z(n4) );
  HS65_LS_IVX9 U41 ( .A(data_in[15]), .Z(n3) );
  HS65_LS_IVX9 U42 ( .A(data_in[6]), .Z(n12) );
  HS65_LS_IVX9 U43 ( .A(data_in[8]), .Z(n10) );
  HS65_LS_IVX9 U44 ( .A(data_in[11]), .Z(n7) );
  HS65_LS_CB4I6X9 U45 ( .A(n2), .B(n1), .C(data_valid), .D(preset), .Z(N19) );
endmodule


module latch_controller_1_11 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_11 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_11 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n7) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_IVX9 U3 ( .A(N0), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_1_x_3 ( preset, .chan_in_f({\chan_in_f[REQ] , \chan_in_f[DATA][34] , 
        \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , 
        \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , 
        \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , 
        \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , 
        \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , 
        \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , 
        \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , 
        \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , 
        \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , 
        \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , 
        \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , 
        \chan_in_f[DATA][0] }), .chan_in_b(\chan_in_b[ACK] ), .chan_out_f({
        \chan_out_f[REQ] , \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , 
        \chan_out_f[DATA][32] , \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , 
        \chan_out_f[DATA][29] , \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , 
        \chan_out_f[DATA][26] , \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , 
        \chan_out_f[DATA][23] , \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , 
        \chan_out_f[DATA][20] , \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , 
        \chan_out_f[DATA][17] , \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , 
        \chan_out_f[DATA][14] , \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , 
        \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , 
        \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , 
        \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , 
        \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), 
    .chan_out_b(\chan_out_b[ACK] ), sel );
  output [4:0] sel;
  input preset, \chan_in_f[REQ] , \chan_in_f[DATA][34] , \chan_in_f[DATA][33] ,
         \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , \chan_in_f[DATA][30] ,
         \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , \chan_in_f[DATA][27] ,
         \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , \chan_in_f[DATA][24] ,
         \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , \chan_in_f[DATA][21] ,
         \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , \chan_in_f[DATA][18] ,
         \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , \chan_in_f[DATA][15] ,
         \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , \chan_in_f[DATA][12] ,
         \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , \chan_in_f[DATA][9] ,
         \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , \chan_in_f[DATA][6] ,
         \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , \chan_in_f[DATA][3] ,
         \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , \chan_in_f[DATA][0] ,
         \chan_out_b[ACK] ;
  output \chan_in_b[ACK] , \chan_out_f[REQ] , \chan_out_f[DATA][34] ,
         \chan_out_f[DATA][33] , \chan_out_f[DATA][32] ,
         \chan_out_f[DATA][31] , \chan_out_f[DATA][30] ,
         \chan_out_f[DATA][29] , \chan_out_f[DATA][28] ,
         \chan_out_f[DATA][27] , \chan_out_f[DATA][26] ,
         \chan_out_f[DATA][25] , \chan_out_f[DATA][24] ,
         \chan_out_f[DATA][23] , \chan_out_f[DATA][22] ,
         \chan_out_f[DATA][21] , \chan_out_f[DATA][20] ,
         \chan_out_f[DATA][19] , \chan_out_f[DATA][18] ,
         \chan_out_f[DATA][17] , \chan_out_f[DATA][16] ,
         \chan_out_f[DATA][15] , \chan_out_f[DATA][14] ,
         \chan_out_f[DATA][13] , \chan_out_f[DATA][12] ,
         \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] ,
         \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] ,
         \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] ,
         \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] ;
  wire   \chan_internal_f[REQ] , \chan_internal_f[DATA][34] ,
         \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] ,
         \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] ,
         \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] ,
         \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] ,
         \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] ,
         \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] ,
         \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] ,
         \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] ,
         \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] ,
         \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] ,
         \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] ,
         \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] ,
         \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] ,
         \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] ,
         \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] ,
         \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] ,
         \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] , req_n, lt_en,
         n1, n2, n3, n4, n5, n6, n7;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign sel[4] = 1'b0;

  hpu_comb_1_x_3 hpu_combinatorial ( .data_valid(lt_en), .data_in({
        \chan_in_f[DATA][34] , \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , 
        \chan_in_f[DATA][31] , \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , 
        \chan_in_f[DATA][28] , \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , 
        \chan_in_f[DATA][25] , \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , 
        \chan_in_f[DATA][22] , \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , 
        \chan_in_f[DATA][19] , \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , 
        \chan_in_f[DATA][16] , \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , 
        \chan_in_f[DATA][13] , \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , 
        \chan_in_f[DATA][10] , \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , 
        \chan_in_f[DATA][7] , \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , 
        \chan_in_f[DATA][4] , \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , 
        \chan_in_f[DATA][1] , \chan_in_f[DATA][0] }), .preset(n7), .data_out({
        \chan_internal_f[DATA][34] , \chan_internal_f[DATA][33] , 
        \chan_internal_f[DATA][32] , \chan_internal_f[DATA][31] , 
        \chan_internal_f[DATA][30] , \chan_internal_f[DATA][29] , 
        \chan_internal_f[DATA][28] , \chan_internal_f[DATA][27] , 
        \chan_internal_f[DATA][26] , \chan_internal_f[DATA][25] , 
        \chan_internal_f[DATA][24] , \chan_internal_f[DATA][23] , 
        \chan_internal_f[DATA][22] , \chan_internal_f[DATA][21] , 
        \chan_internal_f[DATA][20] , \chan_internal_f[DATA][19] , 
        \chan_internal_f[DATA][18] , \chan_internal_f[DATA][17] , 
        \chan_internal_f[DATA][16] , \chan_internal_f[DATA][15] , 
        \chan_internal_f[DATA][14] , \chan_internal_f[DATA][13] , 
        \chan_internal_f[DATA][12] , \chan_internal_f[DATA][11] , 
        \chan_internal_f[DATA][10] , \chan_internal_f[DATA][9] , 
        \chan_internal_f[DATA][8] , \chan_internal_f[DATA][7] , 
        \chan_internal_f[DATA][6] , \chan_internal_f[DATA][5] , 
        \chan_internal_f[DATA][4] , \chan_internal_f[DATA][3] , 
        \chan_internal_f[DATA][2] , \chan_internal_f[DATA][1] , 
        \chan_internal_f[DATA][0] }), .sel({SYNOPSYS_UNCONNECTED__0, sel[3:0]}) );
  channel_latch_1_xxxxxxxxx_11 token_latch ( .preset(n7), .left_in({
        \chan_internal_f[REQ] , \chan_internal_f[DATA][34] , 
        \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] , 
        \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] , 
        \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] , 
        \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] , 
        \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] , 
        \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] , 
        \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] , 
        \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] , 
        \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] , 
        \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] , 
        \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] , 
        \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] , 
        \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] , 
        \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] , 
        \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] , 
        \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] , 
        \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] }), .left_out(
        \chan_in_b[ACK] ), .right_out({\chan_out_f[REQ] , 
        \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , \chan_out_f[DATA][32] , 
        \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , \chan_out_f[DATA][29] , 
        \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , \chan_out_f[DATA][26] , 
        \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , \chan_out_f[DATA][23] , 
        \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , \chan_out_f[DATA][20] , 
        \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , \chan_out_f[DATA][17] , 
        \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , \chan_out_f[DATA][14] , 
        \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , \chan_out_f[DATA][11] , 
        \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , \chan_out_f[DATA][8] , 
        \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , \chan_out_f[DATA][5] , 
        \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , \chan_out_f[DATA][2] , 
        \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), .right_in(
        \chan_out_b[ACK] ), .lt_enable(lt_en) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chan_internal_f[REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(\chan_in_f[REQ] ), .Z(req_n) );
  HS65_LS_BFX9 U1 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U2 ( .A(n3), .Z(n2) );
  HS65_LS_BFX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_BFX9 U4 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U6 ( .A(req_n), .Z(n6) );
  HS65_LS_BFX9 U7 ( .A(preset), .Z(n7) );
endmodule


module sr_latch_1_6 ( s, r, q, qn );
  input s, r;
  output q, qn;
  wire   N3, n1;

  HS65_LS_AND2X4 C9 ( .A(n1), .B(N3), .Z(qn) );
  HS65_LH_NOR2X3 U1 ( .A(r), .B(qn), .Z(q) );
  HS65_LS_IVX9 U2 ( .A(q), .Z(N3) );
  HS65_LS_IVX9 U3 ( .A(s), .Z(n1) );
endmodule


module c_gate_generic_1_5_6 ( preset, \input , \output  );
  input [4:0] \input ;
  input preset;
  output \output ;
  wire   set, reset, n1, n4, n5;

  sr_latch_1_6 latch ( .s(set), .r(reset), .q(\output ) );
  HS65_LS_NOR3X4 U3 ( .A(\input [3]), .B(preset), .C(\input [4]), .Z(n4) );
  HS65_LS_NOR4ABX2 U4 ( .A(n1), .B(n4), .C(\input [2]), .D(\input [1]), .Z(
        reset) );
  HS65_LS_AO31X9 U5 ( .A(n5), .B(\input [3]), .C(\input [4]), .D(preset), .Z(
        set) );
  HS65_LS_IVX9 U6 ( .A(\input [0]), .Z(n1) );
  HS65_LS_AND3X9 U7 ( .A(\input [1]), .B(\input [0]), .C(\input [2]), .Z(n5)
         );
endmodule


module sr_latch_1_5 ( s, r, q, qn );
  input s, r;
  output q, qn;
  wire   N3, n1;

  HS65_LS_AND2X4 C9 ( .A(n1), .B(N3), .Z(qn) );
  HS65_LS_IVX9 U1 ( .A(q), .Z(N3) );
  HS65_LS_IVX9 U2 ( .A(s), .Z(n1) );
  HS65_LS_NOR2X6 U3 ( .A(r), .B(qn), .Z(q) );
endmodule


module c_gate_generic_1_5_5 ( preset, \input , \output  );
  input [4:0] \input ;
  input preset;
  output \output ;
  wire   set, reset, n1, n4, n5;

  sr_latch_1_5 latch ( .s(set), .r(reset), .q(\output ) );
  HS65_LS_NOR3X4 U3 ( .A(\input [3]), .B(preset), .C(\input [4]), .Z(n4) );
  HS65_LS_NOR4ABX2 U4 ( .A(n1), .B(n4), .C(\input [2]), .D(\input [1]), .Z(
        reset) );
  HS65_LS_AO31X9 U5 ( .A(n5), .B(\input [3]), .C(\input [4]), .D(preset), .Z(
        set) );
  HS65_LS_IVX9 U6 ( .A(\input [0]), .Z(n1) );
  HS65_LS_AND3X9 U7 ( .A(\input [1]), .B(\input [0]), .C(\input [2]), .Z(n5)
         );
endmodule


module crossbar_3 ( preset, .switch_sel({\switch_sel[4][4] , 
        \switch_sel[4][3] , \switch_sel[4][2] , \switch_sel[4][1] , 
        \switch_sel[4][0] , \switch_sel[3][4] , \switch_sel[3][3] , 
        \switch_sel[3][2] , \switch_sel[3][1] , \switch_sel[3][0] , 
        \switch_sel[2][4] , \switch_sel[2][3] , \switch_sel[2][2] , 
        \switch_sel[2][1] , \switch_sel[2][0] , \switch_sel[1][4] , 
        \switch_sel[1][3] , \switch_sel[1][2] , \switch_sel[1][1] , 
        \switch_sel[1][0] , \switch_sel[0][4] , \switch_sel[0][3] , 
        \switch_sel[0][2] , \switch_sel[0][1] , \switch_sel[0][0] }), 
    .chs_in_f({\chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] , 
        \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] , 
        \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] , 
        \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] , 
        \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] , 
        \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] , 
        \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] , 
        \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] , 
        \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] , 
        \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] , 
        \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] , 
        \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] , 
        \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] , 
        \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] , \chs_in_f[4][DATA][7] , 
        \chs_in_f[4][DATA][6] , \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] , 
        \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] , \chs_in_f[4][DATA][1] , 
        \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] , \chs_in_f[3][DATA][34] , 
        \chs_in_f[3][DATA][33] , \chs_in_f[3][DATA][32] , 
        \chs_in_f[3][DATA][31] , \chs_in_f[3][DATA][30] , 
        \chs_in_f[3][DATA][29] , \chs_in_f[3][DATA][28] , 
        \chs_in_f[3][DATA][27] , \chs_in_f[3][DATA][26] , 
        \chs_in_f[3][DATA][25] , \chs_in_f[3][DATA][24] , 
        \chs_in_f[3][DATA][23] , \chs_in_f[3][DATA][22] , 
        \chs_in_f[3][DATA][21] , \chs_in_f[3][DATA][20] , 
        \chs_in_f[3][DATA][19] , \chs_in_f[3][DATA][18] , 
        \chs_in_f[3][DATA][17] , \chs_in_f[3][DATA][16] , 
        \chs_in_f[3][DATA][15] , \chs_in_f[3][DATA][14] , 
        \chs_in_f[3][DATA][13] , \chs_in_f[3][DATA][12] , 
        \chs_in_f[3][DATA][11] , \chs_in_f[3][DATA][10] , 
        \chs_in_f[3][DATA][9] , \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] , 
        \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] , \chs_in_f[3][DATA][4] , 
        \chs_in_f[3][DATA][3] , \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] , 
        \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] , 
        \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] , 
        \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] , 
        \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] , 
        \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] , 
        \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] , 
        \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] , 
        \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] , 
        \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] , 
        \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] , 
        \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] , 
        \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] , 
        \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] , 
        \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] , \chs_in_f[2][DATA][7] , 
        \chs_in_f[2][DATA][6] , \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] , 
        \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] , \chs_in_f[2][DATA][1] , 
        \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] , \chs_in_f[1][DATA][34] , 
        \chs_in_f[1][DATA][33] , \chs_in_f[1][DATA][32] , 
        \chs_in_f[1][DATA][31] , \chs_in_f[1][DATA][30] , 
        \chs_in_f[1][DATA][29] , \chs_in_f[1][DATA][28] , 
        \chs_in_f[1][DATA][27] , \chs_in_f[1][DATA][26] , 
        \chs_in_f[1][DATA][25] , \chs_in_f[1][DATA][24] , 
        \chs_in_f[1][DATA][23] , \chs_in_f[1][DATA][22] , 
        \chs_in_f[1][DATA][21] , \chs_in_f[1][DATA][20] , 
        \chs_in_f[1][DATA][19] , \chs_in_f[1][DATA][18] , 
        \chs_in_f[1][DATA][17] , \chs_in_f[1][DATA][16] , 
        \chs_in_f[1][DATA][15] , \chs_in_f[1][DATA][14] , 
        \chs_in_f[1][DATA][13] , \chs_in_f[1][DATA][12] , 
        \chs_in_f[1][DATA][11] , \chs_in_f[1][DATA][10] , 
        \chs_in_f[1][DATA][9] , \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] , 
        \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] , \chs_in_f[1][DATA][4] , 
        \chs_in_f[1][DATA][3] , \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] , 
        \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] , 
        \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] , 
        \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] , 
        \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] , 
        \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] , 
        \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] , 
        \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] , 
        \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] , 
        \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] , 
        \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] , 
        \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] , 
        \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] , 
        \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] , 
        \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] , \chs_in_f[0][DATA][7] , 
        \chs_in_f[0][DATA][6] , \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] , 
        \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] , \chs_in_f[0][DATA][1] , 
        \chs_in_f[0][DATA][0] }), .chs_in_b({\chs_in_b[4][ACK] , 
        \chs_in_b[3][ACK] , \chs_in_b[2][ACK] , \chs_in_b[1][ACK] , 
        \chs_in_b[0][ACK] }), .chs_out_f({\chs_out_f[4][REQ] , 
        \chs_out_f[4][DATA][34] , \chs_out_f[4][DATA][33] , 
        \chs_out_f[4][DATA][32] , \chs_out_f[4][DATA][31] , 
        \chs_out_f[4][DATA][30] , \chs_out_f[4][DATA][29] , 
        \chs_out_f[4][DATA][28] , \chs_out_f[4][DATA][27] , 
        \chs_out_f[4][DATA][26] , \chs_out_f[4][DATA][25] , 
        \chs_out_f[4][DATA][24] , \chs_out_f[4][DATA][23] , 
        \chs_out_f[4][DATA][22] , \chs_out_f[4][DATA][21] , 
        \chs_out_f[4][DATA][20] , \chs_out_f[4][DATA][19] , 
        \chs_out_f[4][DATA][18] , \chs_out_f[4][DATA][17] , 
        \chs_out_f[4][DATA][16] , \chs_out_f[4][DATA][15] , 
        \chs_out_f[4][DATA][14] , \chs_out_f[4][DATA][13] , 
        \chs_out_f[4][DATA][12] , \chs_out_f[4][DATA][11] , 
        \chs_out_f[4][DATA][10] , \chs_out_f[4][DATA][9] , 
        \chs_out_f[4][DATA][8] , \chs_out_f[4][DATA][7] , 
        \chs_out_f[4][DATA][6] , \chs_out_f[4][DATA][5] , 
        \chs_out_f[4][DATA][4] , \chs_out_f[4][DATA][3] , 
        \chs_out_f[4][DATA][2] , \chs_out_f[4][DATA][1] , 
        \chs_out_f[4][DATA][0] , \chs_out_f[3][REQ] , \chs_out_f[3][DATA][34] , 
        \chs_out_f[3][DATA][33] , \chs_out_f[3][DATA][32] , 
        \chs_out_f[3][DATA][31] , \chs_out_f[3][DATA][30] , 
        \chs_out_f[3][DATA][29] , \chs_out_f[3][DATA][28] , 
        \chs_out_f[3][DATA][27] , \chs_out_f[3][DATA][26] , 
        \chs_out_f[3][DATA][25] , \chs_out_f[3][DATA][24] , 
        \chs_out_f[3][DATA][23] , \chs_out_f[3][DATA][22] , 
        \chs_out_f[3][DATA][21] , \chs_out_f[3][DATA][20] , 
        \chs_out_f[3][DATA][19] , \chs_out_f[3][DATA][18] , 
        \chs_out_f[3][DATA][17] , \chs_out_f[3][DATA][16] , 
        \chs_out_f[3][DATA][15] , \chs_out_f[3][DATA][14] , 
        \chs_out_f[3][DATA][13] , \chs_out_f[3][DATA][12] , 
        \chs_out_f[3][DATA][11] , \chs_out_f[3][DATA][10] , 
        \chs_out_f[3][DATA][9] , \chs_out_f[3][DATA][8] , 
        \chs_out_f[3][DATA][7] , \chs_out_f[3][DATA][6] , 
        \chs_out_f[3][DATA][5] , \chs_out_f[3][DATA][4] , 
        \chs_out_f[3][DATA][3] , \chs_out_f[3][DATA][2] , 
        \chs_out_f[3][DATA][1] , \chs_out_f[3][DATA][0] , \chs_out_f[2][REQ] , 
        \chs_out_f[2][DATA][34] , \chs_out_f[2][DATA][33] , 
        \chs_out_f[2][DATA][32] , \chs_out_f[2][DATA][31] , 
        \chs_out_f[2][DATA][30] , \chs_out_f[2][DATA][29] , 
        \chs_out_f[2][DATA][28] , \chs_out_f[2][DATA][27] , 
        \chs_out_f[2][DATA][26] , \chs_out_f[2][DATA][25] , 
        \chs_out_f[2][DATA][24] , \chs_out_f[2][DATA][23] , 
        \chs_out_f[2][DATA][22] , \chs_out_f[2][DATA][21] , 
        \chs_out_f[2][DATA][20] , \chs_out_f[2][DATA][19] , 
        \chs_out_f[2][DATA][18] , \chs_out_f[2][DATA][17] , 
        \chs_out_f[2][DATA][16] , \chs_out_f[2][DATA][15] , 
        \chs_out_f[2][DATA][14] , \chs_out_f[2][DATA][13] , 
        \chs_out_f[2][DATA][12] , \chs_out_f[2][DATA][11] , 
        \chs_out_f[2][DATA][10] , \chs_out_f[2][DATA][9] , 
        \chs_out_f[2][DATA][8] , \chs_out_f[2][DATA][7] , 
        \chs_out_f[2][DATA][6] , \chs_out_f[2][DATA][5] , 
        \chs_out_f[2][DATA][4] , \chs_out_f[2][DATA][3] , 
        \chs_out_f[2][DATA][2] , \chs_out_f[2][DATA][1] , 
        \chs_out_f[2][DATA][0] , \chs_out_f[1][REQ] , \chs_out_f[1][DATA][34] , 
        \chs_out_f[1][DATA][33] , \chs_out_f[1][DATA][32] , 
        \chs_out_f[1][DATA][31] , \chs_out_f[1][DATA][30] , 
        \chs_out_f[1][DATA][29] , \chs_out_f[1][DATA][28] , 
        \chs_out_f[1][DATA][27] , \chs_out_f[1][DATA][26] , 
        \chs_out_f[1][DATA][25] , \chs_out_f[1][DATA][24] , 
        \chs_out_f[1][DATA][23] , \chs_out_f[1][DATA][22] , 
        \chs_out_f[1][DATA][21] , \chs_out_f[1][DATA][20] , 
        \chs_out_f[1][DATA][19] , \chs_out_f[1][DATA][18] , 
        \chs_out_f[1][DATA][17] , \chs_out_f[1][DATA][16] , 
        \chs_out_f[1][DATA][15] , \chs_out_f[1][DATA][14] , 
        \chs_out_f[1][DATA][13] , \chs_out_f[1][DATA][12] , 
        \chs_out_f[1][DATA][11] , \chs_out_f[1][DATA][10] , 
        \chs_out_f[1][DATA][9] , \chs_out_f[1][DATA][8] , 
        \chs_out_f[1][DATA][7] , \chs_out_f[1][DATA][6] , 
        \chs_out_f[1][DATA][5] , \chs_out_f[1][DATA][4] , 
        \chs_out_f[1][DATA][3] , \chs_out_f[1][DATA][2] , 
        \chs_out_f[1][DATA][1] , \chs_out_f[1][DATA][0] , \chs_out_f[0][REQ] , 
        \chs_out_f[0][DATA][34] , \chs_out_f[0][DATA][33] , 
        \chs_out_f[0][DATA][32] , \chs_out_f[0][DATA][31] , 
        \chs_out_f[0][DATA][30] , \chs_out_f[0][DATA][29] , 
        \chs_out_f[0][DATA][28] , \chs_out_f[0][DATA][27] , 
        \chs_out_f[0][DATA][26] , \chs_out_f[0][DATA][25] , 
        \chs_out_f[0][DATA][24] , \chs_out_f[0][DATA][23] , 
        \chs_out_f[0][DATA][22] , \chs_out_f[0][DATA][21] , 
        \chs_out_f[0][DATA][20] , \chs_out_f[0][DATA][19] , 
        \chs_out_f[0][DATA][18] , \chs_out_f[0][DATA][17] , 
        \chs_out_f[0][DATA][16] , \chs_out_f[0][DATA][15] , 
        \chs_out_f[0][DATA][14] , \chs_out_f[0][DATA][13] , 
        \chs_out_f[0][DATA][12] , \chs_out_f[0][DATA][11] , 
        \chs_out_f[0][DATA][10] , \chs_out_f[0][DATA][9] , 
        \chs_out_f[0][DATA][8] , \chs_out_f[0][DATA][7] , 
        \chs_out_f[0][DATA][6] , \chs_out_f[0][DATA][5] , 
        \chs_out_f[0][DATA][4] , \chs_out_f[0][DATA][3] , 
        \chs_out_f[0][DATA][2] , \chs_out_f[0][DATA][1] , 
        \chs_out_f[0][DATA][0] }), .chs_out_b({\chs_out_b[4][ACK] , 
        \chs_out_b[3][ACK] , \chs_out_b[2][ACK] , \chs_out_b[1][ACK] , 
        \chs_out_b[0][ACK] }) );
  input preset, \switch_sel[4][4] , \switch_sel[4][3] , \switch_sel[4][2] ,
         \switch_sel[4][1] , \switch_sel[4][0] , \switch_sel[3][4] ,
         \switch_sel[3][3] , \switch_sel[3][2] , \switch_sel[3][1] ,
         \switch_sel[3][0] , \switch_sel[2][4] , \switch_sel[2][3] ,
         \switch_sel[2][2] , \switch_sel[2][1] , \switch_sel[2][0] ,
         \switch_sel[1][4] , \switch_sel[1][3] , \switch_sel[1][2] ,
         \switch_sel[1][1] , \switch_sel[1][0] , \switch_sel[0][4] ,
         \switch_sel[0][3] , \switch_sel[0][2] , \switch_sel[0][1] ,
         \switch_sel[0][0] , \chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] ,
         \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] ,
         \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] ,
         \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] ,
         \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] ,
         \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] ,
         \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] ,
         \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] ,
         \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] ,
         \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] ,
         \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] ,
         \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] ,
         \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] ,
         \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] ,
         \chs_in_f[4][DATA][7] , \chs_in_f[4][DATA][6] ,
         \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] ,
         \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] ,
         \chs_in_f[4][DATA][1] , \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] ,
         \chs_in_f[3][DATA][34] , \chs_in_f[3][DATA][33] ,
         \chs_in_f[3][DATA][32] , \chs_in_f[3][DATA][31] ,
         \chs_in_f[3][DATA][30] , \chs_in_f[3][DATA][29] ,
         \chs_in_f[3][DATA][28] , \chs_in_f[3][DATA][27] ,
         \chs_in_f[3][DATA][26] , \chs_in_f[3][DATA][25] ,
         \chs_in_f[3][DATA][24] , \chs_in_f[3][DATA][23] ,
         \chs_in_f[3][DATA][22] , \chs_in_f[3][DATA][21] ,
         \chs_in_f[3][DATA][20] , \chs_in_f[3][DATA][19] ,
         \chs_in_f[3][DATA][18] , \chs_in_f[3][DATA][17] ,
         \chs_in_f[3][DATA][16] , \chs_in_f[3][DATA][15] ,
         \chs_in_f[3][DATA][14] , \chs_in_f[3][DATA][13] ,
         \chs_in_f[3][DATA][12] , \chs_in_f[3][DATA][11] ,
         \chs_in_f[3][DATA][10] , \chs_in_f[3][DATA][9] ,
         \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] ,
         \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] ,
         \chs_in_f[3][DATA][4] , \chs_in_f[3][DATA][3] ,
         \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] ,
         \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] ,
         \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] ,
         \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] ,
         \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] ,
         \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] ,
         \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] ,
         \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] ,
         \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] ,
         \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] ,
         \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] ,
         \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] ,
         \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] ,
         \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] ,
         \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] ,
         \chs_in_f[2][DATA][7] , \chs_in_f[2][DATA][6] ,
         \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] ,
         \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] ,
         \chs_in_f[2][DATA][1] , \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] ,
         \chs_in_f[1][DATA][34] , \chs_in_f[1][DATA][33] ,
         \chs_in_f[1][DATA][32] , \chs_in_f[1][DATA][31] ,
         \chs_in_f[1][DATA][30] , \chs_in_f[1][DATA][29] ,
         \chs_in_f[1][DATA][28] , \chs_in_f[1][DATA][27] ,
         \chs_in_f[1][DATA][26] , \chs_in_f[1][DATA][25] ,
         \chs_in_f[1][DATA][24] , \chs_in_f[1][DATA][23] ,
         \chs_in_f[1][DATA][22] , \chs_in_f[1][DATA][21] ,
         \chs_in_f[1][DATA][20] , \chs_in_f[1][DATA][19] ,
         \chs_in_f[1][DATA][18] , \chs_in_f[1][DATA][17] ,
         \chs_in_f[1][DATA][16] , \chs_in_f[1][DATA][15] ,
         \chs_in_f[1][DATA][14] , \chs_in_f[1][DATA][13] ,
         \chs_in_f[1][DATA][12] , \chs_in_f[1][DATA][11] ,
         \chs_in_f[1][DATA][10] , \chs_in_f[1][DATA][9] ,
         \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] ,
         \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] ,
         \chs_in_f[1][DATA][4] , \chs_in_f[1][DATA][3] ,
         \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] ,
         \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] ,
         \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] ,
         \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] ,
         \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] ,
         \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] ,
         \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] ,
         \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] ,
         \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] ,
         \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] ,
         \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] ,
         \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] ,
         \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] ,
         \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] ,
         \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] ,
         \chs_in_f[0][DATA][7] , \chs_in_f[0][DATA][6] ,
         \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] ,
         \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] ,
         \chs_in_f[0][DATA][1] , \chs_in_f[0][DATA][0] , \chs_out_b[4][ACK] ,
         \chs_out_b[3][ACK] , \chs_out_b[2][ACK] , \chs_out_b[1][ACK] ,
         \chs_out_b[0][ACK] ;
  output \chs_in_b[4][ACK] , \chs_in_b[3][ACK] , \chs_in_b[2][ACK] ,
         \chs_in_b[1][ACK] , \chs_in_b[0][ACK] , \chs_out_f[4][REQ] ,
         \chs_out_f[4][DATA][34] , \chs_out_f[4][DATA][33] ,
         \chs_out_f[4][DATA][32] , \chs_out_f[4][DATA][31] ,
         \chs_out_f[4][DATA][30] , \chs_out_f[4][DATA][29] ,
         \chs_out_f[4][DATA][28] , \chs_out_f[4][DATA][27] ,
         \chs_out_f[4][DATA][26] , \chs_out_f[4][DATA][25] ,
         \chs_out_f[4][DATA][24] , \chs_out_f[4][DATA][23] ,
         \chs_out_f[4][DATA][22] , \chs_out_f[4][DATA][21] ,
         \chs_out_f[4][DATA][20] , \chs_out_f[4][DATA][19] ,
         \chs_out_f[4][DATA][18] , \chs_out_f[4][DATA][17] ,
         \chs_out_f[4][DATA][16] , \chs_out_f[4][DATA][15] ,
         \chs_out_f[4][DATA][14] , \chs_out_f[4][DATA][13] ,
         \chs_out_f[4][DATA][12] , \chs_out_f[4][DATA][11] ,
         \chs_out_f[4][DATA][10] , \chs_out_f[4][DATA][9] ,
         \chs_out_f[4][DATA][8] , \chs_out_f[4][DATA][7] ,
         \chs_out_f[4][DATA][6] , \chs_out_f[4][DATA][5] ,
         \chs_out_f[4][DATA][4] , \chs_out_f[4][DATA][3] ,
         \chs_out_f[4][DATA][2] , \chs_out_f[4][DATA][1] ,
         \chs_out_f[4][DATA][0] , \chs_out_f[3][REQ] ,
         \chs_out_f[3][DATA][34] , \chs_out_f[3][DATA][33] ,
         \chs_out_f[3][DATA][32] , \chs_out_f[3][DATA][31] ,
         \chs_out_f[3][DATA][30] , \chs_out_f[3][DATA][29] ,
         \chs_out_f[3][DATA][28] , \chs_out_f[3][DATA][27] ,
         \chs_out_f[3][DATA][26] , \chs_out_f[3][DATA][25] ,
         \chs_out_f[3][DATA][24] , \chs_out_f[3][DATA][23] ,
         \chs_out_f[3][DATA][22] , \chs_out_f[3][DATA][21] ,
         \chs_out_f[3][DATA][20] , \chs_out_f[3][DATA][19] ,
         \chs_out_f[3][DATA][18] , \chs_out_f[3][DATA][17] ,
         \chs_out_f[3][DATA][16] , \chs_out_f[3][DATA][15] ,
         \chs_out_f[3][DATA][14] , \chs_out_f[3][DATA][13] ,
         \chs_out_f[3][DATA][12] , \chs_out_f[3][DATA][11] ,
         \chs_out_f[3][DATA][10] , \chs_out_f[3][DATA][9] ,
         \chs_out_f[3][DATA][8] , \chs_out_f[3][DATA][7] ,
         \chs_out_f[3][DATA][6] , \chs_out_f[3][DATA][5] ,
         \chs_out_f[3][DATA][4] , \chs_out_f[3][DATA][3] ,
         \chs_out_f[3][DATA][2] , \chs_out_f[3][DATA][1] ,
         \chs_out_f[3][DATA][0] , \chs_out_f[2][REQ] ,
         \chs_out_f[2][DATA][34] , \chs_out_f[2][DATA][33] ,
         \chs_out_f[2][DATA][32] , \chs_out_f[2][DATA][31] ,
         \chs_out_f[2][DATA][30] , \chs_out_f[2][DATA][29] ,
         \chs_out_f[2][DATA][28] , \chs_out_f[2][DATA][27] ,
         \chs_out_f[2][DATA][26] , \chs_out_f[2][DATA][25] ,
         \chs_out_f[2][DATA][24] , \chs_out_f[2][DATA][23] ,
         \chs_out_f[2][DATA][22] , \chs_out_f[2][DATA][21] ,
         \chs_out_f[2][DATA][20] , \chs_out_f[2][DATA][19] ,
         \chs_out_f[2][DATA][18] , \chs_out_f[2][DATA][17] ,
         \chs_out_f[2][DATA][16] , \chs_out_f[2][DATA][15] ,
         \chs_out_f[2][DATA][14] , \chs_out_f[2][DATA][13] ,
         \chs_out_f[2][DATA][12] , \chs_out_f[2][DATA][11] ,
         \chs_out_f[2][DATA][10] , \chs_out_f[2][DATA][9] ,
         \chs_out_f[2][DATA][8] , \chs_out_f[2][DATA][7] ,
         \chs_out_f[2][DATA][6] , \chs_out_f[2][DATA][5] ,
         \chs_out_f[2][DATA][4] , \chs_out_f[2][DATA][3] ,
         \chs_out_f[2][DATA][2] , \chs_out_f[2][DATA][1] ,
         \chs_out_f[2][DATA][0] , \chs_out_f[1][REQ] ,
         \chs_out_f[1][DATA][34] , \chs_out_f[1][DATA][33] ,
         \chs_out_f[1][DATA][32] , \chs_out_f[1][DATA][31] ,
         \chs_out_f[1][DATA][30] , \chs_out_f[1][DATA][29] ,
         \chs_out_f[1][DATA][28] , \chs_out_f[1][DATA][27] ,
         \chs_out_f[1][DATA][26] , \chs_out_f[1][DATA][25] ,
         \chs_out_f[1][DATA][24] , \chs_out_f[1][DATA][23] ,
         \chs_out_f[1][DATA][22] , \chs_out_f[1][DATA][21] ,
         \chs_out_f[1][DATA][20] , \chs_out_f[1][DATA][19] ,
         \chs_out_f[1][DATA][18] , \chs_out_f[1][DATA][17] ,
         \chs_out_f[1][DATA][16] , \chs_out_f[1][DATA][15] ,
         \chs_out_f[1][DATA][14] , \chs_out_f[1][DATA][13] ,
         \chs_out_f[1][DATA][12] , \chs_out_f[1][DATA][11] ,
         \chs_out_f[1][DATA][10] , \chs_out_f[1][DATA][9] ,
         \chs_out_f[1][DATA][8] , \chs_out_f[1][DATA][7] ,
         \chs_out_f[1][DATA][6] , \chs_out_f[1][DATA][5] ,
         \chs_out_f[1][DATA][4] , \chs_out_f[1][DATA][3] ,
         \chs_out_f[1][DATA][2] , \chs_out_f[1][DATA][1] ,
         \chs_out_f[1][DATA][0] , \chs_out_f[0][REQ] ,
         \chs_out_f[0][DATA][34] , \chs_out_f[0][DATA][33] ,
         \chs_out_f[0][DATA][32] , \chs_out_f[0][DATA][31] ,
         \chs_out_f[0][DATA][30] , \chs_out_f[0][DATA][29] ,
         \chs_out_f[0][DATA][28] , \chs_out_f[0][DATA][27] ,
         \chs_out_f[0][DATA][26] , \chs_out_f[0][DATA][25] ,
         \chs_out_f[0][DATA][24] , \chs_out_f[0][DATA][23] ,
         \chs_out_f[0][DATA][22] , \chs_out_f[0][DATA][21] ,
         \chs_out_f[0][DATA][20] , \chs_out_f[0][DATA][19] ,
         \chs_out_f[0][DATA][18] , \chs_out_f[0][DATA][17] ,
         \chs_out_f[0][DATA][16] , \chs_out_f[0][DATA][15] ,
         \chs_out_f[0][DATA][14] , \chs_out_f[0][DATA][13] ,
         \chs_out_f[0][DATA][12] , \chs_out_f[0][DATA][11] ,
         \chs_out_f[0][DATA][10] , \chs_out_f[0][DATA][9] ,
         \chs_out_f[0][DATA][8] , \chs_out_f[0][DATA][7] ,
         \chs_out_f[0][DATA][6] , \chs_out_f[0][DATA][5] ,
         \chs_out_f[0][DATA][4] , \chs_out_f[0][DATA][3] ,
         \chs_out_f[0][DATA][2] , \chs_out_f[0][DATA][1] ,
         \chs_out_f[0][DATA][0] ;
  wire   \chs_in_b[4][ACK] , \chs_out_f[4][REQ] , synced_req, del, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510;
  assign \chs_in_b[0][ACK]  = \chs_in_b[4][ACK] ;
  assign \chs_in_b[1][ACK]  = \chs_in_b[4][ACK] ;
  assign \chs_in_b[2][ACK]  = \chs_in_b[4][ACK] ;
  assign \chs_in_b[3][ACK]  = \chs_in_b[4][ACK] ;
  assign \chs_out_f[0][REQ]  = \chs_out_f[4][REQ] ;
  assign \chs_out_f[1][REQ]  = \chs_out_f[4][REQ] ;
  assign \chs_out_f[2][REQ]  = \chs_out_f[4][REQ] ;
  assign \chs_out_f[3][REQ]  = \chs_out_f[4][REQ] ;

  c_gate_generic_1_5_6 c_sync_req ( .preset(preset), .\input ({
        \chs_in_f[4][REQ] , \chs_in_f[3][REQ] , \chs_in_f[2][REQ] , 
        \chs_in_f[1][REQ] , \chs_in_f[0][REQ] }), .\output (synced_req) );
  c_gate_generic_1_5_5 c_sync_ack ( .preset(preset), .\input ({
        \chs_out_b[4][ACK] , \chs_out_b[3][ACK] , \chs_out_b[2][ACK] , 
        \chs_out_b[1][ACK] , \chs_out_b[0][ACK] }), .\output (
        \chs_in_b[4][ACK] ) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chs_out_f[4][REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(synced_req), .Z(del) );
  HS65_LS_IVX9 U2 ( .A(\switch_sel[3][4] ), .Z(n261) );
  HS65_LS_IVX9 U3 ( .A(\switch_sel[3][2] ), .Z(n262) );
  HS65_LS_IVX9 U4 ( .A(\switch_sel[3][1] ), .Z(n263) );
  HS65_LS_IVX9 U5 ( .A(\switch_sel[3][0] ), .Z(n264) );
  HS65_LS_BFX9 U6 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U7 ( .A(del), .Z(n2) );
  HS65_LS_BFX9 U8 ( .A(n258), .Z(n11) );
  HS65_LS_BFX7 U9 ( .A(n257), .Z(n8) );
  HS65_LS_BFX7 U10 ( .A(n256), .Z(n5) );
  HS65_LS_BFX9 U11 ( .A(\switch_sel[0][4] ), .Z(n45) );
  HS65_LS_BFX9 U12 ( .A(\switch_sel[1][4] ), .Z(n61) );
  HS65_LS_BFX9 U13 ( .A(\switch_sel[0][3] ), .Z(n41) );
  HS65_LS_BFX9 U14 ( .A(\switch_sel[1][3] ), .Z(n57) );
  HS65_LS_BFX9 U15 ( .A(\switch_sel[1][2] ), .Z(n53) );
  HS65_LS_BFX9 U16 ( .A(\switch_sel[0][1] ), .Z(n33) );
  HS65_LS_BFX9 U17 ( .A(\switch_sel[1][0] ), .Z(n49) );
  HS65_LS_BFX9 U18 ( .A(n261), .Z(n18) );
  HS65_LS_BFX9 U19 ( .A(n261), .Z(n19) );
  HS65_LS_BFX9 U20 ( .A(n61), .Z(n62) );
  HS65_LS_BFX9 U21 ( .A(n61), .Z(n63) );
  HS65_LS_BFX9 U22 ( .A(n77), .Z(n78) );
  HS65_LS_BFX9 U23 ( .A(n77), .Z(n79) );
  HS65_LS_BFX9 U24 ( .A(n45), .Z(n46) );
  HS65_LS_BFX9 U25 ( .A(n45), .Z(n47) );
  HS65_LS_BFX9 U26 ( .A(n262), .Z(n21) );
  HS65_LS_BFX9 U27 ( .A(n262), .Z(n22) );
  HS65_LS_BFX9 U28 ( .A(n263), .Z(n24) );
  HS65_LS_BFX9 U29 ( .A(n263), .Z(n25) );
  HS65_LS_BFX9 U30 ( .A(n264), .Z(n27) );
  HS65_LS_BFX9 U31 ( .A(n264), .Z(n28) );
  HS65_LS_BFX9 U32 ( .A(n57), .Z(n58) );
  HS65_LS_BFX9 U33 ( .A(n57), .Z(n59) );
  HS65_LS_BFX9 U34 ( .A(n53), .Z(n54) );
  HS65_LS_BFX9 U35 ( .A(n53), .Z(n55) );
  HS65_LS_BFX9 U36 ( .A(n49), .Z(n50) );
  HS65_LS_BFX9 U37 ( .A(n49), .Z(n51) );
  HS65_LS_BFX9 U38 ( .A(n73), .Z(n74) );
  HS65_LS_BFX9 U39 ( .A(n73), .Z(n75) );
  HS65_LS_BFX9 U40 ( .A(n69), .Z(n70) );
  HS65_LS_BFX9 U41 ( .A(n69), .Z(n71) );
  HS65_LS_BFX9 U42 ( .A(n65), .Z(n66) );
  HS65_LS_BFX9 U43 ( .A(n65), .Z(n67) );
  HS65_LS_BFX9 U44 ( .A(n261), .Z(n20) );
  HS65_LS_BFX9 U45 ( .A(n41), .Z(n42) );
  HS65_LS_BFX9 U46 ( .A(n41), .Z(n43) );
  HS65_LS_BFX9 U47 ( .A(n37), .Z(n38) );
  HS65_LS_BFX9 U48 ( .A(n37), .Z(n39) );
  HS65_LS_BFX9 U49 ( .A(n33), .Z(n34) );
  HS65_LS_BFX9 U50 ( .A(n33), .Z(n35) );
  HS65_LS_BFX9 U51 ( .A(n45), .Z(n48) );
  HS65_LS_BFX9 U52 ( .A(n256), .Z(n3) );
  HS65_LS_BFX9 U53 ( .A(n256), .Z(n4) );
  HS65_LS_BFX9 U54 ( .A(n257), .Z(n6) );
  HS65_LS_BFX9 U55 ( .A(n257), .Z(n7) );
  HS65_LS_BFX9 U56 ( .A(n258), .Z(n9) );
  HS65_LS_BFX9 U57 ( .A(n258), .Z(n10) );
  HS65_LS_BFX9 U58 ( .A(n259), .Z(n12) );
  HS65_LS_BFX9 U59 ( .A(n259), .Z(n13) );
  HS65_LS_BFX9 U60 ( .A(n57), .Z(n60) );
  HS65_LS_BFX9 U61 ( .A(n53), .Z(n56) );
  HS65_LS_BFX9 U62 ( .A(n49), .Z(n52) );
  HS65_LS_BFX9 U63 ( .A(n73), .Z(n76) );
  HS65_LS_BFX9 U64 ( .A(n69), .Z(n72) );
  HS65_LS_BFX9 U65 ( .A(n65), .Z(n68) );
  HS65_LS_BFX9 U66 ( .A(n41), .Z(n44) );
  HS65_LS_BFX9 U67 ( .A(n37), .Z(n40) );
  HS65_LS_BFX9 U68 ( .A(n33), .Z(n36) );
  HS65_LS_BFX9 U69 ( .A(n259), .Z(n14) );
  HS65_LS_BFX9 U70 ( .A(n262), .Z(n23) );
  HS65_LS_BFX9 U71 ( .A(n263), .Z(n26) );
  HS65_LS_BFX9 U72 ( .A(n264), .Z(n29) );
  HS65_LS_BFX9 U73 ( .A(n61), .Z(n64) );
  HS65_LS_BFX9 U74 ( .A(n77), .Z(n80) );
  HS65_LS_BFX9 U75 ( .A(n260), .Z(n15) );
  HS65_LS_BFX9 U76 ( .A(n260), .Z(n16) );
  HS65_LS_BFX9 U77 ( .A(n265), .Z(n30) );
  HS65_LS_BFX9 U78 ( .A(n265), .Z(n31) );
  HS65_LS_BFX9 U79 ( .A(n260), .Z(n17) );
  HS65_LS_BFX9 U80 ( .A(n265), .Z(n32) );
  HS65_LS_IVX9 U81 ( .A(\switch_sel[4][3] ), .Z(n256) );
  HS65_LS_IVX9 U82 ( .A(\switch_sel[4][2] ), .Z(n257) );
  HS65_LS_IVX9 U83 ( .A(\switch_sel[4][1] ), .Z(n258) );
  HS65_LS_IVX9 U84 ( .A(\switch_sel[4][0] ), .Z(n259) );
  HS65_LS_AOI222X2 U85 ( .A(\chs_in_f[2][DATA][34] ), .B(n78), .C(
        \chs_in_f[0][DATA][34] ), .D(n48), .E(\chs_in_f[1][DATA][34] ), .F(n62), .Z(n503) );
  HS65_LS_OAI212X5 U86 ( .A(n291), .B(n20), .C(n326), .D(n17), .E(n510), .Z(
        \chs_out_f[4][DATA][9] ) );
  HS65_LS_AOI222X2 U87 ( .A(n78), .B(\chs_in_f[2][DATA][9] ), .C(n48), .D(
        \chs_in_f[0][DATA][9] ), .E(n62), .F(\chs_in_f[1][DATA][9] ), .Z(n510)
         );
  HS65_LS_AOI222X2 U88 ( .A(n76), .B(\chs_in_f[2][DATA][34] ), .C(n44), .D(
        \chs_in_f[0][DATA][34] ), .E(n60), .F(\chs_in_f[1][DATA][34] ), .Z(
        n468) );
  HS65_LS_AOI222X2 U89 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][34] ), 
        .C(n40), .D(\chs_in_f[0][DATA][34] ), .E(n56), .F(
        \chs_in_f[1][DATA][34] ), .Z(n433) );
  HS65_LS_AOI222X2 U90 ( .A(n72), .B(\chs_in_f[2][DATA][34] ), .C(n36), .D(
        \chs_in_f[0][DATA][34] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][34] ), .Z(n398) );
  HS65_LS_AOI222X2 U91 ( .A(n68), .B(\chs_in_f[2][DATA][34] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][34] ), .E(n52), .F(
        \chs_in_f[1][DATA][34] ), .Z(n363) );
  HS65_LS_IVX9 U92 ( .A(\chs_in_f[3][DATA][9] ), .Z(n291) );
  HS65_LS_IVX9 U93 ( .A(\chs_in_f[3][DATA][34] ), .Z(n266) );
  HS65_LS_IVX9 U94 ( .A(\chs_in_f[3][DATA][0] ), .Z(n300) );
  HS65_LS_IVX9 U95 ( .A(\chs_in_f[3][DATA][1] ), .Z(n299) );
  HS65_LS_IVX9 U96 ( .A(\chs_in_f[3][DATA][2] ), .Z(n298) );
  HS65_LS_IVX9 U97 ( .A(\chs_in_f[3][DATA][3] ), .Z(n297) );
  HS65_LS_IVX9 U98 ( .A(\chs_in_f[3][DATA][4] ), .Z(n296) );
  HS65_LS_IVX9 U99 ( .A(\chs_in_f[3][DATA][5] ), .Z(n295) );
  HS65_LS_IVX9 U100 ( .A(\chs_in_f[3][DATA][6] ), .Z(n294) );
  HS65_LS_IVX9 U101 ( .A(\chs_in_f[3][DATA][7] ), .Z(n293) );
  HS65_LS_IVX9 U102 ( .A(\chs_in_f[3][DATA][8] ), .Z(n292) );
  HS65_LS_IVX9 U103 ( .A(\chs_in_f[3][DATA][10] ), .Z(n290) );
  HS65_LS_IVX9 U104 ( .A(\chs_in_f[3][DATA][11] ), .Z(n289) );
  HS65_LS_IVX9 U105 ( .A(\chs_in_f[3][DATA][12] ), .Z(n288) );
  HS65_LS_IVX9 U106 ( .A(\chs_in_f[3][DATA][13] ), .Z(n287) );
  HS65_LS_IVX9 U107 ( .A(\chs_in_f[3][DATA][14] ), .Z(n286) );
  HS65_LS_IVX9 U108 ( .A(\chs_in_f[3][DATA][15] ), .Z(n285) );
  HS65_LS_IVX9 U109 ( .A(\chs_in_f[3][DATA][16] ), .Z(n284) );
  HS65_LS_IVX9 U110 ( .A(\chs_in_f[3][DATA][17] ), .Z(n283) );
  HS65_LS_IVX9 U111 ( .A(\chs_in_f[3][DATA][18] ), .Z(n282) );
  HS65_LS_IVX9 U112 ( .A(\chs_in_f[3][DATA][19] ), .Z(n281) );
  HS65_LS_IVX9 U113 ( .A(\chs_in_f[3][DATA][20] ), .Z(n280) );
  HS65_LS_IVX9 U114 ( .A(\chs_in_f[3][DATA][21] ), .Z(n279) );
  HS65_LS_IVX9 U115 ( .A(\chs_in_f[3][DATA][22] ), .Z(n278) );
  HS65_LS_IVX9 U116 ( .A(\chs_in_f[3][DATA][23] ), .Z(n277) );
  HS65_LS_IVX9 U117 ( .A(\chs_in_f[3][DATA][24] ), .Z(n276) );
  HS65_LS_IVX9 U118 ( .A(\chs_in_f[3][DATA][25] ), .Z(n275) );
  HS65_LS_IVX9 U119 ( .A(\chs_in_f[3][DATA][26] ), .Z(n274) );
  HS65_LS_IVX9 U120 ( .A(\chs_in_f[3][DATA][27] ), .Z(n273) );
  HS65_LS_IVX9 U121 ( .A(\chs_in_f[3][DATA][28] ), .Z(n272) );
  HS65_LS_IVX9 U122 ( .A(\chs_in_f[3][DATA][29] ), .Z(n271) );
  HS65_LS_IVX9 U123 ( .A(\chs_in_f[3][DATA][30] ), .Z(n270) );
  HS65_LS_IVX9 U124 ( .A(\chs_in_f[3][DATA][31] ), .Z(n269) );
  HS65_LS_IVX9 U125 ( .A(\chs_in_f[3][DATA][32] ), .Z(n268) );
  HS65_LS_IVX9 U126 ( .A(\chs_in_f[3][DATA][33] ), .Z(n267) );
  HS65_LS_IVX9 U127 ( .A(\chs_in_f[4][DATA][9] ), .Z(n326) );
  HS65_LS_IVX9 U128 ( .A(\chs_in_f[4][DATA][34] ), .Z(n301) );
  HS65_LS_IVX9 U129 ( .A(\chs_in_f[4][DATA][0] ), .Z(n335) );
  HS65_LS_IVX9 U130 ( .A(\chs_in_f[4][DATA][1] ), .Z(n334) );
  HS65_LS_IVX9 U131 ( .A(\chs_in_f[4][DATA][2] ), .Z(n333) );
  HS65_LS_IVX9 U132 ( .A(\chs_in_f[4][DATA][3] ), .Z(n332) );
  HS65_LS_IVX9 U133 ( .A(\chs_in_f[4][DATA][4] ), .Z(n331) );
  HS65_LS_IVX9 U134 ( .A(\chs_in_f[4][DATA][5] ), .Z(n330) );
  HS65_LS_IVX9 U135 ( .A(\chs_in_f[4][DATA][6] ), .Z(n329) );
  HS65_LS_IVX9 U136 ( .A(\chs_in_f[4][DATA][7] ), .Z(n328) );
  HS65_LS_IVX9 U137 ( .A(\chs_in_f[4][DATA][8] ), .Z(n327) );
  HS65_LS_IVX9 U138 ( .A(\chs_in_f[4][DATA][10] ), .Z(n325) );
  HS65_LS_IVX9 U139 ( .A(\chs_in_f[4][DATA][11] ), .Z(n324) );
  HS65_LS_IVX9 U140 ( .A(\chs_in_f[4][DATA][12] ), .Z(n323) );
  HS65_LS_IVX9 U141 ( .A(\chs_in_f[4][DATA][13] ), .Z(n322) );
  HS65_LS_IVX9 U142 ( .A(\chs_in_f[4][DATA][14] ), .Z(n321) );
  HS65_LS_IVX9 U143 ( .A(\chs_in_f[4][DATA][15] ), .Z(n320) );
  HS65_LS_IVX9 U144 ( .A(\chs_in_f[4][DATA][33] ), .Z(n302) );
  HS65_LS_IVX9 U145 ( .A(\chs_in_f[4][DATA][16] ), .Z(n319) );
  HS65_LS_IVX9 U146 ( .A(\chs_in_f[4][DATA][17] ), .Z(n318) );
  HS65_LS_IVX9 U147 ( .A(\chs_in_f[4][DATA][18] ), .Z(n317) );
  HS65_LS_IVX9 U148 ( .A(\chs_in_f[4][DATA][19] ), .Z(n316) );
  HS65_LS_IVX9 U149 ( .A(\chs_in_f[4][DATA][20] ), .Z(n315) );
  HS65_LS_IVX9 U150 ( .A(\chs_in_f[4][DATA][21] ), .Z(n314) );
  HS65_LS_IVX9 U151 ( .A(\chs_in_f[4][DATA][22] ), .Z(n313) );
  HS65_LS_IVX9 U152 ( .A(\chs_in_f[4][DATA][23] ), .Z(n312) );
  HS65_LS_IVX9 U153 ( .A(\chs_in_f[4][DATA][24] ), .Z(n311) );
  HS65_LS_IVX9 U154 ( .A(\chs_in_f[4][DATA][25] ), .Z(n310) );
  HS65_LS_IVX9 U155 ( .A(\chs_in_f[4][DATA][26] ), .Z(n309) );
  HS65_LS_IVX9 U156 ( .A(\chs_in_f[4][DATA][27] ), .Z(n308) );
  HS65_LS_IVX9 U157 ( .A(\chs_in_f[4][DATA][28] ), .Z(n307) );
  HS65_LS_IVX9 U158 ( .A(\chs_in_f[4][DATA][29] ), .Z(n306) );
  HS65_LS_IVX9 U159 ( .A(\chs_in_f[4][DATA][30] ), .Z(n305) );
  HS65_LS_IVX9 U160 ( .A(\chs_in_f[4][DATA][31] ), .Z(n304) );
  HS65_LS_IVX9 U161 ( .A(\chs_in_f[4][DATA][32] ), .Z(n303) );
  HS65_LS_BFX18 U162 ( .A(\switch_sel[2][4] ), .Z(n77) );
  HS65_LS_BFX18 U163 ( .A(\switch_sel[2][3] ), .Z(n73) );
  HS65_LS_BFX18 U164 ( .A(\switch_sel[0][2] ), .Z(n37) );
  HS65_LS_BFX18 U165 ( .A(\switch_sel[2][1] ), .Z(n69) );
  HS65_LS_BFX18 U166 ( .A(\switch_sel[2][0] ), .Z(n65) );
  HS65_LS_OAI212X5 U167 ( .A(n18), .B(n300), .C(n15), .D(n335), .E(n476), .Z(
        \chs_out_f[4][DATA][0] ) );
  HS65_LS_AOI222X2 U168 ( .A(\chs_in_f[2][DATA][0] ), .B(n80), .C(
        \chs_in_f[0][DATA][0] ), .D(n46), .E(\chs_in_f[1][DATA][0] ), .F(n64), 
        .Z(n476) );
  HS65_LS_OAI212X5 U169 ( .A(n18), .B(n299), .C(n15), .D(n334), .E(n487), .Z(
        \chs_out_f[4][DATA][1] ) );
  HS65_LS_AOI222X2 U170 ( .A(\chs_in_f[2][DATA][1] ), .B(n79), .C(
        \chs_in_f[0][DATA][1] ), .D(n46), .E(\chs_in_f[1][DATA][1] ), .F(n63), 
        .Z(n487) );
  HS65_LS_OAI212X5 U171 ( .A(n19), .B(n298), .C(n16), .D(n333), .E(n498), .Z(
        \chs_out_f[4][DATA][2] ) );
  HS65_LS_AOI222X2 U172 ( .A(\chs_in_f[2][DATA][2] ), .B(n78), .C(
        \chs_in_f[0][DATA][2] ), .D(n47), .E(\chs_in_f[1][DATA][2] ), .F(n62), 
        .Z(n498) );
  HS65_LS_OAI212X5 U173 ( .A(n20), .B(n297), .C(n17), .D(n332), .E(n504), .Z(
        \chs_out_f[4][DATA][3] ) );
  HS65_LS_AOI222X2 U174 ( .A(\chs_in_f[2][DATA][3] ), .B(n78), .C(
        \chs_in_f[0][DATA][3] ), .D(n48), .E(\chs_in_f[1][DATA][3] ), .F(n62), 
        .Z(n504) );
  HS65_LS_OAI212X5 U175 ( .A(n20), .B(n296), .C(n17), .D(n331), .E(n505), .Z(
        \chs_out_f[4][DATA][4] ) );
  HS65_LS_AOI222X2 U176 ( .A(\chs_in_f[2][DATA][4] ), .B(n78), .C(
        \chs_in_f[0][DATA][4] ), .D(n48), .E(\chs_in_f[1][DATA][4] ), .F(n62), 
        .Z(n505) );
  HS65_LS_OAI212X5 U177 ( .A(n20), .B(n295), .C(n17), .D(n330), .E(n506), .Z(
        \chs_out_f[4][DATA][5] ) );
  HS65_LS_AOI222X2 U178 ( .A(\chs_in_f[2][DATA][5] ), .B(n78), .C(
        \chs_in_f[0][DATA][5] ), .D(n48), .E(\chs_in_f[1][DATA][5] ), .F(n62), 
        .Z(n506) );
  HS65_LS_OAI212X5 U179 ( .A(n20), .B(n294), .C(n17), .D(n329), .E(n507), .Z(
        \chs_out_f[4][DATA][6] ) );
  HS65_LS_AOI222X2 U180 ( .A(\chs_in_f[2][DATA][6] ), .B(n78), .C(
        \chs_in_f[0][DATA][6] ), .D(n48), .E(\chs_in_f[1][DATA][6] ), .F(n62), 
        .Z(n507) );
  HS65_LS_OAI212X5 U181 ( .A(n20), .B(n293), .C(n17), .D(n328), .E(n508), .Z(
        \chs_out_f[4][DATA][7] ) );
  HS65_LS_AOI222X2 U182 ( .A(\chs_in_f[2][DATA][7] ), .B(n78), .C(
        \chs_in_f[0][DATA][7] ), .D(n48), .E(\chs_in_f[1][DATA][7] ), .F(n62), 
        .Z(n508) );
  HS65_LS_OAI212X5 U183 ( .A(n20), .B(n292), .C(n17), .D(n327), .E(n509), .Z(
        \chs_out_f[4][DATA][8] ) );
  HS65_LS_AOI222X2 U184 ( .A(\chs_in_f[2][DATA][8] ), .B(n78), .C(
        \chs_in_f[0][DATA][8] ), .D(n48), .E(\chs_in_f[1][DATA][8] ), .F(n62), 
        .Z(n509) );
  HS65_LS_OAI212X5 U185 ( .A(n18), .B(n290), .C(n15), .D(n325), .E(n477), .Z(
        \chs_out_f[4][DATA][10] ) );
  HS65_LS_AOI222X2 U186 ( .A(\chs_in_f[2][DATA][10] ), .B(n80), .C(
        \chs_in_f[0][DATA][10] ), .D(n46), .E(\chs_in_f[1][DATA][10] ), .F(n64), .Z(n477) );
  HS65_LS_OAI212X5 U187 ( .A(n18), .B(n289), .C(n15), .D(n324), .E(n478), .Z(
        \chs_out_f[4][DATA][11] ) );
  HS65_LS_AOI222X2 U188 ( .A(\chs_in_f[2][DATA][11] ), .B(n80), .C(
        \chs_in_f[0][DATA][11] ), .D(n46), .E(\chs_in_f[1][DATA][11] ), .F(n64), .Z(n478) );
  HS65_LS_OAI212X5 U189 ( .A(n18), .B(n288), .C(n15), .D(n323), .E(n479), .Z(
        \chs_out_f[4][DATA][12] ) );
  HS65_LS_AOI222X2 U190 ( .A(\chs_in_f[2][DATA][12] ), .B(n80), .C(
        \chs_in_f[0][DATA][12] ), .D(n46), .E(\chs_in_f[1][DATA][12] ), .F(n64), .Z(n479) );
  HS65_LS_OAI212X5 U191 ( .A(n18), .B(n287), .C(n15), .D(n322), .E(n480), .Z(
        \chs_out_f[4][DATA][13] ) );
  HS65_LS_AOI222X2 U192 ( .A(\chs_in_f[2][DATA][13] ), .B(n80), .C(
        \chs_in_f[0][DATA][13] ), .D(n46), .E(\chs_in_f[1][DATA][13] ), .F(n64), .Z(n480) );
  HS65_LS_OAI212X5 U193 ( .A(n18), .B(n286), .C(n15), .D(n321), .E(n481), .Z(
        \chs_out_f[4][DATA][14] ) );
  HS65_LS_AOI222X2 U194 ( .A(\chs_in_f[2][DATA][14] ), .B(n80), .C(
        \chs_in_f[0][DATA][14] ), .D(n46), .E(\chs_in_f[1][DATA][14] ), .F(n64), .Z(n481) );
  HS65_LS_OAI212X5 U195 ( .A(n18), .B(n285), .C(n15), .D(n320), .E(n482), .Z(
        \chs_out_f[4][DATA][15] ) );
  HS65_LS_AOI222X2 U196 ( .A(\chs_in_f[2][DATA][15] ), .B(n80), .C(
        \chs_in_f[0][DATA][15] ), .D(n46), .E(\chs_in_f[1][DATA][15] ), .F(n64), .Z(n482) );
  HS65_LS_OAI212X5 U197 ( .A(n18), .B(n284), .C(n15), .D(n319), .E(n483), .Z(
        \chs_out_f[4][DATA][16] ) );
  HS65_LS_AOI222X2 U198 ( .A(\chs_in_f[2][DATA][16] ), .B(n80), .C(
        \chs_in_f[0][DATA][16] ), .D(n46), .E(\chs_in_f[1][DATA][16] ), .F(n64), .Z(n483) );
  HS65_LS_OAI212X5 U199 ( .A(n18), .B(n283), .C(n15), .D(n318), .E(n484), .Z(
        \chs_out_f[4][DATA][17] ) );
  HS65_LS_AOI222X2 U200 ( .A(\chs_in_f[2][DATA][17] ), .B(n80), .C(
        \chs_in_f[0][DATA][17] ), .D(n46), .E(\chs_in_f[1][DATA][17] ), .F(n64), .Z(n484) );
  HS65_LS_OAI212X5 U201 ( .A(n18), .B(n282), .C(n15), .D(n317), .E(n485), .Z(
        \chs_out_f[4][DATA][18] ) );
  HS65_LS_AOI222X2 U202 ( .A(\chs_in_f[2][DATA][18] ), .B(n79), .C(
        \chs_in_f[0][DATA][18] ), .D(n46), .E(\chs_in_f[1][DATA][18] ), .F(n63), .Z(n485) );
  HS65_LS_OAI212X5 U203 ( .A(n18), .B(n281), .C(n15), .D(n316), .E(n486), .Z(
        \chs_out_f[4][DATA][19] ) );
  HS65_LS_AOI222X2 U204 ( .A(\chs_in_f[2][DATA][19] ), .B(n79), .C(
        \chs_in_f[0][DATA][19] ), .D(n46), .E(\chs_in_f[1][DATA][19] ), .F(n63), .Z(n486) );
  HS65_LS_OAI212X5 U205 ( .A(n19), .B(n280), .C(n15), .D(n315), .E(n488), .Z(
        \chs_out_f[4][DATA][20] ) );
  HS65_LS_AOI222X2 U206 ( .A(\chs_in_f[2][DATA][20] ), .B(n79), .C(
        \chs_in_f[0][DATA][20] ), .D(n47), .E(\chs_in_f[1][DATA][20] ), .F(n63), .Z(n488) );
  HS65_LS_OAI212X5 U207 ( .A(n19), .B(n279), .C(n16), .D(n314), .E(n489), .Z(
        \chs_out_f[4][DATA][21] ) );
  HS65_LS_AOI222X2 U208 ( .A(\chs_in_f[2][DATA][21] ), .B(n79), .C(
        \chs_in_f[0][DATA][21] ), .D(n47), .E(\chs_in_f[1][DATA][21] ), .F(n63), .Z(n489) );
  HS65_LS_OAI212X5 U209 ( .A(n19), .B(n278), .C(n16), .D(n313), .E(n490), .Z(
        \chs_out_f[4][DATA][22] ) );
  HS65_LS_AOI222X2 U210 ( .A(\chs_in_f[2][DATA][22] ), .B(n79), .C(
        \chs_in_f[0][DATA][22] ), .D(n47), .E(\chs_in_f[1][DATA][22] ), .F(n63), .Z(n490) );
  HS65_LS_OAI212X5 U211 ( .A(n19), .B(n277), .C(n16), .D(n312), .E(n491), .Z(
        \chs_out_f[4][DATA][23] ) );
  HS65_LS_AOI222X2 U212 ( .A(\chs_in_f[2][DATA][23] ), .B(n79), .C(
        \chs_in_f[0][DATA][23] ), .D(n47), .E(\chs_in_f[1][DATA][23] ), .F(n63), .Z(n491) );
  HS65_LS_OAI212X5 U213 ( .A(n19), .B(n276), .C(n16), .D(n311), .E(n492), .Z(
        \chs_out_f[4][DATA][24] ) );
  HS65_LS_AOI222X2 U214 ( .A(\chs_in_f[2][DATA][24] ), .B(n79), .C(
        \chs_in_f[0][DATA][24] ), .D(n47), .E(\chs_in_f[1][DATA][24] ), .F(n63), .Z(n492) );
  HS65_LS_OAI212X5 U215 ( .A(n19), .B(n275), .C(n16), .D(n310), .E(n493), .Z(
        \chs_out_f[4][DATA][25] ) );
  HS65_LS_AOI222X2 U216 ( .A(\chs_in_f[2][DATA][25] ), .B(n79), .C(
        \chs_in_f[0][DATA][25] ), .D(n47), .E(\chs_in_f[1][DATA][25] ), .F(n63), .Z(n493) );
  HS65_LS_OAI212X5 U217 ( .A(n19), .B(n274), .C(n16), .D(n309), .E(n494), .Z(
        \chs_out_f[4][DATA][26] ) );
  HS65_LS_AOI222X2 U218 ( .A(\chs_in_f[2][DATA][26] ), .B(n79), .C(
        \chs_in_f[0][DATA][26] ), .D(n47), .E(\chs_in_f[1][DATA][26] ), .F(n63), .Z(n494) );
  HS65_LS_OAI212X5 U219 ( .A(n19), .B(n273), .C(n16), .D(n308), .E(n495), .Z(
        \chs_out_f[4][DATA][27] ) );
  HS65_LS_AOI222X2 U220 ( .A(\chs_in_f[2][DATA][27] ), .B(n79), .C(
        \chs_in_f[0][DATA][27] ), .D(n47), .E(\chs_in_f[1][DATA][27] ), .F(n63), .Z(n495) );
  HS65_LS_OAI212X5 U221 ( .A(n19), .B(n272), .C(n16), .D(n307), .E(n496), .Z(
        \chs_out_f[4][DATA][28] ) );
  HS65_LS_AOI222X2 U222 ( .A(\chs_in_f[2][DATA][28] ), .B(n79), .C(
        \chs_in_f[0][DATA][28] ), .D(n47), .E(\chs_in_f[1][DATA][28] ), .F(n63), .Z(n496) );
  HS65_LS_OAI212X5 U223 ( .A(n19), .B(n271), .C(n16), .D(n306), .E(n497), .Z(
        \chs_out_f[4][DATA][29] ) );
  HS65_LS_AOI222X2 U224 ( .A(\chs_in_f[2][DATA][29] ), .B(n79), .C(
        \chs_in_f[0][DATA][29] ), .D(n47), .E(\chs_in_f[1][DATA][29] ), .F(n63), .Z(n497) );
  HS65_LS_OAI212X5 U225 ( .A(n19), .B(n270), .C(n16), .D(n305), .E(n499), .Z(
        \chs_out_f[4][DATA][30] ) );
  HS65_LS_AOI222X2 U226 ( .A(\chs_in_f[2][DATA][30] ), .B(n78), .C(
        \chs_in_f[0][DATA][30] ), .D(n47), .E(\chs_in_f[1][DATA][30] ), .F(n62), .Z(n499) );
  HS65_LS_OAI212X5 U227 ( .A(n20), .B(n269), .C(n16), .D(n304), .E(n500), .Z(
        \chs_out_f[4][DATA][31] ) );
  HS65_LS_AOI222X2 U228 ( .A(\chs_in_f[2][DATA][31] ), .B(n78), .C(
        \chs_in_f[0][DATA][31] ), .D(n48), .E(\chs_in_f[1][DATA][31] ), .F(n62), .Z(n500) );
  HS65_LS_OAI212X5 U229 ( .A(n20), .B(n268), .C(n16), .D(n303), .E(n501), .Z(
        \chs_out_f[4][DATA][32] ) );
  HS65_LS_AOI222X2 U230 ( .A(\chs_in_f[2][DATA][32] ), .B(n78), .C(
        \chs_in_f[0][DATA][32] ), .D(n48), .E(\chs_in_f[1][DATA][32] ), .F(n62), .Z(n501) );
  HS65_LS_OAI212X5 U231 ( .A(n20), .B(n267), .C(n17), .D(n302), .E(n502), .Z(
        \chs_out_f[4][DATA][33] ) );
  HS65_LS_AOI222X2 U232 ( .A(\chs_in_f[2][DATA][33] ), .B(n78), .C(
        \chs_in_f[0][DATA][33] ), .D(n48), .E(\chs_in_f[1][DATA][33] ), .F(n62), .Z(n502) );
  HS65_LS_OAI212X5 U233 ( .A(n291), .B(n23), .C(n326), .D(n8), .E(n440), .Z(
        \chs_out_f[2][DATA][9] ) );
  HS65_LS_AOI222X2 U234 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][9] ), 
        .C(n40), .D(\chs_in_f[0][DATA][9] ), .E(n56), .F(
        \chs_in_f[1][DATA][9] ), .Z(n440) );
  HS65_LS_OAI212X5 U235 ( .A(n291), .B(n26), .C(n326), .D(n11), .E(n405), .Z(
        \chs_out_f[1][DATA][9] ) );
  HS65_LS_AOI222X2 U236 ( .A(n72), .B(\chs_in_f[2][DATA][9] ), .C(n36), .D(
        \chs_in_f[0][DATA][9] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][9] ), .Z(n405) );
  HS65_LS_OAI212X5 U237 ( .A(n291), .B(n29), .C(n326), .D(n14), .E(n370), .Z(
        \chs_out_f[0][DATA][9] ) );
  HS65_LS_AOI222X2 U238 ( .A(n68), .B(\chs_in_f[2][DATA][9] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][9] ), .E(n52), .F(
        \chs_in_f[1][DATA][9] ), .Z(n370) );
  HS65_LS_OAI212X5 U239 ( .A(n300), .B(n21), .C(n335), .D(n6), .E(n406), .Z(
        \chs_out_f[2][DATA][0] ) );
  HS65_LS_AOI222X2 U240 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][0] ), 
        .C(n38), .D(\chs_in_f[0][DATA][0] ), .E(n54), .F(
        \chs_in_f[1][DATA][0] ), .Z(n406) );
  HS65_LS_OAI212X5 U241 ( .A(n299), .B(n21), .C(n334), .D(n6), .E(n417), .Z(
        \chs_out_f[2][DATA][1] ) );
  HS65_LS_AOI222X2 U242 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][1] ), 
        .C(n38), .D(\chs_in_f[0][DATA][1] ), .E(n54), .F(
        \chs_in_f[1][DATA][1] ), .Z(n417) );
  HS65_LS_OAI212X5 U243 ( .A(n298), .B(n22), .C(n333), .D(n7), .E(n428), .Z(
        \chs_out_f[2][DATA][2] ) );
  HS65_LS_AOI222X2 U244 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][2] ), 
        .C(n39), .D(\chs_in_f[0][DATA][2] ), .E(n55), .F(
        \chs_in_f[1][DATA][2] ), .Z(n428) );
  HS65_LS_OAI212X5 U245 ( .A(n290), .B(n21), .C(n325), .D(n6), .E(n407), .Z(
        \chs_out_f[2][DATA][10] ) );
  HS65_LS_AOI222X2 U246 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][10] ), 
        .C(n38), .D(\chs_in_f[0][DATA][10] ), .E(n54), .F(
        \chs_in_f[1][DATA][10] ), .Z(n407) );
  HS65_LS_OAI212X5 U247 ( .A(n289), .B(n21), .C(n324), .D(n6), .E(n408), .Z(
        \chs_out_f[2][DATA][11] ) );
  HS65_LS_AOI222X2 U248 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][11] ), 
        .C(n38), .D(\chs_in_f[0][DATA][11] ), .E(n54), .F(
        \chs_in_f[1][DATA][11] ), .Z(n408) );
  HS65_LS_OAI212X5 U249 ( .A(n288), .B(n21), .C(n323), .D(n6), .E(n409), .Z(
        \chs_out_f[2][DATA][12] ) );
  HS65_LS_AOI222X2 U250 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][12] ), 
        .C(n38), .D(\chs_in_f[0][DATA][12] ), .E(n54), .F(
        \chs_in_f[1][DATA][12] ), .Z(n409) );
  HS65_LS_OAI212X5 U251 ( .A(n287), .B(n21), .C(n322), .D(n6), .E(n410), .Z(
        \chs_out_f[2][DATA][13] ) );
  HS65_LS_AOI222X2 U252 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][13] ), 
        .C(n38), .D(\chs_in_f[0][DATA][13] ), .E(n54), .F(
        \chs_in_f[1][DATA][13] ), .Z(n410) );
  HS65_LS_OAI212X5 U253 ( .A(n286), .B(n21), .C(n321), .D(n6), .E(n411), .Z(
        \chs_out_f[2][DATA][14] ) );
  HS65_LS_AOI222X2 U254 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][14] ), 
        .C(n38), .D(\chs_in_f[0][DATA][14] ), .E(n54), .F(
        \chs_in_f[1][DATA][14] ), .Z(n411) );
  HS65_LS_OAI212X5 U255 ( .A(n285), .B(n21), .C(n320), .D(n6), .E(n412), .Z(
        \chs_out_f[2][DATA][15] ) );
  HS65_LS_AOI222X2 U256 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][15] ), 
        .C(n38), .D(\chs_in_f[0][DATA][15] ), .E(n54), .F(
        \chs_in_f[1][DATA][15] ), .Z(n412) );
  HS65_LS_OAI212X5 U257 ( .A(n284), .B(n21), .C(n319), .D(n6), .E(n413), .Z(
        \chs_out_f[2][DATA][16] ) );
  HS65_LS_AOI222X2 U258 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][16] ), 
        .C(n38), .D(\chs_in_f[0][DATA][16] ), .E(n54), .F(
        \chs_in_f[1][DATA][16] ), .Z(n413) );
  HS65_LS_OAI212X5 U259 ( .A(n283), .B(n21), .C(n318), .D(n6), .E(n414), .Z(
        \chs_out_f[2][DATA][17] ) );
  HS65_LS_AOI222X2 U260 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][17] ), 
        .C(n38), .D(\chs_in_f[0][DATA][17] ), .E(n54), .F(
        \chs_in_f[1][DATA][17] ), .Z(n414) );
  HS65_LS_OAI212X5 U261 ( .A(n282), .B(n21), .C(n317), .D(n6), .E(n415), .Z(
        \chs_out_f[2][DATA][18] ) );
  HS65_LS_AOI222X2 U262 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][18] ), 
        .C(n38), .D(\chs_in_f[0][DATA][18] ), .E(n54), .F(
        \chs_in_f[1][DATA][18] ), .Z(n415) );
  HS65_LS_OAI212X5 U263 ( .A(n281), .B(n21), .C(n316), .D(n6), .E(n416), .Z(
        \chs_out_f[2][DATA][19] ) );
  HS65_LS_AOI222X2 U264 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][19] ), 
        .C(n38), .D(\chs_in_f[0][DATA][19] ), .E(n54), .F(
        \chs_in_f[1][DATA][19] ), .Z(n416) );
  HS65_LS_OAI212X5 U265 ( .A(n280), .B(n21), .C(n315), .D(n7), .E(n418), .Z(
        \chs_out_f[2][DATA][20] ) );
  HS65_LS_AOI222X2 U266 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][20] ), 
        .C(n39), .D(\chs_in_f[0][DATA][20] ), .E(n55), .F(
        \chs_in_f[1][DATA][20] ), .Z(n418) );
  HS65_LS_OAI212X5 U267 ( .A(n279), .B(n22), .C(n314), .D(n7), .E(n419), .Z(
        \chs_out_f[2][DATA][21] ) );
  HS65_LS_AOI222X2 U268 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][21] ), 
        .C(n39), .D(\chs_in_f[0][DATA][21] ), .E(n55), .F(
        \chs_in_f[1][DATA][21] ), .Z(n419) );
  HS65_LS_OAI212X5 U269 ( .A(n278), .B(n22), .C(n313), .D(n7), .E(n420), .Z(
        \chs_out_f[2][DATA][22] ) );
  HS65_LS_AOI222X2 U270 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][22] ), 
        .C(n39), .D(\chs_in_f[0][DATA][22] ), .E(n55), .F(
        \chs_in_f[1][DATA][22] ), .Z(n420) );
  HS65_LS_OAI212X5 U271 ( .A(n277), .B(n22), .C(n312), .D(n7), .E(n421), .Z(
        \chs_out_f[2][DATA][23] ) );
  HS65_LS_AOI222X2 U272 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][23] ), 
        .C(n39), .D(\chs_in_f[0][DATA][23] ), .E(n55), .F(
        \chs_in_f[1][DATA][23] ), .Z(n421) );
  HS65_LS_OAI212X5 U273 ( .A(n276), .B(n22), .C(n311), .D(n7), .E(n422), .Z(
        \chs_out_f[2][DATA][24] ) );
  HS65_LS_AOI222X2 U274 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][24] ), 
        .C(n39), .D(\chs_in_f[0][DATA][24] ), .E(n55), .F(
        \chs_in_f[1][DATA][24] ), .Z(n422) );
  HS65_LS_OAI212X5 U275 ( .A(n275), .B(n22), .C(n310), .D(n7), .E(n423), .Z(
        \chs_out_f[2][DATA][25] ) );
  HS65_LS_AOI222X2 U276 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][25] ), 
        .C(n39), .D(\chs_in_f[0][DATA][25] ), .E(n55), .F(
        \chs_in_f[1][DATA][25] ), .Z(n423) );
  HS65_LS_OAI212X5 U277 ( .A(n274), .B(n22), .C(n309), .D(n7), .E(n424), .Z(
        \chs_out_f[2][DATA][26] ) );
  HS65_LS_AOI222X2 U278 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][26] ), 
        .C(n39), .D(\chs_in_f[0][DATA][26] ), .E(n55), .F(
        \chs_in_f[1][DATA][26] ), .Z(n424) );
  HS65_LS_OAI212X5 U279 ( .A(n273), .B(n22), .C(n308), .D(n7), .E(n425), .Z(
        \chs_out_f[2][DATA][27] ) );
  HS65_LS_AOI222X2 U280 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][27] ), 
        .C(n39), .D(\chs_in_f[0][DATA][27] ), .E(n55), .F(
        \chs_in_f[1][DATA][27] ), .Z(n425) );
  HS65_LS_OAI212X5 U281 ( .A(n272), .B(n22), .C(n307), .D(n7), .E(n426), .Z(
        \chs_out_f[2][DATA][28] ) );
  HS65_LS_AOI222X2 U282 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][28] ), 
        .C(n39), .D(\chs_in_f[0][DATA][28] ), .E(n55), .F(
        \chs_in_f[1][DATA][28] ), .Z(n426) );
  HS65_LS_OAI212X5 U283 ( .A(n271), .B(n22), .C(n306), .D(n7), .E(n427), .Z(
        \chs_out_f[2][DATA][29] ) );
  HS65_LS_AOI222X2 U284 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][29] ), 
        .C(n39), .D(\chs_in_f[0][DATA][29] ), .E(n55), .F(
        \chs_in_f[1][DATA][29] ), .Z(n427) );
  HS65_LS_OAI212X5 U285 ( .A(n270), .B(n22), .C(n305), .D(n7), .E(n429), .Z(
        \chs_out_f[2][DATA][30] ) );
  HS65_LS_AOI222X2 U286 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][30] ), 
        .C(n39), .D(\chs_in_f[0][DATA][30] ), .E(n55), .F(
        \chs_in_f[1][DATA][30] ), .Z(n429) );
  HS65_LS_OAI212X5 U287 ( .A(n269), .B(n22), .C(n304), .D(n8), .E(n430), .Z(
        \chs_out_f[2][DATA][31] ) );
  HS65_LS_AOI222X2 U288 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][31] ), 
        .C(n40), .D(\chs_in_f[0][DATA][31] ), .E(n56), .F(
        \chs_in_f[1][DATA][31] ), .Z(n430) );
  HS65_LS_OAI212X5 U289 ( .A(n268), .B(n22), .C(n303), .D(n8), .E(n431), .Z(
        \chs_out_f[2][DATA][32] ) );
  HS65_LS_AOI222X2 U290 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][32] ), 
        .C(n40), .D(\chs_in_f[0][DATA][32] ), .E(n56), .F(
        \chs_in_f[1][DATA][32] ), .Z(n431) );
  HS65_LS_OAI212X5 U291 ( .A(n300), .B(n24), .C(n335), .D(n9), .E(n371), .Z(
        \chs_out_f[1][DATA][0] ) );
  HS65_LS_AOI222X2 U292 ( .A(n70), .B(\chs_in_f[2][DATA][0] ), .C(n34), .D(
        \chs_in_f[0][DATA][0] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][0] ), .Z(n371) );
  HS65_LS_OAI212X5 U293 ( .A(n299), .B(n24), .C(n334), .D(n9), .E(n382), .Z(
        \chs_out_f[1][DATA][1] ) );
  HS65_LS_AOI222X2 U294 ( .A(n70), .B(\chs_in_f[2][DATA][1] ), .C(n34), .D(
        \chs_in_f[0][DATA][1] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][1] ), .Z(n382) );
  HS65_LS_OAI212X5 U295 ( .A(n298), .B(n25), .C(n333), .D(n10), .E(n393), .Z(
        \chs_out_f[1][DATA][2] ) );
  HS65_LS_AOI222X2 U296 ( .A(n71), .B(\chs_in_f[2][DATA][2] ), .C(n35), .D(
        \chs_in_f[0][DATA][2] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][2] ), .Z(n393) );
  HS65_LS_OAI212X5 U297 ( .A(n290), .B(n24), .C(n325), .D(n9), .E(n372), .Z(
        \chs_out_f[1][DATA][10] ) );
  HS65_LS_AOI222X2 U298 ( .A(n70), .B(\chs_in_f[2][DATA][10] ), .C(n34), .D(
        \chs_in_f[0][DATA][10] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][10] ), .Z(n372) );
  HS65_LS_OAI212X5 U299 ( .A(n289), .B(n24), .C(n324), .D(n9), .E(n373), .Z(
        \chs_out_f[1][DATA][11] ) );
  HS65_LS_AOI222X2 U300 ( .A(n70), .B(\chs_in_f[2][DATA][11] ), .C(n34), .D(
        \chs_in_f[0][DATA][11] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][11] ), .Z(n373) );
  HS65_LS_OAI212X5 U301 ( .A(n288), .B(n24), .C(n323), .D(n9), .E(n374), .Z(
        \chs_out_f[1][DATA][12] ) );
  HS65_LS_AOI222X2 U302 ( .A(n70), .B(\chs_in_f[2][DATA][12] ), .C(n34), .D(
        \chs_in_f[0][DATA][12] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][12] ), .Z(n374) );
  HS65_LS_OAI212X5 U303 ( .A(n287), .B(n24), .C(n322), .D(n9), .E(n375), .Z(
        \chs_out_f[1][DATA][13] ) );
  HS65_LS_AOI222X2 U304 ( .A(n70), .B(\chs_in_f[2][DATA][13] ), .C(n34), .D(
        \chs_in_f[0][DATA][13] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][13] ), .Z(n375) );
  HS65_LS_OAI212X5 U305 ( .A(n286), .B(n24), .C(n321), .D(n9), .E(n376), .Z(
        \chs_out_f[1][DATA][14] ) );
  HS65_LS_AOI222X2 U306 ( .A(n70), .B(\chs_in_f[2][DATA][14] ), .C(n34), .D(
        \chs_in_f[0][DATA][14] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][14] ), .Z(n376) );
  HS65_LS_OAI212X5 U307 ( .A(n285), .B(n24), .C(n320), .D(n9), .E(n377), .Z(
        \chs_out_f[1][DATA][15] ) );
  HS65_LS_AOI222X2 U308 ( .A(n70), .B(\chs_in_f[2][DATA][15] ), .C(n34), .D(
        \chs_in_f[0][DATA][15] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][15] ), .Z(n377) );
  HS65_LS_OAI212X5 U309 ( .A(n284), .B(n24), .C(n319), .D(n9), .E(n378), .Z(
        \chs_out_f[1][DATA][16] ) );
  HS65_LS_AOI222X2 U310 ( .A(n70), .B(\chs_in_f[2][DATA][16] ), .C(n34), .D(
        \chs_in_f[0][DATA][16] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][16] ), .Z(n378) );
  HS65_LS_OAI212X5 U311 ( .A(n283), .B(n24), .C(n318), .D(n9), .E(n379), .Z(
        \chs_out_f[1][DATA][17] ) );
  HS65_LS_AOI222X2 U312 ( .A(n70), .B(\chs_in_f[2][DATA][17] ), .C(n34), .D(
        \chs_in_f[0][DATA][17] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][17] ), .Z(n379) );
  HS65_LS_OAI212X5 U313 ( .A(n282), .B(n24), .C(n317), .D(n9), .E(n380), .Z(
        \chs_out_f[1][DATA][18] ) );
  HS65_LS_AOI222X2 U314 ( .A(n70), .B(\chs_in_f[2][DATA][18] ), .C(n34), .D(
        \chs_in_f[0][DATA][18] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][18] ), .Z(n380) );
  HS65_LS_OAI212X5 U315 ( .A(n281), .B(n24), .C(n316), .D(n9), .E(n381), .Z(
        \chs_out_f[1][DATA][19] ) );
  HS65_LS_AOI222X2 U316 ( .A(n70), .B(\chs_in_f[2][DATA][19] ), .C(n34), .D(
        \chs_in_f[0][DATA][19] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][19] ), .Z(n381) );
  HS65_LS_OAI212X5 U317 ( .A(n280), .B(n24), .C(n315), .D(n10), .E(n383), .Z(
        \chs_out_f[1][DATA][20] ) );
  HS65_LS_AOI222X2 U318 ( .A(n71), .B(\chs_in_f[2][DATA][20] ), .C(n35), .D(
        \chs_in_f[0][DATA][20] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][20] ), .Z(n383) );
  HS65_LS_OAI212X5 U319 ( .A(n279), .B(n25), .C(n314), .D(n10), .E(n384), .Z(
        \chs_out_f[1][DATA][21] ) );
  HS65_LS_AOI222X2 U320 ( .A(n71), .B(\chs_in_f[2][DATA][21] ), .C(n35), .D(
        \chs_in_f[0][DATA][21] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][21] ), .Z(n384) );
  HS65_LS_OAI212X5 U321 ( .A(n278), .B(n25), .C(n313), .D(n10), .E(n385), .Z(
        \chs_out_f[1][DATA][22] ) );
  HS65_LS_AOI222X2 U322 ( .A(n71), .B(\chs_in_f[2][DATA][22] ), .C(n35), .D(
        \chs_in_f[0][DATA][22] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][22] ), .Z(n385) );
  HS65_LS_OAI212X5 U323 ( .A(n277), .B(n25), .C(n312), .D(n10), .E(n386), .Z(
        \chs_out_f[1][DATA][23] ) );
  HS65_LS_AOI222X2 U324 ( .A(n71), .B(\chs_in_f[2][DATA][23] ), .C(n35), .D(
        \chs_in_f[0][DATA][23] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][23] ), .Z(n386) );
  HS65_LS_OAI212X5 U325 ( .A(n276), .B(n25), .C(n311), .D(n10), .E(n387), .Z(
        \chs_out_f[1][DATA][24] ) );
  HS65_LS_AOI222X2 U326 ( .A(n71), .B(\chs_in_f[2][DATA][24] ), .C(n35), .D(
        \chs_in_f[0][DATA][24] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][24] ), .Z(n387) );
  HS65_LS_OAI212X5 U327 ( .A(n275), .B(n25), .C(n310), .D(n10), .E(n388), .Z(
        \chs_out_f[1][DATA][25] ) );
  HS65_LS_AOI222X2 U328 ( .A(n71), .B(\chs_in_f[2][DATA][25] ), .C(n35), .D(
        \chs_in_f[0][DATA][25] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][25] ), .Z(n388) );
  HS65_LS_OAI212X5 U329 ( .A(n274), .B(n25), .C(n309), .D(n10), .E(n389), .Z(
        \chs_out_f[1][DATA][26] ) );
  HS65_LS_AOI222X2 U330 ( .A(n71), .B(\chs_in_f[2][DATA][26] ), .C(n35), .D(
        \chs_in_f[0][DATA][26] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][26] ), .Z(n389) );
  HS65_LS_OAI212X5 U331 ( .A(n273), .B(n25), .C(n308), .D(n10), .E(n390), .Z(
        \chs_out_f[1][DATA][27] ) );
  HS65_LS_AOI222X2 U332 ( .A(n71), .B(\chs_in_f[2][DATA][27] ), .C(n35), .D(
        \chs_in_f[0][DATA][27] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][27] ), .Z(n390) );
  HS65_LS_OAI212X5 U333 ( .A(n272), .B(n25), .C(n307), .D(n10), .E(n391), .Z(
        \chs_out_f[1][DATA][28] ) );
  HS65_LS_AOI222X2 U334 ( .A(n71), .B(\chs_in_f[2][DATA][28] ), .C(n35), .D(
        \chs_in_f[0][DATA][28] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][28] ), .Z(n391) );
  HS65_LS_OAI212X5 U335 ( .A(n271), .B(n25), .C(n306), .D(n10), .E(n392), .Z(
        \chs_out_f[1][DATA][29] ) );
  HS65_LS_AOI222X2 U336 ( .A(n71), .B(\chs_in_f[2][DATA][29] ), .C(n35), .D(
        \chs_in_f[0][DATA][29] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][29] ), .Z(n392) );
  HS65_LS_OAI212X5 U337 ( .A(n270), .B(n25), .C(n305), .D(n10), .E(n394), .Z(
        \chs_out_f[1][DATA][30] ) );
  HS65_LS_AOI222X2 U338 ( .A(n71), .B(\chs_in_f[2][DATA][30] ), .C(n35), .D(
        \chs_in_f[0][DATA][30] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][30] ), .Z(n394) );
  HS65_LS_OAI212X5 U339 ( .A(n269), .B(n25), .C(n304), .D(n11), .E(n395), .Z(
        \chs_out_f[1][DATA][31] ) );
  HS65_LS_AOI222X2 U340 ( .A(n72), .B(\chs_in_f[2][DATA][31] ), .C(n36), .D(
        \chs_in_f[0][DATA][31] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][31] ), .Z(n395) );
  HS65_LS_OAI212X5 U341 ( .A(n268), .B(n25), .C(n303), .D(n11), .E(n396), .Z(
        \chs_out_f[1][DATA][32] ) );
  HS65_LS_AOI222X2 U342 ( .A(n72), .B(\chs_in_f[2][DATA][32] ), .C(n36), .D(
        \chs_in_f[0][DATA][32] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][32] ), .Z(n396) );
  HS65_LS_OAI212X5 U343 ( .A(n300), .B(n27), .C(n335), .D(n12), .E(n336), .Z(
        \chs_out_f[0][DATA][0] ) );
  HS65_LS_AOI222X2 U344 ( .A(n66), .B(\chs_in_f[2][DATA][0] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][0] ), .E(n50), .F(
        \chs_in_f[1][DATA][0] ), .Z(n336) );
  HS65_LS_OAI212X5 U345 ( .A(n299), .B(n27), .C(n334), .D(n12), .E(n347), .Z(
        \chs_out_f[0][DATA][1] ) );
  HS65_LS_AOI222X2 U346 ( .A(n66), .B(\chs_in_f[2][DATA][1] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][1] ), .E(n50), .F(
        \chs_in_f[1][DATA][1] ), .Z(n347) );
  HS65_LS_OAI212X5 U347 ( .A(n298), .B(n28), .C(n333), .D(n13), .E(n358), .Z(
        \chs_out_f[0][DATA][2] ) );
  HS65_LS_AOI222X2 U348 ( .A(n67), .B(\chs_in_f[2][DATA][2] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][2] ), .E(n51), .F(
        \chs_in_f[1][DATA][2] ), .Z(n358) );
  HS65_LS_OAI212X5 U349 ( .A(n290), .B(n27), .C(n325), .D(n12), .E(n337), .Z(
        \chs_out_f[0][DATA][10] ) );
  HS65_LS_AOI222X2 U350 ( .A(n66), .B(\chs_in_f[2][DATA][10] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][10] ), .E(n50), .F(
        \chs_in_f[1][DATA][10] ), .Z(n337) );
  HS65_LS_OAI212X5 U351 ( .A(n289), .B(n27), .C(n324), .D(n12), .E(n338), .Z(
        \chs_out_f[0][DATA][11] ) );
  HS65_LS_AOI222X2 U352 ( .A(n66), .B(\chs_in_f[2][DATA][11] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][11] ), .E(n50), .F(
        \chs_in_f[1][DATA][11] ), .Z(n338) );
  HS65_LS_OAI212X5 U353 ( .A(n288), .B(n27), .C(n323), .D(n12), .E(n339), .Z(
        \chs_out_f[0][DATA][12] ) );
  HS65_LS_AOI222X2 U354 ( .A(n66), .B(\chs_in_f[2][DATA][12] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][12] ), .E(n50), .F(
        \chs_in_f[1][DATA][12] ), .Z(n339) );
  HS65_LS_OAI212X5 U355 ( .A(n287), .B(n27), .C(n322), .D(n12), .E(n340), .Z(
        \chs_out_f[0][DATA][13] ) );
  HS65_LS_AOI222X2 U356 ( .A(n66), .B(\chs_in_f[2][DATA][13] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][13] ), .E(n50), .F(
        \chs_in_f[1][DATA][13] ), .Z(n340) );
  HS65_LS_OAI212X5 U357 ( .A(n286), .B(n27), .C(n321), .D(n12), .E(n341), .Z(
        \chs_out_f[0][DATA][14] ) );
  HS65_LS_AOI222X2 U358 ( .A(n66), .B(\chs_in_f[2][DATA][14] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][14] ), .E(n50), .F(
        \chs_in_f[1][DATA][14] ), .Z(n341) );
  HS65_LS_OAI212X5 U359 ( .A(n285), .B(n27), .C(n320), .D(n12), .E(n342), .Z(
        \chs_out_f[0][DATA][15] ) );
  HS65_LS_AOI222X2 U360 ( .A(n66), .B(\chs_in_f[2][DATA][15] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][15] ), .E(n50), .F(
        \chs_in_f[1][DATA][15] ), .Z(n342) );
  HS65_LS_OAI212X5 U361 ( .A(n284), .B(n27), .C(n319), .D(n12), .E(n343), .Z(
        \chs_out_f[0][DATA][16] ) );
  HS65_LS_AOI222X2 U362 ( .A(n66), .B(\chs_in_f[2][DATA][16] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][16] ), .E(n50), .F(
        \chs_in_f[1][DATA][16] ), .Z(n343) );
  HS65_LS_OAI212X5 U363 ( .A(n283), .B(n27), .C(n318), .D(n12), .E(n344), .Z(
        \chs_out_f[0][DATA][17] ) );
  HS65_LS_AOI222X2 U364 ( .A(n66), .B(\chs_in_f[2][DATA][17] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][17] ), .E(n50), .F(
        \chs_in_f[1][DATA][17] ), .Z(n344) );
  HS65_LS_OAI212X5 U365 ( .A(n282), .B(n27), .C(n317), .D(n12), .E(n345), .Z(
        \chs_out_f[0][DATA][18] ) );
  HS65_LS_AOI222X2 U366 ( .A(n66), .B(\chs_in_f[2][DATA][18] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][18] ), .E(n50), .F(
        \chs_in_f[1][DATA][18] ), .Z(n345) );
  HS65_LS_OAI212X5 U367 ( .A(n281), .B(n27), .C(n316), .D(n12), .E(n346), .Z(
        \chs_out_f[0][DATA][19] ) );
  HS65_LS_AOI222X2 U368 ( .A(n66), .B(\chs_in_f[2][DATA][19] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][19] ), .E(n50), .F(
        \chs_in_f[1][DATA][19] ), .Z(n346) );
  HS65_LS_OAI212X5 U369 ( .A(n280), .B(n27), .C(n315), .D(n13), .E(n348), .Z(
        \chs_out_f[0][DATA][20] ) );
  HS65_LS_AOI222X2 U370 ( .A(n67), .B(\chs_in_f[2][DATA][20] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][20] ), .E(n51), .F(
        \chs_in_f[1][DATA][20] ), .Z(n348) );
  HS65_LS_OAI212X5 U371 ( .A(n279), .B(n28), .C(n314), .D(n13), .E(n349), .Z(
        \chs_out_f[0][DATA][21] ) );
  HS65_LS_AOI222X2 U372 ( .A(n67), .B(\chs_in_f[2][DATA][21] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][21] ), .E(n51), .F(
        \chs_in_f[1][DATA][21] ), .Z(n349) );
  HS65_LS_OAI212X5 U373 ( .A(n278), .B(n28), .C(n313), .D(n13), .E(n350), .Z(
        \chs_out_f[0][DATA][22] ) );
  HS65_LS_AOI222X2 U374 ( .A(n67), .B(\chs_in_f[2][DATA][22] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][22] ), .E(n51), .F(
        \chs_in_f[1][DATA][22] ), .Z(n350) );
  HS65_LS_OAI212X5 U375 ( .A(n277), .B(n28), .C(n312), .D(n13), .E(n351), .Z(
        \chs_out_f[0][DATA][23] ) );
  HS65_LS_AOI222X2 U376 ( .A(n67), .B(\chs_in_f[2][DATA][23] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][23] ), .E(n51), .F(
        \chs_in_f[1][DATA][23] ), .Z(n351) );
  HS65_LS_OAI212X5 U377 ( .A(n276), .B(n28), .C(n311), .D(n13), .E(n352), .Z(
        \chs_out_f[0][DATA][24] ) );
  HS65_LS_AOI222X2 U378 ( .A(n67), .B(\chs_in_f[2][DATA][24] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][24] ), .E(n51), .F(
        \chs_in_f[1][DATA][24] ), .Z(n352) );
  HS65_LS_OAI212X5 U379 ( .A(n275), .B(n28), .C(n310), .D(n13), .E(n353), .Z(
        \chs_out_f[0][DATA][25] ) );
  HS65_LS_AOI222X2 U380 ( .A(n67), .B(\chs_in_f[2][DATA][25] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][25] ), .E(n51), .F(
        \chs_in_f[1][DATA][25] ), .Z(n353) );
  HS65_LS_OAI212X5 U381 ( .A(n274), .B(n28), .C(n309), .D(n13), .E(n354), .Z(
        \chs_out_f[0][DATA][26] ) );
  HS65_LS_AOI222X2 U382 ( .A(n67), .B(\chs_in_f[2][DATA][26] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][26] ), .E(n51), .F(
        \chs_in_f[1][DATA][26] ), .Z(n354) );
  HS65_LS_OAI212X5 U383 ( .A(n273), .B(n28), .C(n308), .D(n13), .E(n355), .Z(
        \chs_out_f[0][DATA][27] ) );
  HS65_LS_AOI222X2 U384 ( .A(n67), .B(\chs_in_f[2][DATA][27] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][27] ), .E(n51), .F(
        \chs_in_f[1][DATA][27] ), .Z(n355) );
  HS65_LS_OAI212X5 U385 ( .A(n272), .B(n28), .C(n307), .D(n13), .E(n356), .Z(
        \chs_out_f[0][DATA][28] ) );
  HS65_LS_AOI222X2 U386 ( .A(n67), .B(\chs_in_f[2][DATA][28] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][28] ), .E(n51), .F(
        \chs_in_f[1][DATA][28] ), .Z(n356) );
  HS65_LS_OAI212X5 U387 ( .A(n271), .B(n28), .C(n306), .D(n13), .E(n357), .Z(
        \chs_out_f[0][DATA][29] ) );
  HS65_LS_AOI222X2 U388 ( .A(n67), .B(\chs_in_f[2][DATA][29] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][29] ), .E(n51), .F(
        \chs_in_f[1][DATA][29] ), .Z(n357) );
  HS65_LS_OAI212X5 U389 ( .A(n270), .B(n28), .C(n305), .D(n13), .E(n359), .Z(
        \chs_out_f[0][DATA][30] ) );
  HS65_LS_AOI222X2 U390 ( .A(n67), .B(\chs_in_f[2][DATA][30] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][30] ), .E(n51), .F(
        \chs_in_f[1][DATA][30] ), .Z(n359) );
  HS65_LS_OAI212X5 U391 ( .A(n269), .B(n28), .C(n304), .D(n14), .E(n360), .Z(
        \chs_out_f[0][DATA][31] ) );
  HS65_LS_AOI222X2 U392 ( .A(n68), .B(\chs_in_f[2][DATA][31] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][31] ), .E(n52), .F(
        \chs_in_f[1][DATA][31] ), .Z(n360) );
  HS65_LS_OAI212X5 U393 ( .A(n268), .B(n28), .C(n303), .D(n14), .E(n361), .Z(
        \chs_out_f[0][DATA][32] ) );
  HS65_LS_AOI222X2 U394 ( .A(n68), .B(\chs_in_f[2][DATA][32] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][32] ), .E(n52), .F(
        \chs_in_f[1][DATA][32] ), .Z(n361) );
  HS65_LS_OAI212X5 U395 ( .A(n297), .B(n23), .C(n332), .D(n8), .E(n434), .Z(
        \chs_out_f[2][DATA][3] ) );
  HS65_LS_AOI222X2 U396 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][3] ), 
        .C(n40), .D(\chs_in_f[0][DATA][3] ), .E(n56), .F(
        \chs_in_f[1][DATA][3] ), .Z(n434) );
  HS65_LS_OAI212X5 U397 ( .A(n296), .B(n23), .C(n331), .D(n8), .E(n435), .Z(
        \chs_out_f[2][DATA][4] ) );
  HS65_LS_AOI222X2 U398 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][4] ), 
        .C(n40), .D(\chs_in_f[0][DATA][4] ), .E(n56), .F(
        \chs_in_f[1][DATA][4] ), .Z(n435) );
  HS65_LS_OAI212X5 U399 ( .A(n295), .B(n23), .C(n330), .D(n8), .E(n436), .Z(
        \chs_out_f[2][DATA][5] ) );
  HS65_LS_AOI222X2 U400 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][5] ), 
        .C(n40), .D(\chs_in_f[0][DATA][5] ), .E(n56), .F(
        \chs_in_f[1][DATA][5] ), .Z(n436) );
  HS65_LS_OAI212X5 U401 ( .A(n294), .B(n23), .C(n329), .D(n8), .E(n437), .Z(
        \chs_out_f[2][DATA][6] ) );
  HS65_LS_AOI222X2 U402 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][6] ), 
        .C(n40), .D(\chs_in_f[0][DATA][6] ), .E(n56), .F(
        \chs_in_f[1][DATA][6] ), .Z(n437) );
  HS65_LS_OAI212X5 U403 ( .A(n293), .B(n23), .C(n328), .D(n8), .E(n438), .Z(
        \chs_out_f[2][DATA][7] ) );
  HS65_LS_AOI222X2 U404 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][7] ), 
        .C(n40), .D(\chs_in_f[0][DATA][7] ), .E(n56), .F(
        \chs_in_f[1][DATA][7] ), .Z(n438) );
  HS65_LS_OAI212X5 U405 ( .A(n292), .B(n23), .C(n327), .D(n8), .E(n439), .Z(
        \chs_out_f[2][DATA][8] ) );
  HS65_LS_AOI222X2 U406 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][8] ), 
        .C(n40), .D(\chs_in_f[0][DATA][8] ), .E(n56), .F(
        \chs_in_f[1][DATA][8] ), .Z(n439) );
  HS65_LS_OAI212X5 U407 ( .A(n267), .B(n23), .C(n302), .D(n8), .E(n432), .Z(
        \chs_out_f[2][DATA][33] ) );
  HS65_LS_AOI222X2 U408 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][33] ), 
        .C(n40), .D(\chs_in_f[0][DATA][33] ), .E(n56), .F(
        \chs_in_f[1][DATA][33] ), .Z(n432) );
  HS65_LS_OAI212X5 U409 ( .A(n297), .B(n26), .C(n332), .D(n11), .E(n399), .Z(
        \chs_out_f[1][DATA][3] ) );
  HS65_LS_AOI222X2 U410 ( .A(n72), .B(\chs_in_f[2][DATA][3] ), .C(n36), .D(
        \chs_in_f[0][DATA][3] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][3] ), .Z(n399) );
  HS65_LS_OAI212X5 U411 ( .A(n296), .B(n26), .C(n331), .D(n11), .E(n400), .Z(
        \chs_out_f[1][DATA][4] ) );
  HS65_LS_AOI222X2 U412 ( .A(n72), .B(\chs_in_f[2][DATA][4] ), .C(n36), .D(
        \chs_in_f[0][DATA][4] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][4] ), .Z(n400) );
  HS65_LS_OAI212X5 U413 ( .A(n295), .B(n26), .C(n330), .D(n11), .E(n401), .Z(
        \chs_out_f[1][DATA][5] ) );
  HS65_LS_AOI222X2 U414 ( .A(n72), .B(\chs_in_f[2][DATA][5] ), .C(n36), .D(
        \chs_in_f[0][DATA][5] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][5] ), .Z(n401) );
  HS65_LS_OAI212X5 U415 ( .A(n294), .B(n26), .C(n329), .D(n11), .E(n402), .Z(
        \chs_out_f[1][DATA][6] ) );
  HS65_LS_AOI222X2 U416 ( .A(n72), .B(\chs_in_f[2][DATA][6] ), .C(n36), .D(
        \chs_in_f[0][DATA][6] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][6] ), .Z(n402) );
  HS65_LS_OAI212X5 U417 ( .A(n293), .B(n26), .C(n328), .D(n11), .E(n403), .Z(
        \chs_out_f[1][DATA][7] ) );
  HS65_LS_AOI222X2 U418 ( .A(n72), .B(\chs_in_f[2][DATA][7] ), .C(n36), .D(
        \chs_in_f[0][DATA][7] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][7] ), .Z(n403) );
  HS65_LS_OAI212X5 U419 ( .A(n292), .B(n26), .C(n327), .D(n11), .E(n404), .Z(
        \chs_out_f[1][DATA][8] ) );
  HS65_LS_AOI222X2 U420 ( .A(n72), .B(\chs_in_f[2][DATA][8] ), .C(n36), .D(
        \chs_in_f[0][DATA][8] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][8] ), .Z(n404) );
  HS65_LS_OAI212X5 U421 ( .A(n267), .B(n26), .C(n302), .D(n11), .E(n397), .Z(
        \chs_out_f[1][DATA][33] ) );
  HS65_LS_AOI222X2 U422 ( .A(n72), .B(\chs_in_f[2][DATA][33] ), .C(n36), .D(
        \chs_in_f[0][DATA][33] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][33] ), .Z(n397) );
  HS65_LS_OAI212X5 U423 ( .A(n297), .B(n29), .C(n332), .D(n14), .E(n364), .Z(
        \chs_out_f[0][DATA][3] ) );
  HS65_LS_AOI222X2 U424 ( .A(n68), .B(\chs_in_f[2][DATA][3] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][3] ), .E(n52), .F(
        \chs_in_f[1][DATA][3] ), .Z(n364) );
  HS65_LS_OAI212X5 U425 ( .A(n296), .B(n29), .C(n331), .D(n14), .E(n365), .Z(
        \chs_out_f[0][DATA][4] ) );
  HS65_LS_AOI222X2 U426 ( .A(n68), .B(\chs_in_f[2][DATA][4] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][4] ), .E(n52), .F(
        \chs_in_f[1][DATA][4] ), .Z(n365) );
  HS65_LS_OAI212X5 U427 ( .A(n295), .B(n29), .C(n330), .D(n14), .E(n366), .Z(
        \chs_out_f[0][DATA][5] ) );
  HS65_LS_AOI222X2 U428 ( .A(n68), .B(\chs_in_f[2][DATA][5] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][5] ), .E(n52), .F(
        \chs_in_f[1][DATA][5] ), .Z(n366) );
  HS65_LS_OAI212X5 U429 ( .A(n294), .B(n29), .C(n329), .D(n14), .E(n367), .Z(
        \chs_out_f[0][DATA][6] ) );
  HS65_LS_AOI222X2 U430 ( .A(n68), .B(\chs_in_f[2][DATA][6] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][6] ), .E(n52), .F(
        \chs_in_f[1][DATA][6] ), .Z(n367) );
  HS65_LS_OAI212X5 U431 ( .A(n293), .B(n29), .C(n328), .D(n14), .E(n368), .Z(
        \chs_out_f[0][DATA][7] ) );
  HS65_LS_AOI222X2 U432 ( .A(n68), .B(\chs_in_f[2][DATA][7] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][7] ), .E(n52), .F(
        \chs_in_f[1][DATA][7] ), .Z(n368) );
  HS65_LS_OAI212X5 U433 ( .A(n292), .B(n29), .C(n327), .D(n14), .E(n369), .Z(
        \chs_out_f[0][DATA][8] ) );
  HS65_LS_AOI222X2 U434 ( .A(n68), .B(\chs_in_f[2][DATA][8] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][8] ), .E(n52), .F(
        \chs_in_f[1][DATA][8] ), .Z(n369) );
  HS65_LS_OAI212X5 U435 ( .A(n267), .B(n29), .C(n302), .D(n14), .E(n362), .Z(
        \chs_out_f[0][DATA][33] ) );
  HS65_LS_AOI222X2 U436 ( .A(n68), .B(\chs_in_f[2][DATA][33] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][33] ), .E(n52), .F(
        \chs_in_f[1][DATA][33] ), .Z(n362) );
  HS65_LS_OAI212X5 U437 ( .A(n291), .B(n32), .C(n326), .D(n5), .E(n475), .Z(
        \chs_out_f[3][DATA][9] ) );
  HS65_LS_AOI222X2 U438 ( .A(n76), .B(\chs_in_f[2][DATA][9] ), .C(n44), .D(
        \chs_in_f[0][DATA][9] ), .E(n60), .F(\chs_in_f[1][DATA][9] ), .Z(n475)
         );
  HS65_LS_OAI212X5 U439 ( .A(n300), .B(n30), .C(n335), .D(n3), .E(n441), .Z(
        \chs_out_f[3][DATA][0] ) );
  HS65_LS_AOI222X2 U440 ( .A(n74), .B(\chs_in_f[2][DATA][0] ), .C(n42), .D(
        \chs_in_f[0][DATA][0] ), .E(n58), .F(\chs_in_f[1][DATA][0] ), .Z(n441)
         );
  HS65_LS_OAI212X5 U441 ( .A(n299), .B(n30), .C(n334), .D(n3), .E(n452), .Z(
        \chs_out_f[3][DATA][1] ) );
  HS65_LS_AOI222X2 U442 ( .A(n74), .B(\chs_in_f[2][DATA][1] ), .C(n42), .D(
        \chs_in_f[0][DATA][1] ), .E(n58), .F(\chs_in_f[1][DATA][1] ), .Z(n452)
         );
  HS65_LS_OAI212X5 U443 ( .A(n298), .B(n31), .C(n333), .D(n4), .E(n463), .Z(
        \chs_out_f[3][DATA][2] ) );
  HS65_LS_AOI222X2 U444 ( .A(n75), .B(\chs_in_f[2][DATA][2] ), .C(n43), .D(
        \chs_in_f[0][DATA][2] ), .E(n59), .F(\chs_in_f[1][DATA][2] ), .Z(n463)
         );
  HS65_LS_OAI212X5 U445 ( .A(n297), .B(n32), .C(n332), .D(n5), .E(n469), .Z(
        \chs_out_f[3][DATA][3] ) );
  HS65_LS_AOI222X2 U446 ( .A(n76), .B(\chs_in_f[2][DATA][3] ), .C(n44), .D(
        \chs_in_f[0][DATA][3] ), .E(n60), .F(\chs_in_f[1][DATA][3] ), .Z(n469)
         );
  HS65_LS_OAI212X5 U447 ( .A(n296), .B(n32), .C(n331), .D(n5), .E(n470), .Z(
        \chs_out_f[3][DATA][4] ) );
  HS65_LS_AOI222X2 U448 ( .A(n76), .B(\chs_in_f[2][DATA][4] ), .C(n44), .D(
        \chs_in_f[0][DATA][4] ), .E(n60), .F(\chs_in_f[1][DATA][4] ), .Z(n470)
         );
  HS65_LS_OAI212X5 U449 ( .A(n295), .B(n32), .C(n330), .D(n5), .E(n471), .Z(
        \chs_out_f[3][DATA][5] ) );
  HS65_LS_AOI222X2 U450 ( .A(n76), .B(\chs_in_f[2][DATA][5] ), .C(n44), .D(
        \chs_in_f[0][DATA][5] ), .E(n60), .F(\chs_in_f[1][DATA][5] ), .Z(n471)
         );
  HS65_LS_OAI212X5 U451 ( .A(n294), .B(n32), .C(n329), .D(n5), .E(n472), .Z(
        \chs_out_f[3][DATA][6] ) );
  HS65_LS_AOI222X2 U452 ( .A(n76), .B(\chs_in_f[2][DATA][6] ), .C(n44), .D(
        \chs_in_f[0][DATA][6] ), .E(n60), .F(\chs_in_f[1][DATA][6] ), .Z(n472)
         );
  HS65_LS_OAI212X5 U453 ( .A(n293), .B(n32), .C(n328), .D(n5), .E(n473), .Z(
        \chs_out_f[3][DATA][7] ) );
  HS65_LS_AOI222X2 U454 ( .A(n76), .B(\chs_in_f[2][DATA][7] ), .C(n44), .D(
        \chs_in_f[0][DATA][7] ), .E(n60), .F(\chs_in_f[1][DATA][7] ), .Z(n473)
         );
  HS65_LS_OAI212X5 U455 ( .A(n292), .B(n32), .C(n327), .D(n5), .E(n474), .Z(
        \chs_out_f[3][DATA][8] ) );
  HS65_LS_AOI222X2 U456 ( .A(n76), .B(\chs_in_f[2][DATA][8] ), .C(n44), .D(
        \chs_in_f[0][DATA][8] ), .E(n60), .F(\chs_in_f[1][DATA][8] ), .Z(n474)
         );
  HS65_LS_OAI212X5 U457 ( .A(n290), .B(n30), .C(n325), .D(n3), .E(n442), .Z(
        \chs_out_f[3][DATA][10] ) );
  HS65_LS_AOI222X2 U458 ( .A(n74), .B(\chs_in_f[2][DATA][10] ), .C(n42), .D(
        \chs_in_f[0][DATA][10] ), .E(n58), .F(\chs_in_f[1][DATA][10] ), .Z(
        n442) );
  HS65_LS_OAI212X5 U459 ( .A(n289), .B(n30), .C(n324), .D(n3), .E(n443), .Z(
        \chs_out_f[3][DATA][11] ) );
  HS65_LS_AOI222X2 U460 ( .A(n74), .B(\chs_in_f[2][DATA][11] ), .C(n42), .D(
        \chs_in_f[0][DATA][11] ), .E(n58), .F(\chs_in_f[1][DATA][11] ), .Z(
        n443) );
  HS65_LS_OAI212X5 U461 ( .A(n288), .B(n30), .C(n323), .D(n3), .E(n444), .Z(
        \chs_out_f[3][DATA][12] ) );
  HS65_LS_AOI222X2 U462 ( .A(n74), .B(\chs_in_f[2][DATA][12] ), .C(n42), .D(
        \chs_in_f[0][DATA][12] ), .E(n58), .F(\chs_in_f[1][DATA][12] ), .Z(
        n444) );
  HS65_LS_OAI212X5 U463 ( .A(n287), .B(n30), .C(n322), .D(n3), .E(n445), .Z(
        \chs_out_f[3][DATA][13] ) );
  HS65_LS_AOI222X2 U464 ( .A(n74), .B(\chs_in_f[2][DATA][13] ), .C(n42), .D(
        \chs_in_f[0][DATA][13] ), .E(n58), .F(\chs_in_f[1][DATA][13] ), .Z(
        n445) );
  HS65_LS_OAI212X5 U465 ( .A(n286), .B(n30), .C(n321), .D(n3), .E(n446), .Z(
        \chs_out_f[3][DATA][14] ) );
  HS65_LS_AOI222X2 U466 ( .A(n74), .B(\chs_in_f[2][DATA][14] ), .C(n42), .D(
        \chs_in_f[0][DATA][14] ), .E(n58), .F(\chs_in_f[1][DATA][14] ), .Z(
        n446) );
  HS65_LS_OAI212X5 U467 ( .A(n285), .B(n30), .C(n320), .D(n3), .E(n447), .Z(
        \chs_out_f[3][DATA][15] ) );
  HS65_LS_AOI222X2 U468 ( .A(n74), .B(\chs_in_f[2][DATA][15] ), .C(n42), .D(
        \chs_in_f[0][DATA][15] ), .E(n58), .F(\chs_in_f[1][DATA][15] ), .Z(
        n447) );
  HS65_LS_OAI212X5 U469 ( .A(n284), .B(n30), .C(n319), .D(n3), .E(n448), .Z(
        \chs_out_f[3][DATA][16] ) );
  HS65_LS_AOI222X2 U470 ( .A(n74), .B(\chs_in_f[2][DATA][16] ), .C(n42), .D(
        \chs_in_f[0][DATA][16] ), .E(n58), .F(\chs_in_f[1][DATA][16] ), .Z(
        n448) );
  HS65_LS_OAI212X5 U471 ( .A(n283), .B(n30), .C(n318), .D(n3), .E(n449), .Z(
        \chs_out_f[3][DATA][17] ) );
  HS65_LS_AOI222X2 U472 ( .A(n74), .B(\chs_in_f[2][DATA][17] ), .C(n42), .D(
        \chs_in_f[0][DATA][17] ), .E(n58), .F(\chs_in_f[1][DATA][17] ), .Z(
        n449) );
  HS65_LS_OAI212X5 U473 ( .A(n282), .B(n30), .C(n317), .D(n3), .E(n450), .Z(
        \chs_out_f[3][DATA][18] ) );
  HS65_LS_AOI222X2 U474 ( .A(n74), .B(\chs_in_f[2][DATA][18] ), .C(n42), .D(
        \chs_in_f[0][DATA][18] ), .E(n58), .F(\chs_in_f[1][DATA][18] ), .Z(
        n450) );
  HS65_LS_OAI212X5 U475 ( .A(n281), .B(n30), .C(n316), .D(n3), .E(n451), .Z(
        \chs_out_f[3][DATA][19] ) );
  HS65_LS_AOI222X2 U476 ( .A(n74), .B(\chs_in_f[2][DATA][19] ), .C(n42), .D(
        \chs_in_f[0][DATA][19] ), .E(n58), .F(\chs_in_f[1][DATA][19] ), .Z(
        n451) );
  HS65_LS_OAI212X5 U477 ( .A(n280), .B(n30), .C(n315), .D(n4), .E(n453), .Z(
        \chs_out_f[3][DATA][20] ) );
  HS65_LS_AOI222X2 U478 ( .A(n75), .B(\chs_in_f[2][DATA][20] ), .C(n43), .D(
        \chs_in_f[0][DATA][20] ), .E(n59), .F(\chs_in_f[1][DATA][20] ), .Z(
        n453) );
  HS65_LS_OAI212X5 U479 ( .A(n279), .B(n31), .C(n314), .D(n4), .E(n454), .Z(
        \chs_out_f[3][DATA][21] ) );
  HS65_LS_AOI222X2 U480 ( .A(n75), .B(\chs_in_f[2][DATA][21] ), .C(n43), .D(
        \chs_in_f[0][DATA][21] ), .E(n59), .F(\chs_in_f[1][DATA][21] ), .Z(
        n454) );
  HS65_LS_OAI212X5 U481 ( .A(n278), .B(n31), .C(n313), .D(n4), .E(n455), .Z(
        \chs_out_f[3][DATA][22] ) );
  HS65_LS_AOI222X2 U482 ( .A(n75), .B(\chs_in_f[2][DATA][22] ), .C(n43), .D(
        \chs_in_f[0][DATA][22] ), .E(n59), .F(\chs_in_f[1][DATA][22] ), .Z(
        n455) );
  HS65_LS_OAI212X5 U483 ( .A(n277), .B(n31), .C(n312), .D(n4), .E(n456), .Z(
        \chs_out_f[3][DATA][23] ) );
  HS65_LS_AOI222X2 U484 ( .A(n75), .B(\chs_in_f[2][DATA][23] ), .C(n43), .D(
        \chs_in_f[0][DATA][23] ), .E(n59), .F(\chs_in_f[1][DATA][23] ), .Z(
        n456) );
  HS65_LS_OAI212X5 U485 ( .A(n276), .B(n31), .C(n311), .D(n4), .E(n457), .Z(
        \chs_out_f[3][DATA][24] ) );
  HS65_LS_AOI222X2 U486 ( .A(n75), .B(\chs_in_f[2][DATA][24] ), .C(n43), .D(
        \chs_in_f[0][DATA][24] ), .E(n59), .F(\chs_in_f[1][DATA][24] ), .Z(
        n457) );
  HS65_LS_OAI212X5 U487 ( .A(n275), .B(n31), .C(n310), .D(n4), .E(n458), .Z(
        \chs_out_f[3][DATA][25] ) );
  HS65_LS_AOI222X2 U488 ( .A(n75), .B(\chs_in_f[2][DATA][25] ), .C(n43), .D(
        \chs_in_f[0][DATA][25] ), .E(n59), .F(\chs_in_f[1][DATA][25] ), .Z(
        n458) );
  HS65_LS_OAI212X5 U489 ( .A(n274), .B(n31), .C(n309), .D(n4), .E(n459), .Z(
        \chs_out_f[3][DATA][26] ) );
  HS65_LS_AOI222X2 U490 ( .A(n75), .B(\chs_in_f[2][DATA][26] ), .C(n43), .D(
        \chs_in_f[0][DATA][26] ), .E(n59), .F(\chs_in_f[1][DATA][26] ), .Z(
        n459) );
  HS65_LS_OAI212X5 U491 ( .A(n273), .B(n31), .C(n308), .D(n4), .E(n460), .Z(
        \chs_out_f[3][DATA][27] ) );
  HS65_LS_AOI222X2 U492 ( .A(n75), .B(\chs_in_f[2][DATA][27] ), .C(n43), .D(
        \chs_in_f[0][DATA][27] ), .E(n59), .F(\chs_in_f[1][DATA][27] ), .Z(
        n460) );
  HS65_LS_OAI212X5 U493 ( .A(n272), .B(n31), .C(n307), .D(n4), .E(n461), .Z(
        \chs_out_f[3][DATA][28] ) );
  HS65_LS_AOI222X2 U494 ( .A(n75), .B(\chs_in_f[2][DATA][28] ), .C(n43), .D(
        \chs_in_f[0][DATA][28] ), .E(n59), .F(\chs_in_f[1][DATA][28] ), .Z(
        n461) );
  HS65_LS_OAI212X5 U495 ( .A(n271), .B(n31), .C(n306), .D(n4), .E(n462), .Z(
        \chs_out_f[3][DATA][29] ) );
  HS65_LS_AOI222X2 U496 ( .A(n75), .B(\chs_in_f[2][DATA][29] ), .C(n43), .D(
        \chs_in_f[0][DATA][29] ), .E(n59), .F(\chs_in_f[1][DATA][29] ), .Z(
        n462) );
  HS65_LS_OAI212X5 U497 ( .A(n270), .B(n31), .C(n305), .D(n4), .E(n464), .Z(
        \chs_out_f[3][DATA][30] ) );
  HS65_LS_AOI222X2 U498 ( .A(n75), .B(\chs_in_f[2][DATA][30] ), .C(n43), .D(
        \chs_in_f[0][DATA][30] ), .E(n59), .F(\chs_in_f[1][DATA][30] ), .Z(
        n464) );
  HS65_LS_OAI212X5 U499 ( .A(n269), .B(n31), .C(n304), .D(n5), .E(n465), .Z(
        \chs_out_f[3][DATA][31] ) );
  HS65_LS_AOI222X2 U500 ( .A(n76), .B(\chs_in_f[2][DATA][31] ), .C(n44), .D(
        \chs_in_f[0][DATA][31] ), .E(n60), .F(\chs_in_f[1][DATA][31] ), .Z(
        n465) );
  HS65_LS_OAI212X5 U501 ( .A(n268), .B(n31), .C(n303), .D(n5), .E(n466), .Z(
        \chs_out_f[3][DATA][32] ) );
  HS65_LS_AOI222X2 U502 ( .A(n76), .B(\chs_in_f[2][DATA][32] ), .C(n44), .D(
        \chs_in_f[0][DATA][32] ), .E(n60), .F(\chs_in_f[1][DATA][32] ), .Z(
        n466) );
  HS65_LS_OAI212X5 U503 ( .A(n267), .B(n32), .C(n302), .D(n5), .E(n467), .Z(
        \chs_out_f[3][DATA][33] ) );
  HS65_LS_AOI222X2 U504 ( .A(n76), .B(\chs_in_f[2][DATA][33] ), .C(n44), .D(
        \chs_in_f[0][DATA][33] ), .E(n60), .F(\chs_in_f[1][DATA][33] ), .Z(
        n467) );
  HS65_LS_OAI212X5 U505 ( .A(n20), .B(n266), .C(n17), .D(n301), .E(n503), .Z(
        \chs_out_f[4][DATA][34] ) );
  HS65_LS_OAI212X5 U506 ( .A(n266), .B(n32), .C(n301), .D(n5), .E(n468), .Z(
        \chs_out_f[3][DATA][34] ) );
  HS65_LS_OAI212X5 U507 ( .A(n266), .B(n23), .C(n301), .D(n8), .E(n433), .Z(
        \chs_out_f[2][DATA][34] ) );
  HS65_LS_OAI212X5 U508 ( .A(n266), .B(n26), .C(n301), .D(n11), .E(n398), .Z(
        \chs_out_f[1][DATA][34] ) );
  HS65_LS_OAI212X5 U509 ( .A(n266), .B(n29), .C(n301), .D(n14), .E(n363), .Z(
        \chs_out_f[0][DATA][34] ) );
  HS65_LS_IVX9 U510 ( .A(\switch_sel[4][4] ), .Z(n260) );
  HS65_LS_IVX9 U511 ( .A(\switch_sel[3][3] ), .Z(n265) );
endmodule


module latch_controller_0_15 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_0_000000000_15 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, n3, n5, n6, n7, n8, n9, n10;
  assign N0 = preset;

  latch_controller_0_15 controller ( .preset(n6), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLQX9 type_out_reg ( .D(N4), .GN(n8), .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U8 ( .A(\left_in[DATA][34] ), .B(n3), .Z(n9) );
  HS65_LS_AND2X4 U7 ( .A(1'b0), .B(n7), .Z(n10) );
  HS65_LS_OR2X9 U9 ( .A(n10), .B(n9), .Z(N4) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(N39), .Q(\right_out[DATA][33] )
         );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(N38), .Q(\right_out[DATA][32] )
         );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(N37), .Q(\right_out[DATA][31] )
         );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(N36), .Q(\right_out[DATA][30] )
         );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(N35), .Q(\right_out[DATA][29] )
         );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(N34), .Q(\right_out[DATA][28] )
         );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(N33), .Q(\right_out[DATA][27] )
         );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(N32), .Q(\right_out[DATA][26] )
         );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(N31), .Q(\right_out[DATA][25] )
         );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(N30), .Q(\right_out[DATA][24] )
         );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(N29), .Q(\right_out[DATA][23] )
         );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(N28), .Q(\right_out[DATA][22] )
         );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(N27), .Q(\right_out[DATA][21] )
         );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(N26), .Q(\right_out[DATA][20] )
         );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(N25), .Q(\right_out[DATA][19] )
         );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(N24), .Q(\right_out[DATA][18] )
         );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(N23), .Q(\right_out[DATA][17] )
         );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(N22), .Q(\right_out[DATA][16] )
         );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(N21), .Q(\right_out[DATA][15] )
         );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(N20), .Q(\right_out[DATA][14] )
         );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(N19), .Q(\right_out[DATA][13] )
         );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(N18), .Q(\right_out[DATA][12] )
         );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(N17), .Q(\right_out[DATA][11] )
         );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(N16), .Q(\right_out[DATA][10] )
         );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(N15), .Q(\right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(N14), .Q(\right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(N13), .Q(\right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(N12), .Q(\right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(N11), .Q(\right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(N10), .Q(\right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(N9), .Q(\right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(N8), .Q(\right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(N7), .Q(\right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(N6), .Q(\right_out[DATA][0] ) );
  HS65_LS_BFX9 U3 ( .A(N0), .Z(n6) );
  HS65_LS_IVX9 U4 ( .A(n6), .Z(n3) );
  HS65_LS_IVX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_NOR2X6 U6 ( .A(lt_enable), .B(n7), .Z(n8) );
  HS65_LS_AND2X4 U10 ( .A(\left_in[DATA][9] ), .B(n3), .Z(N15) );
  HS65_LS_AND2X4 U11 ( .A(\left_in[DATA][0] ), .B(n3), .Z(N6) );
  HS65_LS_AND2X4 U12 ( .A(\left_in[DATA][1] ), .B(n5), .Z(N7) );
  HS65_LS_AND2X4 U13 ( .A(\left_in[DATA][2] ), .B(n3), .Z(N8) );
  HS65_LS_AND2X4 U14 ( .A(\left_in[DATA][3] ), .B(n5), .Z(N9) );
  HS65_LS_AND2X4 U15 ( .A(\left_in[DATA][4] ), .B(n3), .Z(N10) );
  HS65_LS_AND2X4 U16 ( .A(\left_in[DATA][5] ), .B(n3), .Z(N11) );
  HS65_LS_AND2X4 U17 ( .A(\left_in[DATA][6] ), .B(n3), .Z(N12) );
  HS65_LS_AND2X4 U18 ( .A(\left_in[DATA][7] ), .B(n3), .Z(N13) );
  HS65_LS_AND2X4 U19 ( .A(\left_in[DATA][8] ), .B(n3), .Z(N14) );
  HS65_LS_AND2X4 U20 ( .A(\left_in[DATA][10] ), .B(n3), .Z(N16) );
  HS65_LS_AND2X4 U21 ( .A(\left_in[DATA][11] ), .B(n3), .Z(N17) );
  HS65_LS_AND2X4 U22 ( .A(\left_in[DATA][12] ), .B(n3), .Z(N18) );
  HS65_LS_AND2X4 U23 ( .A(\left_in[DATA][13] ), .B(n3), .Z(N19) );
  HS65_LS_AND2X4 U24 ( .A(\left_in[DATA][14] ), .B(n3), .Z(N20) );
  HS65_LS_AND2X4 U25 ( .A(\left_in[DATA][15] ), .B(n3), .Z(N21) );
  HS65_LS_AND2X4 U26 ( .A(\left_in[DATA][16] ), .B(n3), .Z(N22) );
  HS65_LS_AND2X4 U27 ( .A(\left_in[DATA][17] ), .B(n5), .Z(N23) );
  HS65_LS_AND2X4 U28 ( .A(\left_in[DATA][18] ), .B(n5), .Z(N24) );
  HS65_LS_AND2X4 U29 ( .A(\left_in[DATA][19] ), .B(n5), .Z(N25) );
  HS65_LS_AND2X4 U30 ( .A(\left_in[DATA][20] ), .B(n5), .Z(N26) );
  HS65_LS_AND2X4 U31 ( .A(\left_in[DATA][21] ), .B(n5), .Z(N27) );
  HS65_LS_AND2X4 U32 ( .A(\left_in[DATA][22] ), .B(n5), .Z(N28) );
  HS65_LS_AND2X4 U33 ( .A(\left_in[DATA][23] ), .B(n5), .Z(N29) );
  HS65_LS_AND2X4 U34 ( .A(\left_in[DATA][24] ), .B(n5), .Z(N30) );
  HS65_LS_AND2X4 U35 ( .A(\left_in[DATA][25] ), .B(n5), .Z(N31) );
  HS65_LS_AND2X4 U36 ( .A(\left_in[DATA][26] ), .B(n5), .Z(N32) );
  HS65_LS_AND2X4 U37 ( .A(\left_in[DATA][27] ), .B(n5), .Z(N33) );
  HS65_LS_AND2X4 U38 ( .A(\left_in[DATA][28] ), .B(n5), .Z(N34) );
  HS65_LS_AND2X4 U39 ( .A(\left_in[DATA][29] ), .B(n5), .Z(N35) );
  HS65_LS_AND2X4 U40 ( .A(\left_in[DATA][30] ), .B(n3), .Z(N36) );
  HS65_LS_AND2X4 U41 ( .A(\left_in[DATA][31] ), .B(n5), .Z(N37) );
  HS65_LS_AND2X4 U42 ( .A(\left_in[DATA][32] ), .B(n3), .Z(N38) );
  HS65_LS_AND2X4 U43 ( .A(\left_in[DATA][33] ), .B(n5), .Z(N39) );
  HS65_LS_BFX9 U44 ( .A(N0), .Z(n7) );
  HS65_LS_NAND2X7 U45 ( .A(\right_out[DATA][34] ), .B(n8), .Z(N5) );
endmodule


module latch_controller_0_14 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_0_000000000_14 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, n3, n5, n6, n7, n8, n9, n10;
  assign N0 = preset;

  latch_controller_0_14 controller ( .preset(n6), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLQX9 type_out_reg ( .D(N4), .GN(n8), .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(1'b0), .B(n7), .Z(n10) );
  HS65_LS_OR2X9 U9 ( .A(n10), .B(n9), .Z(N4) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(N39), .Q(\right_out[DATA][33] )
         );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(N38), .Q(\right_out[DATA][32] )
         );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(N37), .Q(\right_out[DATA][31] )
         );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(N36), .Q(\right_out[DATA][30] )
         );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(N35), .Q(\right_out[DATA][29] )
         );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(N34), .Q(\right_out[DATA][28] )
         );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(N33), .Q(\right_out[DATA][27] )
         );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(N32), .Q(\right_out[DATA][26] )
         );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(N31), .Q(\right_out[DATA][25] )
         );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(N30), .Q(\right_out[DATA][24] )
         );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(N29), .Q(\right_out[DATA][23] )
         );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(N28), .Q(\right_out[DATA][22] )
         );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(N27), .Q(\right_out[DATA][21] )
         );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(N26), .Q(\right_out[DATA][20] )
         );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(N25), .Q(\right_out[DATA][19] )
         );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(N24), .Q(\right_out[DATA][18] )
         );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(N23), .Q(\right_out[DATA][17] )
         );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(N22), .Q(\right_out[DATA][16] )
         );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(N21), .Q(\right_out[DATA][15] )
         );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(N20), .Q(\right_out[DATA][14] )
         );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(N19), .Q(\right_out[DATA][13] )
         );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(N18), .Q(\right_out[DATA][12] )
         );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(N17), .Q(\right_out[DATA][11] )
         );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(N16), .Q(\right_out[DATA][10] )
         );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(N15), .Q(\right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(N14), .Q(\right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(N13), .Q(\right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(N12), .Q(\right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(N11), .Q(\right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(N10), .Q(\right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(N9), .Q(\right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(N8), .Q(\right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(N7), .Q(\right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(N6), .Q(\right_out[DATA][0] ) );
  HS65_LS_AND2X4 U8 ( .A(\left_in[DATA][34] ), .B(n5), .Z(n9) );
  HS65_LS_AND2X4 U3 ( .A(\left_in[DATA][3] ), .B(n3), .Z(N9) );
  HS65_LS_AND2X4 U4 ( .A(\left_in[DATA][4] ), .B(n3), .Z(N10) );
  HS65_LS_AND2X4 U5 ( .A(\left_in[DATA][5] ), .B(n3), .Z(N11) );
  HS65_LS_AND2X4 U6 ( .A(\left_in[DATA][6] ), .B(n3), .Z(N12) );
  HS65_LS_AND2X4 U10 ( .A(\left_in[DATA][7] ), .B(n3), .Z(N13) );
  HS65_LS_AND2X4 U11 ( .A(\left_in[DATA][8] ), .B(n3), .Z(N14) );
  HS65_LS_AND2X4 U12 ( .A(\left_in[DATA][9] ), .B(n3), .Z(N15) );
  HS65_LS_AND2X4 U13 ( .A(\left_in[DATA][33] ), .B(n5), .Z(N39) );
  HS65_LS_AND2X4 U14 ( .A(\left_in[DATA][0] ), .B(n3), .Z(N6) );
  HS65_LS_AND2X4 U15 ( .A(\left_in[DATA][1] ), .B(n5), .Z(N7) );
  HS65_LS_AND2X4 U16 ( .A(\left_in[DATA][2] ), .B(n3), .Z(N8) );
  HS65_LS_AND2X4 U17 ( .A(\left_in[DATA][10] ), .B(n3), .Z(N16) );
  HS65_LS_AND2X4 U18 ( .A(\left_in[DATA][11] ), .B(n3), .Z(N17) );
  HS65_LS_AND2X4 U19 ( .A(\left_in[DATA][12] ), .B(n3), .Z(N18) );
  HS65_LS_AND2X4 U20 ( .A(\left_in[DATA][13] ), .B(n3), .Z(N19) );
  HS65_LS_AND2X4 U21 ( .A(\left_in[DATA][14] ), .B(n3), .Z(N20) );
  HS65_LS_AND2X4 U22 ( .A(\left_in[DATA][15] ), .B(n3), .Z(N21) );
  HS65_LS_BFX9 U23 ( .A(N0), .Z(n6) );
  HS65_LS_IVX9 U24 ( .A(n6), .Z(n3) );
  HS65_LS_IVX9 U25 ( .A(n6), .Z(n5) );
  HS65_LS_NOR2X6 U26 ( .A(lt_enable), .B(n7), .Z(n8) );
  HS65_LS_AND2X4 U27 ( .A(\left_in[DATA][16] ), .B(n3), .Z(N22) );
  HS65_LS_AND2X4 U28 ( .A(\left_in[DATA][17] ), .B(n5), .Z(N23) );
  HS65_LS_AND2X4 U29 ( .A(\left_in[DATA][18] ), .B(n5), .Z(N24) );
  HS65_LS_AND2X4 U30 ( .A(\left_in[DATA][19] ), .B(n5), .Z(N25) );
  HS65_LS_AND2X4 U31 ( .A(\left_in[DATA][20] ), .B(n5), .Z(N26) );
  HS65_LS_AND2X4 U32 ( .A(\left_in[DATA][21] ), .B(n5), .Z(N27) );
  HS65_LS_AND2X4 U33 ( .A(\left_in[DATA][22] ), .B(n5), .Z(N28) );
  HS65_LS_AND2X4 U34 ( .A(\left_in[DATA][23] ), .B(n5), .Z(N29) );
  HS65_LS_AND2X4 U35 ( .A(\left_in[DATA][24] ), .B(n5), .Z(N30) );
  HS65_LS_AND2X4 U36 ( .A(\left_in[DATA][25] ), .B(n5), .Z(N31) );
  HS65_LS_AND2X4 U37 ( .A(\left_in[DATA][26] ), .B(n5), .Z(N32) );
  HS65_LS_AND2X4 U38 ( .A(\left_in[DATA][27] ), .B(n5), .Z(N33) );
  HS65_LS_AND2X4 U39 ( .A(\left_in[DATA][28] ), .B(n5), .Z(N34) );
  HS65_LS_AND2X4 U40 ( .A(\left_in[DATA][29] ), .B(n5), .Z(N35) );
  HS65_LS_AND2X4 U41 ( .A(\left_in[DATA][30] ), .B(n3), .Z(N36) );
  HS65_LS_AND2X4 U42 ( .A(\left_in[DATA][31] ), .B(n5), .Z(N37) );
  HS65_LS_AND2X4 U43 ( .A(\left_in[DATA][32] ), .B(n3), .Z(N38) );
  HS65_LS_BFX9 U44 ( .A(N0), .Z(n7) );
  HS65_LS_NAND2X7 U45 ( .A(\right_out[DATA][34] ), .B(n8), .Z(N5) );
endmodule


module latch_controller_0_13 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_0_000000000_13 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, n3, n5, n6, n7, n8, n9, n10;
  assign N0 = preset;

  latch_controller_0_13 controller ( .preset(n6), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLQX9 type_out_reg ( .D(N4), .GN(n8), .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U8 ( .A(\left_in[DATA][34] ), .B(n3), .Z(n9) );
  HS65_LS_AND2X4 U7 ( .A(1'b0), .B(n7), .Z(n10) );
  HS65_LS_OR2X9 U9 ( .A(n10), .B(n9), .Z(N4) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(N39), .Q(\right_out[DATA][33] )
         );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(N38), .Q(\right_out[DATA][32] )
         );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(N37), .Q(\right_out[DATA][31] )
         );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(N36), .Q(\right_out[DATA][30] )
         );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(N35), .Q(\right_out[DATA][29] )
         );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(N34), .Q(\right_out[DATA][28] )
         );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(N33), .Q(\right_out[DATA][27] )
         );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(N32), .Q(\right_out[DATA][26] )
         );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(N31), .Q(\right_out[DATA][25] )
         );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(N30), .Q(\right_out[DATA][24] )
         );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(N29), .Q(\right_out[DATA][23] )
         );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(N28), .Q(\right_out[DATA][22] )
         );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(N27), .Q(\right_out[DATA][21] )
         );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(N26), .Q(\right_out[DATA][20] )
         );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(N25), .Q(\right_out[DATA][19] )
         );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(N24), .Q(\right_out[DATA][18] )
         );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(N23), .Q(\right_out[DATA][17] )
         );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(N22), .Q(\right_out[DATA][16] )
         );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(N21), .Q(\right_out[DATA][15] )
         );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(N20), .Q(\right_out[DATA][14] )
         );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(N19), .Q(\right_out[DATA][13] )
         );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(N18), .Q(\right_out[DATA][12] )
         );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(N17), .Q(\right_out[DATA][11] )
         );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(N16), .Q(\right_out[DATA][10] )
         );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(N15), .Q(\right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(N14), .Q(\right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(N13), .Q(\right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(N12), .Q(\right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(N11), .Q(\right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(N10), .Q(\right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(N9), .Q(\right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(N8), .Q(\right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(N7), .Q(\right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(N6), .Q(\right_out[DATA][0] ) );
  HS65_LS_AND2X4 U3 ( .A(\left_in[DATA][0] ), .B(n3), .Z(N6) );
  HS65_LS_AND2X4 U4 ( .A(\left_in[DATA][1] ), .B(n5), .Z(N7) );
  HS65_LS_AND2X4 U5 ( .A(\left_in[DATA][2] ), .B(n3), .Z(N8) );
  HS65_LS_AND2X4 U6 ( .A(\left_in[DATA][10] ), .B(n3), .Z(N16) );
  HS65_LS_AND2X4 U10 ( .A(\left_in[DATA][11] ), .B(n3), .Z(N17) );
  HS65_LS_AND2X4 U11 ( .A(\left_in[DATA][12] ), .B(n3), .Z(N18) );
  HS65_LS_AND2X4 U12 ( .A(\left_in[DATA][13] ), .B(n3), .Z(N19) );
  HS65_LS_AND2X4 U13 ( .A(\left_in[DATA][14] ), .B(n3), .Z(N20) );
  HS65_LS_AND2X4 U14 ( .A(\left_in[DATA][15] ), .B(n3), .Z(N21) );
  HS65_LS_AND2X4 U15 ( .A(\left_in[DATA][4] ), .B(n3), .Z(N10) );
  HS65_LS_AND2X4 U16 ( .A(\left_in[DATA][5] ), .B(n3), .Z(N11) );
  HS65_LS_AND2X4 U17 ( .A(\left_in[DATA][6] ), .B(n3), .Z(N12) );
  HS65_LS_AND2X4 U18 ( .A(\left_in[DATA][7] ), .B(n3), .Z(N13) );
  HS65_LS_AND2X4 U19 ( .A(\left_in[DATA][8] ), .B(n3), .Z(N14) );
  HS65_LS_AND2X4 U20 ( .A(\left_in[DATA][9] ), .B(n3), .Z(N15) );
  HS65_LS_AND2X4 U21 ( .A(\left_in[DATA][3] ), .B(n5), .Z(N9) );
  HS65_LS_AND2X4 U22 ( .A(\left_in[DATA][33] ), .B(n3), .Z(N39) );
  HS65_LS_BFX9 U23 ( .A(N0), .Z(n6) );
  HS65_LS_IVX9 U24 ( .A(n6), .Z(n3) );
  HS65_LS_IVX9 U25 ( .A(n6), .Z(n5) );
  HS65_LS_NOR2X6 U26 ( .A(lt_enable), .B(n7), .Z(n8) );
  HS65_LS_AND2X4 U27 ( .A(\left_in[DATA][16] ), .B(n3), .Z(N22) );
  HS65_LS_AND2X4 U28 ( .A(\left_in[DATA][17] ), .B(n5), .Z(N23) );
  HS65_LS_AND2X4 U29 ( .A(\left_in[DATA][18] ), .B(n5), .Z(N24) );
  HS65_LS_AND2X4 U30 ( .A(\left_in[DATA][19] ), .B(n5), .Z(N25) );
  HS65_LS_AND2X4 U31 ( .A(\left_in[DATA][20] ), .B(n5), .Z(N26) );
  HS65_LS_AND2X4 U32 ( .A(\left_in[DATA][21] ), .B(n5), .Z(N27) );
  HS65_LS_AND2X4 U33 ( .A(\left_in[DATA][22] ), .B(n5), .Z(N28) );
  HS65_LS_AND2X4 U34 ( .A(\left_in[DATA][23] ), .B(n5), .Z(N29) );
  HS65_LS_AND2X4 U35 ( .A(\left_in[DATA][24] ), .B(n5), .Z(N30) );
  HS65_LS_AND2X4 U36 ( .A(\left_in[DATA][25] ), .B(n5), .Z(N31) );
  HS65_LS_AND2X4 U37 ( .A(\left_in[DATA][26] ), .B(n5), .Z(N32) );
  HS65_LS_AND2X4 U38 ( .A(\left_in[DATA][27] ), .B(n5), .Z(N33) );
  HS65_LS_AND2X4 U39 ( .A(\left_in[DATA][28] ), .B(n5), .Z(N34) );
  HS65_LS_AND2X4 U40 ( .A(\left_in[DATA][29] ), .B(n5), .Z(N35) );
  HS65_LS_AND2X4 U41 ( .A(\left_in[DATA][30] ), .B(n5), .Z(N36) );
  HS65_LS_AND2X4 U42 ( .A(\left_in[DATA][31] ), .B(n3), .Z(N37) );
  HS65_LS_AND2X4 U43 ( .A(\left_in[DATA][32] ), .B(n5), .Z(N38) );
  HS65_LS_BFX9 U44 ( .A(N0), .Z(n7) );
  HS65_LS_NAND2X7 U45 ( .A(\right_out[DATA][34] ), .B(n8), .Z(N5) );
endmodule


module latch_controller_0_12 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_0_000000000_12 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, n3, n5, n6, n7, n8, n9, n10;
  assign N0 = preset;

  latch_controller_0_12 controller ( .preset(n6), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLQX9 type_out_reg ( .D(N4), .GN(n8), .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U8 ( .A(\left_in[DATA][34] ), .B(n3), .Z(n9) );
  HS65_LS_AND2X4 U7 ( .A(1'b0), .B(n7), .Z(n10) );
  HS65_LS_OR2X9 U9 ( .A(n10), .B(n9), .Z(N4) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(N39), .Q(\right_out[DATA][33] )
         );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(N38), .Q(\right_out[DATA][32] )
         );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(N37), .Q(\right_out[DATA][31] )
         );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(N36), .Q(\right_out[DATA][30] )
         );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(N35), .Q(\right_out[DATA][29] )
         );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(N34), .Q(\right_out[DATA][28] )
         );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(N33), .Q(\right_out[DATA][27] )
         );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(N32), .Q(\right_out[DATA][26] )
         );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(N31), .Q(\right_out[DATA][25] )
         );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(N30), .Q(\right_out[DATA][24] )
         );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(N29), .Q(\right_out[DATA][23] )
         );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(N28), .Q(\right_out[DATA][22] )
         );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(N27), .Q(\right_out[DATA][21] )
         );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(N26), .Q(\right_out[DATA][20] )
         );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(N25), .Q(\right_out[DATA][19] )
         );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(N24), .Q(\right_out[DATA][18] )
         );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(N23), .Q(\right_out[DATA][17] )
         );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(N22), .Q(\right_out[DATA][16] )
         );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(N21), .Q(\right_out[DATA][15] )
         );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(N20), .Q(\right_out[DATA][14] )
         );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(N19), .Q(\right_out[DATA][13] )
         );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(N18), .Q(\right_out[DATA][12] )
         );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(N17), .Q(\right_out[DATA][11] )
         );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(N16), .Q(\right_out[DATA][10] )
         );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(N15), .Q(\right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(N14), .Q(\right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(N13), .Q(\right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(N12), .Q(\right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(N11), .Q(\right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(N10), .Q(\right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(N9), .Q(\right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(N8), .Q(\right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(N7), .Q(\right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(N6), .Q(\right_out[DATA][0] ) );
  HS65_LS_AND2X4 U3 ( .A(\left_in[DATA][0] ), .B(n3), .Z(N6) );
  HS65_LS_AND2X4 U4 ( .A(\left_in[DATA][1] ), .B(n5), .Z(N7) );
  HS65_LS_AND2X4 U5 ( .A(\left_in[DATA][2] ), .B(n3), .Z(N8) );
  HS65_LS_AND2X4 U6 ( .A(\left_in[DATA][10] ), .B(n3), .Z(N16) );
  HS65_LS_AND2X4 U10 ( .A(\left_in[DATA][11] ), .B(n3), .Z(N17) );
  HS65_LS_AND2X4 U11 ( .A(\left_in[DATA][12] ), .B(n3), .Z(N18) );
  HS65_LS_AND2X4 U12 ( .A(\left_in[DATA][13] ), .B(n3), .Z(N19) );
  HS65_LS_AND2X4 U13 ( .A(\left_in[DATA][14] ), .B(n3), .Z(N20) );
  HS65_LS_AND2X4 U14 ( .A(\left_in[DATA][15] ), .B(n3), .Z(N21) );
  HS65_LS_AND2X4 U15 ( .A(\left_in[DATA][4] ), .B(n3), .Z(N10) );
  HS65_LS_AND2X4 U16 ( .A(\left_in[DATA][5] ), .B(n3), .Z(N11) );
  HS65_LS_AND2X4 U17 ( .A(\left_in[DATA][6] ), .B(n3), .Z(N12) );
  HS65_LS_AND2X4 U18 ( .A(\left_in[DATA][7] ), .B(n3), .Z(N13) );
  HS65_LS_AND2X4 U19 ( .A(\left_in[DATA][8] ), .B(n3), .Z(N14) );
  HS65_LS_AND2X4 U20 ( .A(\left_in[DATA][9] ), .B(n3), .Z(N15) );
  HS65_LS_AND2X4 U21 ( .A(\left_in[DATA][3] ), .B(n5), .Z(N9) );
  HS65_LS_AND2X4 U22 ( .A(\left_in[DATA][33] ), .B(n3), .Z(N39) );
  HS65_LS_BFX9 U23 ( .A(N0), .Z(n6) );
  HS65_LS_IVX9 U24 ( .A(n6), .Z(n3) );
  HS65_LS_IVX9 U25 ( .A(n6), .Z(n5) );
  HS65_LS_NOR2X6 U26 ( .A(lt_enable), .B(n7), .Z(n8) );
  HS65_LS_AND2X4 U27 ( .A(\left_in[DATA][16] ), .B(n3), .Z(N22) );
  HS65_LS_AND2X4 U28 ( .A(\left_in[DATA][17] ), .B(n5), .Z(N23) );
  HS65_LS_AND2X4 U29 ( .A(\left_in[DATA][18] ), .B(n5), .Z(N24) );
  HS65_LS_AND2X4 U30 ( .A(\left_in[DATA][19] ), .B(n5), .Z(N25) );
  HS65_LS_AND2X4 U31 ( .A(\left_in[DATA][20] ), .B(n5), .Z(N26) );
  HS65_LS_AND2X4 U32 ( .A(\left_in[DATA][21] ), .B(n5), .Z(N27) );
  HS65_LS_AND2X4 U33 ( .A(\left_in[DATA][22] ), .B(n5), .Z(N28) );
  HS65_LS_AND2X4 U34 ( .A(\left_in[DATA][23] ), .B(n5), .Z(N29) );
  HS65_LS_AND2X4 U35 ( .A(\left_in[DATA][24] ), .B(n5), .Z(N30) );
  HS65_LS_AND2X4 U36 ( .A(\left_in[DATA][25] ), .B(n5), .Z(N31) );
  HS65_LS_AND2X4 U37 ( .A(\left_in[DATA][26] ), .B(n5), .Z(N32) );
  HS65_LS_AND2X4 U38 ( .A(\left_in[DATA][27] ), .B(n5), .Z(N33) );
  HS65_LS_AND2X4 U39 ( .A(\left_in[DATA][28] ), .B(n5), .Z(N34) );
  HS65_LS_AND2X4 U40 ( .A(\left_in[DATA][29] ), .B(n5), .Z(N35) );
  HS65_LS_AND2X4 U41 ( .A(\left_in[DATA][30] ), .B(n5), .Z(N36) );
  HS65_LS_AND2X4 U42 ( .A(\left_in[DATA][31] ), .B(n3), .Z(N37) );
  HS65_LS_AND2X4 U43 ( .A(\left_in[DATA][32] ), .B(n5), .Z(N38) );
  HS65_LS_BFX9 U44 ( .A(N0), .Z(n7) );
  HS65_LS_NAND2X7 U45 ( .A(\right_out[DATA][34] ), .B(n8), .Z(N5) );
endmodule


module latch_controller_0_11 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_0_000000000_11 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, n3, n5, n6, n7, n8, n9, n10;
  assign N0 = preset;

  latch_controller_0_11 controller ( .preset(n6), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLQX9 type_out_reg ( .D(N4), .GN(n8), .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U8 ( .A(\left_in[DATA][34] ), .B(n3), .Z(n9) );
  HS65_LS_AND2X4 U7 ( .A(1'b0), .B(n7), .Z(n10) );
  HS65_LS_OR2X9 U9 ( .A(n10), .B(n9), .Z(N4) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(N39), .Q(\right_out[DATA][33] )
         );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(N38), .Q(\right_out[DATA][32] )
         );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(N37), .Q(\right_out[DATA][31] )
         );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(N36), .Q(\right_out[DATA][30] )
         );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(N35), .Q(\right_out[DATA][29] )
         );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(N34), .Q(\right_out[DATA][28] )
         );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(N33), .Q(\right_out[DATA][27] )
         );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(N32), .Q(\right_out[DATA][26] )
         );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(N31), .Q(\right_out[DATA][25] )
         );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(N30), .Q(\right_out[DATA][24] )
         );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(N29), .Q(\right_out[DATA][23] )
         );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(N28), .Q(\right_out[DATA][22] )
         );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(N27), .Q(\right_out[DATA][21] )
         );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(N26), .Q(\right_out[DATA][20] )
         );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(N25), .Q(\right_out[DATA][19] )
         );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(N24), .Q(\right_out[DATA][18] )
         );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(N23), .Q(\right_out[DATA][17] )
         );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(N22), .Q(\right_out[DATA][16] )
         );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(N21), .Q(\right_out[DATA][15] )
         );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(N20), .Q(\right_out[DATA][14] )
         );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(N19), .Q(\right_out[DATA][13] )
         );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(N18), .Q(\right_out[DATA][12] )
         );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(N17), .Q(\right_out[DATA][11] )
         );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(N16), .Q(\right_out[DATA][10] )
         );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(N15), .Q(\right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(N14), .Q(\right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(N13), .Q(\right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(N12), .Q(\right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(N11), .Q(\right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(N10), .Q(\right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(N9), .Q(\right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(N8), .Q(\right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(N7), .Q(\right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(N6), .Q(\right_out[DATA][0] ) );
  HS65_LS_AND2X4 U3 ( .A(\left_in[DATA][4] ), .B(n3), .Z(N10) );
  HS65_LS_AND2X4 U4 ( .A(\left_in[DATA][5] ), .B(n3), .Z(N11) );
  HS65_LS_AND2X4 U5 ( .A(\left_in[DATA][6] ), .B(n3), .Z(N12) );
  HS65_LS_AND2X4 U6 ( .A(\left_in[DATA][7] ), .B(n3), .Z(N13) );
  HS65_LS_AND2X4 U10 ( .A(\left_in[DATA][8] ), .B(n3), .Z(N14) );
  HS65_LS_AND2X4 U11 ( .A(\left_in[DATA][9] ), .B(n3), .Z(N15) );
  HS65_LS_AND2X4 U12 ( .A(\left_in[DATA][10] ), .B(n3), .Z(N16) );
  HS65_LS_AND2X4 U13 ( .A(\left_in[DATA][11] ), .B(n3), .Z(N17) );
  HS65_LS_AND2X4 U14 ( .A(\left_in[DATA][12] ), .B(n3), .Z(N18) );
  HS65_LS_AND2X4 U15 ( .A(\left_in[DATA][13] ), .B(n3), .Z(N19) );
  HS65_LS_AND2X4 U16 ( .A(\left_in[DATA][14] ), .B(n3), .Z(N20) );
  HS65_LS_AND2X4 U17 ( .A(\left_in[DATA][15] ), .B(n3), .Z(N21) );
  HS65_LS_AND2X4 U18 ( .A(\left_in[DATA][0] ), .B(n3), .Z(N6) );
  HS65_LS_AND2X4 U19 ( .A(\left_in[DATA][1] ), .B(n5), .Z(N7) );
  HS65_LS_AND2X4 U20 ( .A(\left_in[DATA][2] ), .B(n3), .Z(N8) );
  HS65_LS_AND2X4 U21 ( .A(\left_in[DATA][3] ), .B(n5), .Z(N9) );
  HS65_LS_AND2X4 U22 ( .A(\left_in[DATA][33] ), .B(n3), .Z(N39) );
  HS65_LS_BFX9 U23 ( .A(N0), .Z(n6) );
  HS65_LS_IVX9 U24 ( .A(n6), .Z(n3) );
  HS65_LS_IVX9 U25 ( .A(n6), .Z(n5) );
  HS65_LS_NOR2X6 U26 ( .A(lt_enable), .B(n7), .Z(n8) );
  HS65_LS_AND2X4 U27 ( .A(\left_in[DATA][16] ), .B(n3), .Z(N22) );
  HS65_LS_AND2X4 U28 ( .A(\left_in[DATA][17] ), .B(n5), .Z(N23) );
  HS65_LS_AND2X4 U29 ( .A(\left_in[DATA][18] ), .B(n5), .Z(N24) );
  HS65_LS_AND2X4 U30 ( .A(\left_in[DATA][19] ), .B(n5), .Z(N25) );
  HS65_LS_AND2X4 U31 ( .A(\left_in[DATA][20] ), .B(n5), .Z(N26) );
  HS65_LS_AND2X4 U32 ( .A(\left_in[DATA][21] ), .B(n5), .Z(N27) );
  HS65_LS_AND2X4 U33 ( .A(\left_in[DATA][22] ), .B(n5), .Z(N28) );
  HS65_LS_AND2X4 U34 ( .A(\left_in[DATA][23] ), .B(n5), .Z(N29) );
  HS65_LS_AND2X4 U35 ( .A(\left_in[DATA][24] ), .B(n5), .Z(N30) );
  HS65_LS_AND2X4 U36 ( .A(\left_in[DATA][25] ), .B(n5), .Z(N31) );
  HS65_LS_AND2X4 U37 ( .A(\left_in[DATA][26] ), .B(n5), .Z(N32) );
  HS65_LS_AND2X4 U38 ( .A(\left_in[DATA][27] ), .B(n5), .Z(N33) );
  HS65_LS_AND2X4 U39 ( .A(\left_in[DATA][28] ), .B(n5), .Z(N34) );
  HS65_LS_AND2X4 U40 ( .A(\left_in[DATA][29] ), .B(n5), .Z(N35) );
  HS65_LS_AND2X4 U41 ( .A(\left_in[DATA][30] ), .B(n5), .Z(N36) );
  HS65_LS_AND2X4 U42 ( .A(\left_in[DATA][31] ), .B(n3), .Z(N37) );
  HS65_LS_AND2X4 U43 ( .A(\left_in[DATA][32] ), .B(n5), .Z(N38) );
  HS65_LS_BFX9 U44 ( .A(N0), .Z(n7) );
  HS65_LS_NAND2X7 U45 ( .A(\right_out[DATA][34] ), .B(n8), .Z(N5) );
endmodule


module crossbar_stage_3 ( preset, .switch_sel({\switch_sel[4][4] , 
        \switch_sel[4][3] , \switch_sel[4][2] , \switch_sel[4][1] , 
        \switch_sel[4][0] , \switch_sel[3][4] , \switch_sel[3][3] , 
        \switch_sel[3][2] , \switch_sel[3][1] , \switch_sel[3][0] , 
        \switch_sel[2][4] , \switch_sel[2][3] , \switch_sel[2][2] , 
        \switch_sel[2][1] , \switch_sel[2][0] , \switch_sel[1][4] , 
        \switch_sel[1][3] , \switch_sel[1][2] , \switch_sel[1][1] , 
        \switch_sel[1][0] , \switch_sel[0][4] , \switch_sel[0][3] , 
        \switch_sel[0][2] , \switch_sel[0][1] , \switch_sel[0][0] }), 
    .chs_in_f({\chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] , 
        \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] , 
        \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] , 
        \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] , 
        \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] , 
        \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] , 
        \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] , 
        \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] , 
        \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] , 
        \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] , 
        \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] , 
        \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] , 
        \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] , 
        \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] , \chs_in_f[4][DATA][7] , 
        \chs_in_f[4][DATA][6] , \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] , 
        \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] , \chs_in_f[4][DATA][1] , 
        \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] , \chs_in_f[3][DATA][34] , 
        \chs_in_f[3][DATA][33] , \chs_in_f[3][DATA][32] , 
        \chs_in_f[3][DATA][31] , \chs_in_f[3][DATA][30] , 
        \chs_in_f[3][DATA][29] , \chs_in_f[3][DATA][28] , 
        \chs_in_f[3][DATA][27] , \chs_in_f[3][DATA][26] , 
        \chs_in_f[3][DATA][25] , \chs_in_f[3][DATA][24] , 
        \chs_in_f[3][DATA][23] , \chs_in_f[3][DATA][22] , 
        \chs_in_f[3][DATA][21] , \chs_in_f[3][DATA][20] , 
        \chs_in_f[3][DATA][19] , \chs_in_f[3][DATA][18] , 
        \chs_in_f[3][DATA][17] , \chs_in_f[3][DATA][16] , 
        \chs_in_f[3][DATA][15] , \chs_in_f[3][DATA][14] , 
        \chs_in_f[3][DATA][13] , \chs_in_f[3][DATA][12] , 
        \chs_in_f[3][DATA][11] , \chs_in_f[3][DATA][10] , 
        \chs_in_f[3][DATA][9] , \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] , 
        \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] , \chs_in_f[3][DATA][4] , 
        \chs_in_f[3][DATA][3] , \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] , 
        \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] , 
        \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] , 
        \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] , 
        \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] , 
        \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] , 
        \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] , 
        \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] , 
        \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] , 
        \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] , 
        \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] , 
        \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] , 
        \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] , 
        \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] , 
        \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] , \chs_in_f[2][DATA][7] , 
        \chs_in_f[2][DATA][6] , \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] , 
        \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] , \chs_in_f[2][DATA][1] , 
        \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] , \chs_in_f[1][DATA][34] , 
        \chs_in_f[1][DATA][33] , \chs_in_f[1][DATA][32] , 
        \chs_in_f[1][DATA][31] , \chs_in_f[1][DATA][30] , 
        \chs_in_f[1][DATA][29] , \chs_in_f[1][DATA][28] , 
        \chs_in_f[1][DATA][27] , \chs_in_f[1][DATA][26] , 
        \chs_in_f[1][DATA][25] , \chs_in_f[1][DATA][24] , 
        \chs_in_f[1][DATA][23] , \chs_in_f[1][DATA][22] , 
        \chs_in_f[1][DATA][21] , \chs_in_f[1][DATA][20] , 
        \chs_in_f[1][DATA][19] , \chs_in_f[1][DATA][18] , 
        \chs_in_f[1][DATA][17] , \chs_in_f[1][DATA][16] , 
        \chs_in_f[1][DATA][15] , \chs_in_f[1][DATA][14] , 
        \chs_in_f[1][DATA][13] , \chs_in_f[1][DATA][12] , 
        \chs_in_f[1][DATA][11] , \chs_in_f[1][DATA][10] , 
        \chs_in_f[1][DATA][9] , \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] , 
        \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] , \chs_in_f[1][DATA][4] , 
        \chs_in_f[1][DATA][3] , \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] , 
        \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] , 
        \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] , 
        \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] , 
        \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] , 
        \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] , 
        \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] , 
        \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] , 
        \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] , 
        \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] , 
        \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] , 
        \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] , 
        \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] , 
        \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] , 
        \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] , \chs_in_f[0][DATA][7] , 
        \chs_in_f[0][DATA][6] , \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] , 
        \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] , \chs_in_f[0][DATA][1] , 
        \chs_in_f[0][DATA][0] }), .chs_in_b({\chs_in_b[4][ACK] , 
        \chs_in_b[3][ACK] , \chs_in_b[2][ACK] , \chs_in_b[1][ACK] , 
        \chs_in_b[0][ACK] }), .latches_out_f({\latches_out_f[4][REQ] , 
        \latches_out_f[4][DATA][34] , \latches_out_f[4][DATA][33] , 
        \latches_out_f[4][DATA][32] , \latches_out_f[4][DATA][31] , 
        \latches_out_f[4][DATA][30] , \latches_out_f[4][DATA][29] , 
        \latches_out_f[4][DATA][28] , \latches_out_f[4][DATA][27] , 
        \latches_out_f[4][DATA][26] , \latches_out_f[4][DATA][25] , 
        \latches_out_f[4][DATA][24] , \latches_out_f[4][DATA][23] , 
        \latches_out_f[4][DATA][22] , \latches_out_f[4][DATA][21] , 
        \latches_out_f[4][DATA][20] , \latches_out_f[4][DATA][19] , 
        \latches_out_f[4][DATA][18] , \latches_out_f[4][DATA][17] , 
        \latches_out_f[4][DATA][16] , \latches_out_f[4][DATA][15] , 
        \latches_out_f[4][DATA][14] , \latches_out_f[4][DATA][13] , 
        \latches_out_f[4][DATA][12] , \latches_out_f[4][DATA][11] , 
        \latches_out_f[4][DATA][10] , \latches_out_f[4][DATA][9] , 
        \latches_out_f[4][DATA][8] , \latches_out_f[4][DATA][7] , 
        \latches_out_f[4][DATA][6] , \latches_out_f[4][DATA][5] , 
        \latches_out_f[4][DATA][4] , \latches_out_f[4][DATA][3] , 
        \latches_out_f[4][DATA][2] , \latches_out_f[4][DATA][1] , 
        \latches_out_f[4][DATA][0] , \latches_out_f[3][REQ] , 
        \latches_out_f[3][DATA][34] , \latches_out_f[3][DATA][33] , 
        \latches_out_f[3][DATA][32] , \latches_out_f[3][DATA][31] , 
        \latches_out_f[3][DATA][30] , \latches_out_f[3][DATA][29] , 
        \latches_out_f[3][DATA][28] , \latches_out_f[3][DATA][27] , 
        \latches_out_f[3][DATA][26] , \latches_out_f[3][DATA][25] , 
        \latches_out_f[3][DATA][24] , \latches_out_f[3][DATA][23] , 
        \latches_out_f[3][DATA][22] , \latches_out_f[3][DATA][21] , 
        \latches_out_f[3][DATA][20] , \latches_out_f[3][DATA][19] , 
        \latches_out_f[3][DATA][18] , \latches_out_f[3][DATA][17] , 
        \latches_out_f[3][DATA][16] , \latches_out_f[3][DATA][15] , 
        \latches_out_f[3][DATA][14] , \latches_out_f[3][DATA][13] , 
        \latches_out_f[3][DATA][12] , \latches_out_f[3][DATA][11] , 
        \latches_out_f[3][DATA][10] , \latches_out_f[3][DATA][9] , 
        \latches_out_f[3][DATA][8] , \latches_out_f[3][DATA][7] , 
        \latches_out_f[3][DATA][6] , \latches_out_f[3][DATA][5] , 
        \latches_out_f[3][DATA][4] , \latches_out_f[3][DATA][3] , 
        \latches_out_f[3][DATA][2] , \latches_out_f[3][DATA][1] , 
        \latches_out_f[3][DATA][0] , \latches_out_f[2][REQ] , 
        \latches_out_f[2][DATA][34] , \latches_out_f[2][DATA][33] , 
        \latches_out_f[2][DATA][32] , \latches_out_f[2][DATA][31] , 
        \latches_out_f[2][DATA][30] , \latches_out_f[2][DATA][29] , 
        \latches_out_f[2][DATA][28] , \latches_out_f[2][DATA][27] , 
        \latches_out_f[2][DATA][26] , \latches_out_f[2][DATA][25] , 
        \latches_out_f[2][DATA][24] , \latches_out_f[2][DATA][23] , 
        \latches_out_f[2][DATA][22] , \latches_out_f[2][DATA][21] , 
        \latches_out_f[2][DATA][20] , \latches_out_f[2][DATA][19] , 
        \latches_out_f[2][DATA][18] , \latches_out_f[2][DATA][17] , 
        \latches_out_f[2][DATA][16] , \latches_out_f[2][DATA][15] , 
        \latches_out_f[2][DATA][14] , \latches_out_f[2][DATA][13] , 
        \latches_out_f[2][DATA][12] , \latches_out_f[2][DATA][11] , 
        \latches_out_f[2][DATA][10] , \latches_out_f[2][DATA][9] , 
        \latches_out_f[2][DATA][8] , \latches_out_f[2][DATA][7] , 
        \latches_out_f[2][DATA][6] , \latches_out_f[2][DATA][5] , 
        \latches_out_f[2][DATA][4] , \latches_out_f[2][DATA][3] , 
        \latches_out_f[2][DATA][2] , \latches_out_f[2][DATA][1] , 
        \latches_out_f[2][DATA][0] , \latches_out_f[1][REQ] , 
        \latches_out_f[1][DATA][34] , \latches_out_f[1][DATA][33] , 
        \latches_out_f[1][DATA][32] , \latches_out_f[1][DATA][31] , 
        \latches_out_f[1][DATA][30] , \latches_out_f[1][DATA][29] , 
        \latches_out_f[1][DATA][28] , \latches_out_f[1][DATA][27] , 
        \latches_out_f[1][DATA][26] , \latches_out_f[1][DATA][25] , 
        \latches_out_f[1][DATA][24] , \latches_out_f[1][DATA][23] , 
        \latches_out_f[1][DATA][22] , \latches_out_f[1][DATA][21] , 
        \latches_out_f[1][DATA][20] , \latches_out_f[1][DATA][19] , 
        \latches_out_f[1][DATA][18] , \latches_out_f[1][DATA][17] , 
        \latches_out_f[1][DATA][16] , \latches_out_f[1][DATA][15] , 
        \latches_out_f[1][DATA][14] , \latches_out_f[1][DATA][13] , 
        \latches_out_f[1][DATA][12] , \latches_out_f[1][DATA][11] , 
        \latches_out_f[1][DATA][10] , \latches_out_f[1][DATA][9] , 
        \latches_out_f[1][DATA][8] , \latches_out_f[1][DATA][7] , 
        \latches_out_f[1][DATA][6] , \latches_out_f[1][DATA][5] , 
        \latches_out_f[1][DATA][4] , \latches_out_f[1][DATA][3] , 
        \latches_out_f[1][DATA][2] , \latches_out_f[1][DATA][1] , 
        \latches_out_f[1][DATA][0] , \latches_out_f[0][REQ] , 
        \latches_out_f[0][DATA][34] , \latches_out_f[0][DATA][33] , 
        \latches_out_f[0][DATA][32] , \latches_out_f[0][DATA][31] , 
        \latches_out_f[0][DATA][30] , \latches_out_f[0][DATA][29] , 
        \latches_out_f[0][DATA][28] , \latches_out_f[0][DATA][27] , 
        \latches_out_f[0][DATA][26] , \latches_out_f[0][DATA][25] , 
        \latches_out_f[0][DATA][24] , \latches_out_f[0][DATA][23] , 
        \latches_out_f[0][DATA][22] , \latches_out_f[0][DATA][21] , 
        \latches_out_f[0][DATA][20] , \latches_out_f[0][DATA][19] , 
        \latches_out_f[0][DATA][18] , \latches_out_f[0][DATA][17] , 
        \latches_out_f[0][DATA][16] , \latches_out_f[0][DATA][15] , 
        \latches_out_f[0][DATA][14] , \latches_out_f[0][DATA][13] , 
        \latches_out_f[0][DATA][12] , \latches_out_f[0][DATA][11] , 
        \latches_out_f[0][DATA][10] , \latches_out_f[0][DATA][9] , 
        \latches_out_f[0][DATA][8] , \latches_out_f[0][DATA][7] , 
        \latches_out_f[0][DATA][6] , \latches_out_f[0][DATA][5] , 
        \latches_out_f[0][DATA][4] , \latches_out_f[0][DATA][3] , 
        \latches_out_f[0][DATA][2] , \latches_out_f[0][DATA][1] , 
        \latches_out_f[0][DATA][0] }), .latches_out_b({\latches_out_b[4][ACK] , 
        \latches_out_b[3][ACK] , \latches_out_b[2][ACK] , 
        \latches_out_b[1][ACK] , \latches_out_b[0][ACK] }) );
  input preset, \switch_sel[4][4] , \switch_sel[4][3] , \switch_sel[4][2] ,
         \switch_sel[4][1] , \switch_sel[4][0] , \switch_sel[3][4] ,
         \switch_sel[3][3] , \switch_sel[3][2] , \switch_sel[3][1] ,
         \switch_sel[3][0] , \switch_sel[2][4] , \switch_sel[2][3] ,
         \switch_sel[2][2] , \switch_sel[2][1] , \switch_sel[2][0] ,
         \switch_sel[1][4] , \switch_sel[1][3] , \switch_sel[1][2] ,
         \switch_sel[1][1] , \switch_sel[1][0] , \switch_sel[0][4] ,
         \switch_sel[0][3] , \switch_sel[0][2] , \switch_sel[0][1] ,
         \switch_sel[0][0] , \chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] ,
         \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] ,
         \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] ,
         \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] ,
         \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] ,
         \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] ,
         \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] ,
         \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] ,
         \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] ,
         \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] ,
         \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] ,
         \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] ,
         \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] ,
         \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] ,
         \chs_in_f[4][DATA][7] , \chs_in_f[4][DATA][6] ,
         \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] ,
         \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] ,
         \chs_in_f[4][DATA][1] , \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] ,
         \chs_in_f[3][DATA][34] , \chs_in_f[3][DATA][33] ,
         \chs_in_f[3][DATA][32] , \chs_in_f[3][DATA][31] ,
         \chs_in_f[3][DATA][30] , \chs_in_f[3][DATA][29] ,
         \chs_in_f[3][DATA][28] , \chs_in_f[3][DATA][27] ,
         \chs_in_f[3][DATA][26] , \chs_in_f[3][DATA][25] ,
         \chs_in_f[3][DATA][24] , \chs_in_f[3][DATA][23] ,
         \chs_in_f[3][DATA][22] , \chs_in_f[3][DATA][21] ,
         \chs_in_f[3][DATA][20] , \chs_in_f[3][DATA][19] ,
         \chs_in_f[3][DATA][18] , \chs_in_f[3][DATA][17] ,
         \chs_in_f[3][DATA][16] , \chs_in_f[3][DATA][15] ,
         \chs_in_f[3][DATA][14] , \chs_in_f[3][DATA][13] ,
         \chs_in_f[3][DATA][12] , \chs_in_f[3][DATA][11] ,
         \chs_in_f[3][DATA][10] , \chs_in_f[3][DATA][9] ,
         \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] ,
         \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] ,
         \chs_in_f[3][DATA][4] , \chs_in_f[3][DATA][3] ,
         \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] ,
         \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] ,
         \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] ,
         \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] ,
         \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] ,
         \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] ,
         \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] ,
         \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] ,
         \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] ,
         \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] ,
         \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] ,
         \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] ,
         \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] ,
         \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] ,
         \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] ,
         \chs_in_f[2][DATA][7] , \chs_in_f[2][DATA][6] ,
         \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] ,
         \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] ,
         \chs_in_f[2][DATA][1] , \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] ,
         \chs_in_f[1][DATA][34] , \chs_in_f[1][DATA][33] ,
         \chs_in_f[1][DATA][32] , \chs_in_f[1][DATA][31] ,
         \chs_in_f[1][DATA][30] , \chs_in_f[1][DATA][29] ,
         \chs_in_f[1][DATA][28] , \chs_in_f[1][DATA][27] ,
         \chs_in_f[1][DATA][26] , \chs_in_f[1][DATA][25] ,
         \chs_in_f[1][DATA][24] , \chs_in_f[1][DATA][23] ,
         \chs_in_f[1][DATA][22] , \chs_in_f[1][DATA][21] ,
         \chs_in_f[1][DATA][20] , \chs_in_f[1][DATA][19] ,
         \chs_in_f[1][DATA][18] , \chs_in_f[1][DATA][17] ,
         \chs_in_f[1][DATA][16] , \chs_in_f[1][DATA][15] ,
         \chs_in_f[1][DATA][14] , \chs_in_f[1][DATA][13] ,
         \chs_in_f[1][DATA][12] , \chs_in_f[1][DATA][11] ,
         \chs_in_f[1][DATA][10] , \chs_in_f[1][DATA][9] ,
         \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] ,
         \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] ,
         \chs_in_f[1][DATA][4] , \chs_in_f[1][DATA][3] ,
         \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] ,
         \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] ,
         \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] ,
         \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] ,
         \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] ,
         \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] ,
         \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] ,
         \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] ,
         \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] ,
         \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] ,
         \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] ,
         \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] ,
         \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] ,
         \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] ,
         \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] ,
         \chs_in_f[0][DATA][7] , \chs_in_f[0][DATA][6] ,
         \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] ,
         \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] ,
         \chs_in_f[0][DATA][1] , \chs_in_f[0][DATA][0] ,
         \latches_out_b[4][ACK] , \latches_out_b[3][ACK] ,
         \latches_out_b[2][ACK] , \latches_out_b[1][ACK] ,
         \latches_out_b[0][ACK] ;
  output \chs_in_b[4][ACK] , \chs_in_b[3][ACK] , \chs_in_b[2][ACK] ,
         \chs_in_b[1][ACK] , \chs_in_b[0][ACK] , \latches_out_f[4][REQ] ,
         \latches_out_f[4][DATA][34] , \latches_out_f[4][DATA][33] ,
         \latches_out_f[4][DATA][32] , \latches_out_f[4][DATA][31] ,
         \latches_out_f[4][DATA][30] , \latches_out_f[4][DATA][29] ,
         \latches_out_f[4][DATA][28] , \latches_out_f[4][DATA][27] ,
         \latches_out_f[4][DATA][26] , \latches_out_f[4][DATA][25] ,
         \latches_out_f[4][DATA][24] , \latches_out_f[4][DATA][23] ,
         \latches_out_f[4][DATA][22] , \latches_out_f[4][DATA][21] ,
         \latches_out_f[4][DATA][20] , \latches_out_f[4][DATA][19] ,
         \latches_out_f[4][DATA][18] , \latches_out_f[4][DATA][17] ,
         \latches_out_f[4][DATA][16] , \latches_out_f[4][DATA][15] ,
         \latches_out_f[4][DATA][14] , \latches_out_f[4][DATA][13] ,
         \latches_out_f[4][DATA][12] , \latches_out_f[4][DATA][11] ,
         \latches_out_f[4][DATA][10] , \latches_out_f[4][DATA][9] ,
         \latches_out_f[4][DATA][8] , \latches_out_f[4][DATA][7] ,
         \latches_out_f[4][DATA][6] , \latches_out_f[4][DATA][5] ,
         \latches_out_f[4][DATA][4] , \latches_out_f[4][DATA][3] ,
         \latches_out_f[4][DATA][2] , \latches_out_f[4][DATA][1] ,
         \latches_out_f[4][DATA][0] , \latches_out_f[3][REQ] ,
         \latches_out_f[3][DATA][34] , \latches_out_f[3][DATA][33] ,
         \latches_out_f[3][DATA][32] , \latches_out_f[3][DATA][31] ,
         \latches_out_f[3][DATA][30] , \latches_out_f[3][DATA][29] ,
         \latches_out_f[3][DATA][28] , \latches_out_f[3][DATA][27] ,
         \latches_out_f[3][DATA][26] , \latches_out_f[3][DATA][25] ,
         \latches_out_f[3][DATA][24] , \latches_out_f[3][DATA][23] ,
         \latches_out_f[3][DATA][22] , \latches_out_f[3][DATA][21] ,
         \latches_out_f[3][DATA][20] , \latches_out_f[3][DATA][19] ,
         \latches_out_f[3][DATA][18] , \latches_out_f[3][DATA][17] ,
         \latches_out_f[3][DATA][16] , \latches_out_f[3][DATA][15] ,
         \latches_out_f[3][DATA][14] , \latches_out_f[3][DATA][13] ,
         \latches_out_f[3][DATA][12] , \latches_out_f[3][DATA][11] ,
         \latches_out_f[3][DATA][10] , \latches_out_f[3][DATA][9] ,
         \latches_out_f[3][DATA][8] , \latches_out_f[3][DATA][7] ,
         \latches_out_f[3][DATA][6] , \latches_out_f[3][DATA][5] ,
         \latches_out_f[3][DATA][4] , \latches_out_f[3][DATA][3] ,
         \latches_out_f[3][DATA][2] , \latches_out_f[3][DATA][1] ,
         \latches_out_f[3][DATA][0] , \latches_out_f[2][REQ] ,
         \latches_out_f[2][DATA][34] , \latches_out_f[2][DATA][33] ,
         \latches_out_f[2][DATA][32] , \latches_out_f[2][DATA][31] ,
         \latches_out_f[2][DATA][30] , \latches_out_f[2][DATA][29] ,
         \latches_out_f[2][DATA][28] , \latches_out_f[2][DATA][27] ,
         \latches_out_f[2][DATA][26] , \latches_out_f[2][DATA][25] ,
         \latches_out_f[2][DATA][24] , \latches_out_f[2][DATA][23] ,
         \latches_out_f[2][DATA][22] , \latches_out_f[2][DATA][21] ,
         \latches_out_f[2][DATA][20] , \latches_out_f[2][DATA][19] ,
         \latches_out_f[2][DATA][18] , \latches_out_f[2][DATA][17] ,
         \latches_out_f[2][DATA][16] , \latches_out_f[2][DATA][15] ,
         \latches_out_f[2][DATA][14] , \latches_out_f[2][DATA][13] ,
         \latches_out_f[2][DATA][12] , \latches_out_f[2][DATA][11] ,
         \latches_out_f[2][DATA][10] , \latches_out_f[2][DATA][9] ,
         \latches_out_f[2][DATA][8] , \latches_out_f[2][DATA][7] ,
         \latches_out_f[2][DATA][6] , \latches_out_f[2][DATA][5] ,
         \latches_out_f[2][DATA][4] , \latches_out_f[2][DATA][3] ,
         \latches_out_f[2][DATA][2] , \latches_out_f[2][DATA][1] ,
         \latches_out_f[2][DATA][0] , \latches_out_f[1][REQ] ,
         \latches_out_f[1][DATA][34] , \latches_out_f[1][DATA][33] ,
         \latches_out_f[1][DATA][32] , \latches_out_f[1][DATA][31] ,
         \latches_out_f[1][DATA][30] , \latches_out_f[1][DATA][29] ,
         \latches_out_f[1][DATA][28] , \latches_out_f[1][DATA][27] ,
         \latches_out_f[1][DATA][26] , \latches_out_f[1][DATA][25] ,
         \latches_out_f[1][DATA][24] , \latches_out_f[1][DATA][23] ,
         \latches_out_f[1][DATA][22] , \latches_out_f[1][DATA][21] ,
         \latches_out_f[1][DATA][20] , \latches_out_f[1][DATA][19] ,
         \latches_out_f[1][DATA][18] , \latches_out_f[1][DATA][17] ,
         \latches_out_f[1][DATA][16] , \latches_out_f[1][DATA][15] ,
         \latches_out_f[1][DATA][14] , \latches_out_f[1][DATA][13] ,
         \latches_out_f[1][DATA][12] , \latches_out_f[1][DATA][11] ,
         \latches_out_f[1][DATA][10] , \latches_out_f[1][DATA][9] ,
         \latches_out_f[1][DATA][8] , \latches_out_f[1][DATA][7] ,
         \latches_out_f[1][DATA][6] , \latches_out_f[1][DATA][5] ,
         \latches_out_f[1][DATA][4] , \latches_out_f[1][DATA][3] ,
         \latches_out_f[1][DATA][2] , \latches_out_f[1][DATA][1] ,
         \latches_out_f[1][DATA][0] , \latches_out_f[0][REQ] ,
         \latches_out_f[0][DATA][34] , \latches_out_f[0][DATA][33] ,
         \latches_out_f[0][DATA][32] , \latches_out_f[0][DATA][31] ,
         \latches_out_f[0][DATA][30] , \latches_out_f[0][DATA][29] ,
         \latches_out_f[0][DATA][28] , \latches_out_f[0][DATA][27] ,
         \latches_out_f[0][DATA][26] , \latches_out_f[0][DATA][25] ,
         \latches_out_f[0][DATA][24] , \latches_out_f[0][DATA][23] ,
         \latches_out_f[0][DATA][22] , \latches_out_f[0][DATA][21] ,
         \latches_out_f[0][DATA][20] , \latches_out_f[0][DATA][19] ,
         \latches_out_f[0][DATA][18] , \latches_out_f[0][DATA][17] ,
         \latches_out_f[0][DATA][16] , \latches_out_f[0][DATA][15] ,
         \latches_out_f[0][DATA][14] , \latches_out_f[0][DATA][13] ,
         \latches_out_f[0][DATA][12] , \latches_out_f[0][DATA][11] ,
         \latches_out_f[0][DATA][10] , \latches_out_f[0][DATA][9] ,
         \latches_out_f[0][DATA][8] , \latches_out_f[0][DATA][7] ,
         \latches_out_f[0][DATA][6] , \latches_out_f[0][DATA][5] ,
         \latches_out_f[0][DATA][4] , \latches_out_f[0][DATA][3] ,
         \latches_out_f[0][DATA][2] , \latches_out_f[0][DATA][1] ,
         \latches_out_f[0][DATA][0] ;
  wire   \latches_in_f[4][REQ] , \latches_in_f[4][DATA][34] ,
         \latches_in_f[4][DATA][33] , \latches_in_f[4][DATA][32] ,
         \latches_in_f[4][DATA][31] , \latches_in_f[4][DATA][30] ,
         \latches_in_f[4][DATA][29] , \latches_in_f[4][DATA][28] ,
         \latches_in_f[4][DATA][27] , \latches_in_f[4][DATA][26] ,
         \latches_in_f[4][DATA][25] , \latches_in_f[4][DATA][24] ,
         \latches_in_f[4][DATA][23] , \latches_in_f[4][DATA][22] ,
         \latches_in_f[4][DATA][21] , \latches_in_f[4][DATA][20] ,
         \latches_in_f[4][DATA][19] , \latches_in_f[4][DATA][18] ,
         \latches_in_f[4][DATA][17] , \latches_in_f[4][DATA][16] ,
         \latches_in_f[4][DATA][15] , \latches_in_f[4][DATA][14] ,
         \latches_in_f[4][DATA][13] , \latches_in_f[4][DATA][12] ,
         \latches_in_f[4][DATA][11] , \latches_in_f[4][DATA][10] ,
         \latches_in_f[4][DATA][9] , \latches_in_f[4][DATA][8] ,
         \latches_in_f[4][DATA][7] , \latches_in_f[4][DATA][6] ,
         \latches_in_f[4][DATA][5] , \latches_in_f[4][DATA][4] ,
         \latches_in_f[4][DATA][3] , \latches_in_f[4][DATA][2] ,
         \latches_in_f[4][DATA][1] , \latches_in_f[4][DATA][0] ,
         \latches_in_f[3][REQ] , \latches_in_f[3][DATA][34] ,
         \latches_in_f[3][DATA][33] , \latches_in_f[3][DATA][32] ,
         \latches_in_f[3][DATA][31] , \latches_in_f[3][DATA][30] ,
         \latches_in_f[3][DATA][29] , \latches_in_f[3][DATA][28] ,
         \latches_in_f[3][DATA][27] , \latches_in_f[3][DATA][26] ,
         \latches_in_f[3][DATA][25] , \latches_in_f[3][DATA][24] ,
         \latches_in_f[3][DATA][23] , \latches_in_f[3][DATA][22] ,
         \latches_in_f[3][DATA][21] , \latches_in_f[3][DATA][20] ,
         \latches_in_f[3][DATA][19] , \latches_in_f[3][DATA][18] ,
         \latches_in_f[3][DATA][17] , \latches_in_f[3][DATA][16] ,
         \latches_in_f[3][DATA][15] , \latches_in_f[3][DATA][14] ,
         \latches_in_f[3][DATA][13] , \latches_in_f[3][DATA][12] ,
         \latches_in_f[3][DATA][11] , \latches_in_f[3][DATA][10] ,
         \latches_in_f[3][DATA][9] , \latches_in_f[3][DATA][8] ,
         \latches_in_f[3][DATA][7] , \latches_in_f[3][DATA][6] ,
         \latches_in_f[3][DATA][5] , \latches_in_f[3][DATA][4] ,
         \latches_in_f[3][DATA][3] , \latches_in_f[3][DATA][2] ,
         \latches_in_f[3][DATA][1] , \latches_in_f[3][DATA][0] ,
         \latches_in_f[2][REQ] , \latches_in_f[2][DATA][34] ,
         \latches_in_f[2][DATA][33] , \latches_in_f[2][DATA][32] ,
         \latches_in_f[2][DATA][31] , \latches_in_f[2][DATA][30] ,
         \latches_in_f[2][DATA][29] , \latches_in_f[2][DATA][28] ,
         \latches_in_f[2][DATA][27] , \latches_in_f[2][DATA][26] ,
         \latches_in_f[2][DATA][25] , \latches_in_f[2][DATA][24] ,
         \latches_in_f[2][DATA][23] , \latches_in_f[2][DATA][22] ,
         \latches_in_f[2][DATA][21] , \latches_in_f[2][DATA][20] ,
         \latches_in_f[2][DATA][19] , \latches_in_f[2][DATA][18] ,
         \latches_in_f[2][DATA][17] , \latches_in_f[2][DATA][16] ,
         \latches_in_f[2][DATA][15] , \latches_in_f[2][DATA][14] ,
         \latches_in_f[2][DATA][13] , \latches_in_f[2][DATA][12] ,
         \latches_in_f[2][DATA][11] , \latches_in_f[2][DATA][10] ,
         \latches_in_f[2][DATA][9] , \latches_in_f[2][DATA][8] ,
         \latches_in_f[2][DATA][7] , \latches_in_f[2][DATA][6] ,
         \latches_in_f[2][DATA][5] , \latches_in_f[2][DATA][4] ,
         \latches_in_f[2][DATA][3] , \latches_in_f[2][DATA][2] ,
         \latches_in_f[2][DATA][1] , \latches_in_f[2][DATA][0] ,
         \latches_in_f[1][REQ] , \latches_in_f[1][DATA][34] ,
         \latches_in_f[1][DATA][33] , \latches_in_f[1][DATA][32] ,
         \latches_in_f[1][DATA][31] , \latches_in_f[1][DATA][30] ,
         \latches_in_f[1][DATA][29] , \latches_in_f[1][DATA][28] ,
         \latches_in_f[1][DATA][27] , \latches_in_f[1][DATA][26] ,
         \latches_in_f[1][DATA][25] , \latches_in_f[1][DATA][24] ,
         \latches_in_f[1][DATA][23] , \latches_in_f[1][DATA][22] ,
         \latches_in_f[1][DATA][21] , \latches_in_f[1][DATA][20] ,
         \latches_in_f[1][DATA][19] , \latches_in_f[1][DATA][18] ,
         \latches_in_f[1][DATA][17] , \latches_in_f[1][DATA][16] ,
         \latches_in_f[1][DATA][15] , \latches_in_f[1][DATA][14] ,
         \latches_in_f[1][DATA][13] , \latches_in_f[1][DATA][12] ,
         \latches_in_f[1][DATA][11] , \latches_in_f[1][DATA][10] ,
         \latches_in_f[1][DATA][9] , \latches_in_f[1][DATA][8] ,
         \latches_in_f[1][DATA][7] , \latches_in_f[1][DATA][6] ,
         \latches_in_f[1][DATA][5] , \latches_in_f[1][DATA][4] ,
         \latches_in_f[1][DATA][3] , \latches_in_f[1][DATA][2] ,
         \latches_in_f[1][DATA][1] , \latches_in_f[1][DATA][0] ,
         \latches_in_f[0][REQ] , \latches_in_f[0][DATA][34] ,
         \latches_in_f[0][DATA][33] , \latches_in_f[0][DATA][32] ,
         \latches_in_f[0][DATA][31] , \latches_in_f[0][DATA][30] ,
         \latches_in_f[0][DATA][29] , \latches_in_f[0][DATA][28] ,
         \latches_in_f[0][DATA][27] , \latches_in_f[0][DATA][26] ,
         \latches_in_f[0][DATA][25] , \latches_in_f[0][DATA][24] ,
         \latches_in_f[0][DATA][23] , \latches_in_f[0][DATA][22] ,
         \latches_in_f[0][DATA][21] , \latches_in_f[0][DATA][20] ,
         \latches_in_f[0][DATA][19] , \latches_in_f[0][DATA][18] ,
         \latches_in_f[0][DATA][17] , \latches_in_f[0][DATA][16] ,
         \latches_in_f[0][DATA][15] , \latches_in_f[0][DATA][14] ,
         \latches_in_f[0][DATA][13] , \latches_in_f[0][DATA][12] ,
         \latches_in_f[0][DATA][11] , \latches_in_f[0][DATA][10] ,
         \latches_in_f[0][DATA][9] , \latches_in_f[0][DATA][8] ,
         \latches_in_f[0][DATA][7] , \latches_in_f[0][DATA][6] ,
         \latches_in_f[0][DATA][5] , \latches_in_f[0][DATA][4] ,
         \latches_in_f[0][DATA][3] , \latches_in_f[0][DATA][2] ,
         \latches_in_f[0][DATA][1] , \latches_in_f[0][DATA][0] ,
         \latches_in_b[4][ACK] , \latches_in_b[3][ACK] ,
         \latches_in_b[2][ACK] , \latches_in_b[1][ACK] ,
         \latches_in_b[0][ACK] , n1;

  crossbar_3 crossbar ( .preset(n1), .switch_sel({\switch_sel[4][4] , 
        \switch_sel[4][3] , \switch_sel[4][2] , \switch_sel[4][1] , 
        \switch_sel[4][0] , \switch_sel[3][4] , \switch_sel[3][3] , 
        \switch_sel[3][2] , \switch_sel[3][1] , \switch_sel[3][0] , 
        \switch_sel[2][4] , \switch_sel[2][3] , \switch_sel[2][2] , 
        \switch_sel[2][1] , \switch_sel[2][0] , \switch_sel[1][4] , 
        \switch_sel[1][3] , \switch_sel[1][2] , \switch_sel[1][1] , 
        \switch_sel[1][0] , \switch_sel[0][4] , \switch_sel[0][3] , 
        \switch_sel[0][2] , \switch_sel[0][1] , \switch_sel[0][0] }), 
        .chs_in_f({\chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] , 
        \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] , 
        \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] , 
        \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] , 
        \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] , 
        \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] , 
        \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] , 
        \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] , 
        \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] , 
        \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] , 
        \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] , 
        \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] , 
        \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] , 
        \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] , \chs_in_f[4][DATA][7] , 
        \chs_in_f[4][DATA][6] , \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] , 
        \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] , \chs_in_f[4][DATA][1] , 
        \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] , \chs_in_f[3][DATA][34] , 
        \chs_in_f[3][DATA][33] , \chs_in_f[3][DATA][32] , 
        \chs_in_f[3][DATA][31] , \chs_in_f[3][DATA][30] , 
        \chs_in_f[3][DATA][29] , \chs_in_f[3][DATA][28] , 
        \chs_in_f[3][DATA][27] , \chs_in_f[3][DATA][26] , 
        \chs_in_f[3][DATA][25] , \chs_in_f[3][DATA][24] , 
        \chs_in_f[3][DATA][23] , \chs_in_f[3][DATA][22] , 
        \chs_in_f[3][DATA][21] , \chs_in_f[3][DATA][20] , 
        \chs_in_f[3][DATA][19] , \chs_in_f[3][DATA][18] , 
        \chs_in_f[3][DATA][17] , \chs_in_f[3][DATA][16] , 
        \chs_in_f[3][DATA][15] , \chs_in_f[3][DATA][14] , 
        \chs_in_f[3][DATA][13] , \chs_in_f[3][DATA][12] , 
        \chs_in_f[3][DATA][11] , \chs_in_f[3][DATA][10] , 
        \chs_in_f[3][DATA][9] , \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] , 
        \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] , \chs_in_f[3][DATA][4] , 
        \chs_in_f[3][DATA][3] , \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] , 
        \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] , 
        \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] , 
        \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] , 
        \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] , 
        \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] , 
        \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] , 
        \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] , 
        \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] , 
        \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] , 
        \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] , 
        \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] , 
        \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] , 
        \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] , 
        \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] , \chs_in_f[2][DATA][7] , 
        \chs_in_f[2][DATA][6] , \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] , 
        \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] , \chs_in_f[2][DATA][1] , 
        \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] , \chs_in_f[1][DATA][34] , 
        \chs_in_f[1][DATA][33] , \chs_in_f[1][DATA][32] , 
        \chs_in_f[1][DATA][31] , \chs_in_f[1][DATA][30] , 
        \chs_in_f[1][DATA][29] , \chs_in_f[1][DATA][28] , 
        \chs_in_f[1][DATA][27] , \chs_in_f[1][DATA][26] , 
        \chs_in_f[1][DATA][25] , \chs_in_f[1][DATA][24] , 
        \chs_in_f[1][DATA][23] , \chs_in_f[1][DATA][22] , 
        \chs_in_f[1][DATA][21] , \chs_in_f[1][DATA][20] , 
        \chs_in_f[1][DATA][19] , \chs_in_f[1][DATA][18] , 
        \chs_in_f[1][DATA][17] , \chs_in_f[1][DATA][16] , 
        \chs_in_f[1][DATA][15] , \chs_in_f[1][DATA][14] , 
        \chs_in_f[1][DATA][13] , \chs_in_f[1][DATA][12] , 
        \chs_in_f[1][DATA][11] , \chs_in_f[1][DATA][10] , 
        \chs_in_f[1][DATA][9] , \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] , 
        \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] , \chs_in_f[1][DATA][4] , 
        \chs_in_f[1][DATA][3] , \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] , 
        \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] , 
        \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] , 
        \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] , 
        \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] , 
        \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] , 
        \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] , 
        \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] , 
        \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] , 
        \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] , 
        \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] , 
        \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] , 
        \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] , 
        \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] , 
        \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] , \chs_in_f[0][DATA][7] , 
        \chs_in_f[0][DATA][6] , \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] , 
        \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] , \chs_in_f[0][DATA][1] , 
        \chs_in_f[0][DATA][0] }), .chs_in_b({\chs_in_b[4][ACK] , 
        \chs_in_b[3][ACK] , \chs_in_b[2][ACK] , \chs_in_b[1][ACK] , 
        \chs_in_b[0][ACK] }), .chs_out_f({\latches_in_f[4][REQ] , 
        \latches_in_f[4][DATA][34] , \latches_in_f[4][DATA][33] , 
        \latches_in_f[4][DATA][32] , \latches_in_f[4][DATA][31] , 
        \latches_in_f[4][DATA][30] , \latches_in_f[4][DATA][29] , 
        \latches_in_f[4][DATA][28] , \latches_in_f[4][DATA][27] , 
        \latches_in_f[4][DATA][26] , \latches_in_f[4][DATA][25] , 
        \latches_in_f[4][DATA][24] , \latches_in_f[4][DATA][23] , 
        \latches_in_f[4][DATA][22] , \latches_in_f[4][DATA][21] , 
        \latches_in_f[4][DATA][20] , \latches_in_f[4][DATA][19] , 
        \latches_in_f[4][DATA][18] , \latches_in_f[4][DATA][17] , 
        \latches_in_f[4][DATA][16] , \latches_in_f[4][DATA][15] , 
        \latches_in_f[4][DATA][14] , \latches_in_f[4][DATA][13] , 
        \latches_in_f[4][DATA][12] , \latches_in_f[4][DATA][11] , 
        \latches_in_f[4][DATA][10] , \latches_in_f[4][DATA][9] , 
        \latches_in_f[4][DATA][8] , \latches_in_f[4][DATA][7] , 
        \latches_in_f[4][DATA][6] , \latches_in_f[4][DATA][5] , 
        \latches_in_f[4][DATA][4] , \latches_in_f[4][DATA][3] , 
        \latches_in_f[4][DATA][2] , \latches_in_f[4][DATA][1] , 
        \latches_in_f[4][DATA][0] , \latches_in_f[3][REQ] , 
        \latches_in_f[3][DATA][34] , \latches_in_f[3][DATA][33] , 
        \latches_in_f[3][DATA][32] , \latches_in_f[3][DATA][31] , 
        \latches_in_f[3][DATA][30] , \latches_in_f[3][DATA][29] , 
        \latches_in_f[3][DATA][28] , \latches_in_f[3][DATA][27] , 
        \latches_in_f[3][DATA][26] , \latches_in_f[3][DATA][25] , 
        \latches_in_f[3][DATA][24] , \latches_in_f[3][DATA][23] , 
        \latches_in_f[3][DATA][22] , \latches_in_f[3][DATA][21] , 
        \latches_in_f[3][DATA][20] , \latches_in_f[3][DATA][19] , 
        \latches_in_f[3][DATA][18] , \latches_in_f[3][DATA][17] , 
        \latches_in_f[3][DATA][16] , \latches_in_f[3][DATA][15] , 
        \latches_in_f[3][DATA][14] , \latches_in_f[3][DATA][13] , 
        \latches_in_f[3][DATA][12] , \latches_in_f[3][DATA][11] , 
        \latches_in_f[3][DATA][10] , \latches_in_f[3][DATA][9] , 
        \latches_in_f[3][DATA][8] , \latches_in_f[3][DATA][7] , 
        \latches_in_f[3][DATA][6] , \latches_in_f[3][DATA][5] , 
        \latches_in_f[3][DATA][4] , \latches_in_f[3][DATA][3] , 
        \latches_in_f[3][DATA][2] , \latches_in_f[3][DATA][1] , 
        \latches_in_f[3][DATA][0] , \latches_in_f[2][REQ] , 
        \latches_in_f[2][DATA][34] , \latches_in_f[2][DATA][33] , 
        \latches_in_f[2][DATA][32] , \latches_in_f[2][DATA][31] , 
        \latches_in_f[2][DATA][30] , \latches_in_f[2][DATA][29] , 
        \latches_in_f[2][DATA][28] , \latches_in_f[2][DATA][27] , 
        \latches_in_f[2][DATA][26] , \latches_in_f[2][DATA][25] , 
        \latches_in_f[2][DATA][24] , \latches_in_f[2][DATA][23] , 
        \latches_in_f[2][DATA][22] , \latches_in_f[2][DATA][21] , 
        \latches_in_f[2][DATA][20] , \latches_in_f[2][DATA][19] , 
        \latches_in_f[2][DATA][18] , \latches_in_f[2][DATA][17] , 
        \latches_in_f[2][DATA][16] , \latches_in_f[2][DATA][15] , 
        \latches_in_f[2][DATA][14] , \latches_in_f[2][DATA][13] , 
        \latches_in_f[2][DATA][12] , \latches_in_f[2][DATA][11] , 
        \latches_in_f[2][DATA][10] , \latches_in_f[2][DATA][9] , 
        \latches_in_f[2][DATA][8] , \latches_in_f[2][DATA][7] , 
        \latches_in_f[2][DATA][6] , \latches_in_f[2][DATA][5] , 
        \latches_in_f[2][DATA][4] , \latches_in_f[2][DATA][3] , 
        \latches_in_f[2][DATA][2] , \latches_in_f[2][DATA][1] , 
        \latches_in_f[2][DATA][0] , \latches_in_f[1][REQ] , 
        \latches_in_f[1][DATA][34] , \latches_in_f[1][DATA][33] , 
        \latches_in_f[1][DATA][32] , \latches_in_f[1][DATA][31] , 
        \latches_in_f[1][DATA][30] , \latches_in_f[1][DATA][29] , 
        \latches_in_f[1][DATA][28] , \latches_in_f[1][DATA][27] , 
        \latches_in_f[1][DATA][26] , \latches_in_f[1][DATA][25] , 
        \latches_in_f[1][DATA][24] , \latches_in_f[1][DATA][23] , 
        \latches_in_f[1][DATA][22] , \latches_in_f[1][DATA][21] , 
        \latches_in_f[1][DATA][20] , \latches_in_f[1][DATA][19] , 
        \latches_in_f[1][DATA][18] , \latches_in_f[1][DATA][17] , 
        \latches_in_f[1][DATA][16] , \latches_in_f[1][DATA][15] , 
        \latches_in_f[1][DATA][14] , \latches_in_f[1][DATA][13] , 
        \latches_in_f[1][DATA][12] , \latches_in_f[1][DATA][11] , 
        \latches_in_f[1][DATA][10] , \latches_in_f[1][DATA][9] , 
        \latches_in_f[1][DATA][8] , \latches_in_f[1][DATA][7] , 
        \latches_in_f[1][DATA][6] , \latches_in_f[1][DATA][5] , 
        \latches_in_f[1][DATA][4] , \latches_in_f[1][DATA][3] , 
        \latches_in_f[1][DATA][2] , \latches_in_f[1][DATA][1] , 
        \latches_in_f[1][DATA][0] , \latches_in_f[0][REQ] , 
        \latches_in_f[0][DATA][34] , \latches_in_f[0][DATA][33] , 
        \latches_in_f[0][DATA][32] , \latches_in_f[0][DATA][31] , 
        \latches_in_f[0][DATA][30] , \latches_in_f[0][DATA][29] , 
        \latches_in_f[0][DATA][28] , \latches_in_f[0][DATA][27] , 
        \latches_in_f[0][DATA][26] , \latches_in_f[0][DATA][25] , 
        \latches_in_f[0][DATA][24] , \latches_in_f[0][DATA][23] , 
        \latches_in_f[0][DATA][22] , \latches_in_f[0][DATA][21] , 
        \latches_in_f[0][DATA][20] , \latches_in_f[0][DATA][19] , 
        \latches_in_f[0][DATA][18] , \latches_in_f[0][DATA][17] , 
        \latches_in_f[0][DATA][16] , \latches_in_f[0][DATA][15] , 
        \latches_in_f[0][DATA][14] , \latches_in_f[0][DATA][13] , 
        \latches_in_f[0][DATA][12] , \latches_in_f[0][DATA][11] , 
        \latches_in_f[0][DATA][10] , \latches_in_f[0][DATA][9] , 
        \latches_in_f[0][DATA][8] , \latches_in_f[0][DATA][7] , 
        \latches_in_f[0][DATA][6] , \latches_in_f[0][DATA][5] , 
        \latches_in_f[0][DATA][4] , \latches_in_f[0][DATA][3] , 
        \latches_in_f[0][DATA][2] , \latches_in_f[0][DATA][1] , 
        \latches_in_f[0][DATA][0] }), .chs_out_b({\latches_in_b[4][ACK] , 
        \latches_in_b[3][ACK] , \latches_in_b[2][ACK] , \latches_in_b[1][ACK] , 
        \latches_in_b[0][ACK] }) );
  channel_latch_0_000000000_15 ch_latch_4 ( .preset(n1), .left_in({
        \latches_in_f[4][REQ] , \latches_in_f[4][DATA][34] , 
        \latches_in_f[4][DATA][33] , \latches_in_f[4][DATA][32] , 
        \latches_in_f[4][DATA][31] , \latches_in_f[4][DATA][30] , 
        \latches_in_f[4][DATA][29] , \latches_in_f[4][DATA][28] , 
        \latches_in_f[4][DATA][27] , \latches_in_f[4][DATA][26] , 
        \latches_in_f[4][DATA][25] , \latches_in_f[4][DATA][24] , 
        \latches_in_f[4][DATA][23] , \latches_in_f[4][DATA][22] , 
        \latches_in_f[4][DATA][21] , \latches_in_f[4][DATA][20] , 
        \latches_in_f[4][DATA][19] , \latches_in_f[4][DATA][18] , 
        \latches_in_f[4][DATA][17] , \latches_in_f[4][DATA][16] , 
        \latches_in_f[4][DATA][15] , \latches_in_f[4][DATA][14] , 
        \latches_in_f[4][DATA][13] , \latches_in_f[4][DATA][12] , 
        \latches_in_f[4][DATA][11] , \latches_in_f[4][DATA][10] , 
        \latches_in_f[4][DATA][9] , \latches_in_f[4][DATA][8] , 
        \latches_in_f[4][DATA][7] , \latches_in_f[4][DATA][6] , 
        \latches_in_f[4][DATA][5] , \latches_in_f[4][DATA][4] , 
        \latches_in_f[4][DATA][3] , \latches_in_f[4][DATA][2] , 
        \latches_in_f[4][DATA][1] , \latches_in_f[4][DATA][0] }), .left_out(
        \latches_in_b[4][ACK] ), .right_out({\latches_out_f[4][REQ] , 
        \latches_out_f[4][DATA][34] , \latches_out_f[4][DATA][33] , 
        \latches_out_f[4][DATA][32] , \latches_out_f[4][DATA][31] , 
        \latches_out_f[4][DATA][30] , \latches_out_f[4][DATA][29] , 
        \latches_out_f[4][DATA][28] , \latches_out_f[4][DATA][27] , 
        \latches_out_f[4][DATA][26] , \latches_out_f[4][DATA][25] , 
        \latches_out_f[4][DATA][24] , \latches_out_f[4][DATA][23] , 
        \latches_out_f[4][DATA][22] , \latches_out_f[4][DATA][21] , 
        \latches_out_f[4][DATA][20] , \latches_out_f[4][DATA][19] , 
        \latches_out_f[4][DATA][18] , \latches_out_f[4][DATA][17] , 
        \latches_out_f[4][DATA][16] , \latches_out_f[4][DATA][15] , 
        \latches_out_f[4][DATA][14] , \latches_out_f[4][DATA][13] , 
        \latches_out_f[4][DATA][12] , \latches_out_f[4][DATA][11] , 
        \latches_out_f[4][DATA][10] , \latches_out_f[4][DATA][9] , 
        \latches_out_f[4][DATA][8] , \latches_out_f[4][DATA][7] , 
        \latches_out_f[4][DATA][6] , \latches_out_f[4][DATA][5] , 
        \latches_out_f[4][DATA][4] , \latches_out_f[4][DATA][3] , 
        \latches_out_f[4][DATA][2] , \latches_out_f[4][DATA][1] , 
        \latches_out_f[4][DATA][0] }), .right_in(\latches_out_b[4][ACK] ) );
  channel_latch_0_000000000_14 ch_latch_3 ( .preset(n1), .left_in({
        \latches_in_f[3][REQ] , \latches_in_f[3][DATA][34] , 
        \latches_in_f[3][DATA][33] , \latches_in_f[3][DATA][32] , 
        \latches_in_f[3][DATA][31] , \latches_in_f[3][DATA][30] , 
        \latches_in_f[3][DATA][29] , \latches_in_f[3][DATA][28] , 
        \latches_in_f[3][DATA][27] , \latches_in_f[3][DATA][26] , 
        \latches_in_f[3][DATA][25] , \latches_in_f[3][DATA][24] , 
        \latches_in_f[3][DATA][23] , \latches_in_f[3][DATA][22] , 
        \latches_in_f[3][DATA][21] , \latches_in_f[3][DATA][20] , 
        \latches_in_f[3][DATA][19] , \latches_in_f[3][DATA][18] , 
        \latches_in_f[3][DATA][17] , \latches_in_f[3][DATA][16] , 
        \latches_in_f[3][DATA][15] , \latches_in_f[3][DATA][14] , 
        \latches_in_f[3][DATA][13] , \latches_in_f[3][DATA][12] , 
        \latches_in_f[3][DATA][11] , \latches_in_f[3][DATA][10] , 
        \latches_in_f[3][DATA][9] , \latches_in_f[3][DATA][8] , 
        \latches_in_f[3][DATA][7] , \latches_in_f[3][DATA][6] , 
        \latches_in_f[3][DATA][5] , \latches_in_f[3][DATA][4] , 
        \latches_in_f[3][DATA][3] , \latches_in_f[3][DATA][2] , 
        \latches_in_f[3][DATA][1] , \latches_in_f[3][DATA][0] }), .left_out(
        \latches_in_b[3][ACK] ), .right_out({\latches_out_f[3][REQ] , 
        \latches_out_f[3][DATA][34] , \latches_out_f[3][DATA][33] , 
        \latches_out_f[3][DATA][32] , \latches_out_f[3][DATA][31] , 
        \latches_out_f[3][DATA][30] , \latches_out_f[3][DATA][29] , 
        \latches_out_f[3][DATA][28] , \latches_out_f[3][DATA][27] , 
        \latches_out_f[3][DATA][26] , \latches_out_f[3][DATA][25] , 
        \latches_out_f[3][DATA][24] , \latches_out_f[3][DATA][23] , 
        \latches_out_f[3][DATA][22] , \latches_out_f[3][DATA][21] , 
        \latches_out_f[3][DATA][20] , \latches_out_f[3][DATA][19] , 
        \latches_out_f[3][DATA][18] , \latches_out_f[3][DATA][17] , 
        \latches_out_f[3][DATA][16] , \latches_out_f[3][DATA][15] , 
        \latches_out_f[3][DATA][14] , \latches_out_f[3][DATA][13] , 
        \latches_out_f[3][DATA][12] , \latches_out_f[3][DATA][11] , 
        \latches_out_f[3][DATA][10] , \latches_out_f[3][DATA][9] , 
        \latches_out_f[3][DATA][8] , \latches_out_f[3][DATA][7] , 
        \latches_out_f[3][DATA][6] , \latches_out_f[3][DATA][5] , 
        \latches_out_f[3][DATA][4] , \latches_out_f[3][DATA][3] , 
        \latches_out_f[3][DATA][2] , \latches_out_f[3][DATA][1] , 
        \latches_out_f[3][DATA][0] }), .right_in(\latches_out_b[3][ACK] ) );
  channel_latch_0_000000000_13 ch_latch_2 ( .preset(n1), .left_in({
        \latches_in_f[2][REQ] , \latches_in_f[2][DATA][34] , 
        \latches_in_f[2][DATA][33] , \latches_in_f[2][DATA][32] , 
        \latches_in_f[2][DATA][31] , \latches_in_f[2][DATA][30] , 
        \latches_in_f[2][DATA][29] , \latches_in_f[2][DATA][28] , 
        \latches_in_f[2][DATA][27] , \latches_in_f[2][DATA][26] , 
        \latches_in_f[2][DATA][25] , \latches_in_f[2][DATA][24] , 
        \latches_in_f[2][DATA][23] , \latches_in_f[2][DATA][22] , 
        \latches_in_f[2][DATA][21] , \latches_in_f[2][DATA][20] , 
        \latches_in_f[2][DATA][19] , \latches_in_f[2][DATA][18] , 
        \latches_in_f[2][DATA][17] , \latches_in_f[2][DATA][16] , 
        \latches_in_f[2][DATA][15] , \latches_in_f[2][DATA][14] , 
        \latches_in_f[2][DATA][13] , \latches_in_f[2][DATA][12] , 
        \latches_in_f[2][DATA][11] , \latches_in_f[2][DATA][10] , 
        \latches_in_f[2][DATA][9] , \latches_in_f[2][DATA][8] , 
        \latches_in_f[2][DATA][7] , \latches_in_f[2][DATA][6] , 
        \latches_in_f[2][DATA][5] , \latches_in_f[2][DATA][4] , 
        \latches_in_f[2][DATA][3] , \latches_in_f[2][DATA][2] , 
        \latches_in_f[2][DATA][1] , \latches_in_f[2][DATA][0] }), .left_out(
        \latches_in_b[2][ACK] ), .right_out({\latches_out_f[2][REQ] , 
        \latches_out_f[2][DATA][34] , \latches_out_f[2][DATA][33] , 
        \latches_out_f[2][DATA][32] , \latches_out_f[2][DATA][31] , 
        \latches_out_f[2][DATA][30] , \latches_out_f[2][DATA][29] , 
        \latches_out_f[2][DATA][28] , \latches_out_f[2][DATA][27] , 
        \latches_out_f[2][DATA][26] , \latches_out_f[2][DATA][25] , 
        \latches_out_f[2][DATA][24] , \latches_out_f[2][DATA][23] , 
        \latches_out_f[2][DATA][22] , \latches_out_f[2][DATA][21] , 
        \latches_out_f[2][DATA][20] , \latches_out_f[2][DATA][19] , 
        \latches_out_f[2][DATA][18] , \latches_out_f[2][DATA][17] , 
        \latches_out_f[2][DATA][16] , \latches_out_f[2][DATA][15] , 
        \latches_out_f[2][DATA][14] , \latches_out_f[2][DATA][13] , 
        \latches_out_f[2][DATA][12] , \latches_out_f[2][DATA][11] , 
        \latches_out_f[2][DATA][10] , \latches_out_f[2][DATA][9] , 
        \latches_out_f[2][DATA][8] , \latches_out_f[2][DATA][7] , 
        \latches_out_f[2][DATA][6] , \latches_out_f[2][DATA][5] , 
        \latches_out_f[2][DATA][4] , \latches_out_f[2][DATA][3] , 
        \latches_out_f[2][DATA][2] , \latches_out_f[2][DATA][1] , 
        \latches_out_f[2][DATA][0] }), .right_in(\latches_out_b[2][ACK] ) );
  channel_latch_0_000000000_12 ch_latch_1 ( .preset(n1), .left_in({
        \latches_in_f[1][REQ] , \latches_in_f[1][DATA][34] , 
        \latches_in_f[1][DATA][33] , \latches_in_f[1][DATA][32] , 
        \latches_in_f[1][DATA][31] , \latches_in_f[1][DATA][30] , 
        \latches_in_f[1][DATA][29] , \latches_in_f[1][DATA][28] , 
        \latches_in_f[1][DATA][27] , \latches_in_f[1][DATA][26] , 
        \latches_in_f[1][DATA][25] , \latches_in_f[1][DATA][24] , 
        \latches_in_f[1][DATA][23] , \latches_in_f[1][DATA][22] , 
        \latches_in_f[1][DATA][21] , \latches_in_f[1][DATA][20] , 
        \latches_in_f[1][DATA][19] , \latches_in_f[1][DATA][18] , 
        \latches_in_f[1][DATA][17] , \latches_in_f[1][DATA][16] , 
        \latches_in_f[1][DATA][15] , \latches_in_f[1][DATA][14] , 
        \latches_in_f[1][DATA][13] , \latches_in_f[1][DATA][12] , 
        \latches_in_f[1][DATA][11] , \latches_in_f[1][DATA][10] , 
        \latches_in_f[1][DATA][9] , \latches_in_f[1][DATA][8] , 
        \latches_in_f[1][DATA][7] , \latches_in_f[1][DATA][6] , 
        \latches_in_f[1][DATA][5] , \latches_in_f[1][DATA][4] , 
        \latches_in_f[1][DATA][3] , \latches_in_f[1][DATA][2] , 
        \latches_in_f[1][DATA][1] , \latches_in_f[1][DATA][0] }), .left_out(
        \latches_in_b[1][ACK] ), .right_out({\latches_out_f[1][REQ] , 
        \latches_out_f[1][DATA][34] , \latches_out_f[1][DATA][33] , 
        \latches_out_f[1][DATA][32] , \latches_out_f[1][DATA][31] , 
        \latches_out_f[1][DATA][30] , \latches_out_f[1][DATA][29] , 
        \latches_out_f[1][DATA][28] , \latches_out_f[1][DATA][27] , 
        \latches_out_f[1][DATA][26] , \latches_out_f[1][DATA][25] , 
        \latches_out_f[1][DATA][24] , \latches_out_f[1][DATA][23] , 
        \latches_out_f[1][DATA][22] , \latches_out_f[1][DATA][21] , 
        \latches_out_f[1][DATA][20] , \latches_out_f[1][DATA][19] , 
        \latches_out_f[1][DATA][18] , \latches_out_f[1][DATA][17] , 
        \latches_out_f[1][DATA][16] , \latches_out_f[1][DATA][15] , 
        \latches_out_f[1][DATA][14] , \latches_out_f[1][DATA][13] , 
        \latches_out_f[1][DATA][12] , \latches_out_f[1][DATA][11] , 
        \latches_out_f[1][DATA][10] , \latches_out_f[1][DATA][9] , 
        \latches_out_f[1][DATA][8] , \latches_out_f[1][DATA][7] , 
        \latches_out_f[1][DATA][6] , \latches_out_f[1][DATA][5] , 
        \latches_out_f[1][DATA][4] , \latches_out_f[1][DATA][3] , 
        \latches_out_f[1][DATA][2] , \latches_out_f[1][DATA][1] , 
        \latches_out_f[1][DATA][0] }), .right_in(\latches_out_b[1][ACK] ) );
  channel_latch_0_000000000_11 ch_latch_0 ( .preset(n1), .left_in({
        \latches_in_f[0][REQ] , \latches_in_f[0][DATA][34] , 
        \latches_in_f[0][DATA][33] , \latches_in_f[0][DATA][32] , 
        \latches_in_f[0][DATA][31] , \latches_in_f[0][DATA][30] , 
        \latches_in_f[0][DATA][29] , \latches_in_f[0][DATA][28] , 
        \latches_in_f[0][DATA][27] , \latches_in_f[0][DATA][26] , 
        \latches_in_f[0][DATA][25] , \latches_in_f[0][DATA][24] , 
        \latches_in_f[0][DATA][23] , \latches_in_f[0][DATA][22] , 
        \latches_in_f[0][DATA][21] , \latches_in_f[0][DATA][20] , 
        \latches_in_f[0][DATA][19] , \latches_in_f[0][DATA][18] , 
        \latches_in_f[0][DATA][17] , \latches_in_f[0][DATA][16] , 
        \latches_in_f[0][DATA][15] , \latches_in_f[0][DATA][14] , 
        \latches_in_f[0][DATA][13] , \latches_in_f[0][DATA][12] , 
        \latches_in_f[0][DATA][11] , \latches_in_f[0][DATA][10] , 
        \latches_in_f[0][DATA][9] , \latches_in_f[0][DATA][8] , 
        \latches_in_f[0][DATA][7] , \latches_in_f[0][DATA][6] , 
        \latches_in_f[0][DATA][5] , \latches_in_f[0][DATA][4] , 
        \latches_in_f[0][DATA][3] , \latches_in_f[0][DATA][2] , 
        \latches_in_f[0][DATA][1] , \latches_in_f[0][DATA][0] }), .left_out(
        \latches_in_b[0][ACK] ), .right_out({\latches_out_f[0][REQ] , 
        \latches_out_f[0][DATA][34] , \latches_out_f[0][DATA][33] , 
        \latches_out_f[0][DATA][32] , \latches_out_f[0][DATA][31] , 
        \latches_out_f[0][DATA][30] , \latches_out_f[0][DATA][29] , 
        \latches_out_f[0][DATA][28] , \latches_out_f[0][DATA][27] , 
        \latches_out_f[0][DATA][26] , \latches_out_f[0][DATA][25] , 
        \latches_out_f[0][DATA][24] , \latches_out_f[0][DATA][23] , 
        \latches_out_f[0][DATA][22] , \latches_out_f[0][DATA][21] , 
        \latches_out_f[0][DATA][20] , \latches_out_f[0][DATA][19] , 
        \latches_out_f[0][DATA][18] , \latches_out_f[0][DATA][17] , 
        \latches_out_f[0][DATA][16] , \latches_out_f[0][DATA][15] , 
        \latches_out_f[0][DATA][14] , \latches_out_f[0][DATA][13] , 
        \latches_out_f[0][DATA][12] , \latches_out_f[0][DATA][11] , 
        \latches_out_f[0][DATA][10] , \latches_out_f[0][DATA][9] , 
        \latches_out_f[0][DATA][8] , \latches_out_f[0][DATA][7] , 
        \latches_out_f[0][DATA][6] , \latches_out_f[0][DATA][5] , 
        \latches_out_f[0][DATA][4] , \latches_out_f[0][DATA][3] , 
        \latches_out_f[0][DATA][2] , \latches_out_f[0][DATA][1] , 
        \latches_out_f[0][DATA][0] }), .right_in(\latches_out_b[0][ACK] ) );
  HS65_LS_BFX9 U1 ( .A(preset), .Z(n1) );
endmodule


module noc_switch_3 ( preset, .north_in_f({\north_in_f[REQ] , 
        \north_in_f[DATA][34] , \north_in_f[DATA][33] , \north_in_f[DATA][32] , 
        \north_in_f[DATA][31] , \north_in_f[DATA][30] , \north_in_f[DATA][29] , 
        \north_in_f[DATA][28] , \north_in_f[DATA][27] , \north_in_f[DATA][26] , 
        \north_in_f[DATA][25] , \north_in_f[DATA][24] , \north_in_f[DATA][23] , 
        \north_in_f[DATA][22] , \north_in_f[DATA][21] , \north_in_f[DATA][20] , 
        \north_in_f[DATA][19] , \north_in_f[DATA][18] , \north_in_f[DATA][17] , 
        \north_in_f[DATA][16] , \north_in_f[DATA][15] , \north_in_f[DATA][14] , 
        \north_in_f[DATA][13] , \north_in_f[DATA][12] , \north_in_f[DATA][11] , 
        \north_in_f[DATA][10] , \north_in_f[DATA][9] , \north_in_f[DATA][8] , 
        \north_in_f[DATA][7] , \north_in_f[DATA][6] , \north_in_f[DATA][5] , 
        \north_in_f[DATA][4] , \north_in_f[DATA][3] , \north_in_f[DATA][2] , 
        \north_in_f[DATA][1] , \north_in_f[DATA][0] }), .north_in_b(
        \north_in_b[ACK] ), .east_in_f({\east_in_f[REQ] , 
        \east_in_f[DATA][34] , \east_in_f[DATA][33] , \east_in_f[DATA][32] , 
        \east_in_f[DATA][31] , \east_in_f[DATA][30] , \east_in_f[DATA][29] , 
        \east_in_f[DATA][28] , \east_in_f[DATA][27] , \east_in_f[DATA][26] , 
        \east_in_f[DATA][25] , \east_in_f[DATA][24] , \east_in_f[DATA][23] , 
        \east_in_f[DATA][22] , \east_in_f[DATA][21] , \east_in_f[DATA][20] , 
        \east_in_f[DATA][19] , \east_in_f[DATA][18] , \east_in_f[DATA][17] , 
        \east_in_f[DATA][16] , \east_in_f[DATA][15] , \east_in_f[DATA][14] , 
        \east_in_f[DATA][13] , \east_in_f[DATA][12] , \east_in_f[DATA][11] , 
        \east_in_f[DATA][10] , \east_in_f[DATA][9] , \east_in_f[DATA][8] , 
        \east_in_f[DATA][7] , \east_in_f[DATA][6] , \east_in_f[DATA][5] , 
        \east_in_f[DATA][4] , \east_in_f[DATA][3] , \east_in_f[DATA][2] , 
        \east_in_f[DATA][1] , \east_in_f[DATA][0] }), .east_in_b(
        \east_in_b[ACK] ), .south_in_f({\south_in_f[REQ] , 
        \south_in_f[DATA][34] , \south_in_f[DATA][33] , \south_in_f[DATA][32] , 
        \south_in_f[DATA][31] , \south_in_f[DATA][30] , \south_in_f[DATA][29] , 
        \south_in_f[DATA][28] , \south_in_f[DATA][27] , \south_in_f[DATA][26] , 
        \south_in_f[DATA][25] , \south_in_f[DATA][24] , \south_in_f[DATA][23] , 
        \south_in_f[DATA][22] , \south_in_f[DATA][21] , \south_in_f[DATA][20] , 
        \south_in_f[DATA][19] , \south_in_f[DATA][18] , \south_in_f[DATA][17] , 
        \south_in_f[DATA][16] , \south_in_f[DATA][15] , \south_in_f[DATA][14] , 
        \south_in_f[DATA][13] , \south_in_f[DATA][12] , \south_in_f[DATA][11] , 
        \south_in_f[DATA][10] , \south_in_f[DATA][9] , \south_in_f[DATA][8] , 
        \south_in_f[DATA][7] , \south_in_f[DATA][6] , \south_in_f[DATA][5] , 
        \south_in_f[DATA][4] , \south_in_f[DATA][3] , \south_in_f[DATA][2] , 
        \south_in_f[DATA][1] , \south_in_f[DATA][0] }), .south_in_b(
        \south_in_b[ACK] ), .west_in_f({\west_in_f[REQ] , 
        \west_in_f[DATA][34] , \west_in_f[DATA][33] , \west_in_f[DATA][32] , 
        \west_in_f[DATA][31] , \west_in_f[DATA][30] , \west_in_f[DATA][29] , 
        \west_in_f[DATA][28] , \west_in_f[DATA][27] , \west_in_f[DATA][26] , 
        \west_in_f[DATA][25] , \west_in_f[DATA][24] , \west_in_f[DATA][23] , 
        \west_in_f[DATA][22] , \west_in_f[DATA][21] , \west_in_f[DATA][20] , 
        \west_in_f[DATA][19] , \west_in_f[DATA][18] , \west_in_f[DATA][17] , 
        \west_in_f[DATA][16] , \west_in_f[DATA][15] , \west_in_f[DATA][14] , 
        \west_in_f[DATA][13] , \west_in_f[DATA][12] , \west_in_f[DATA][11] , 
        \west_in_f[DATA][10] , \west_in_f[DATA][9] , \west_in_f[DATA][8] , 
        \west_in_f[DATA][7] , \west_in_f[DATA][6] , \west_in_f[DATA][5] , 
        \west_in_f[DATA][4] , \west_in_f[DATA][3] , \west_in_f[DATA][2] , 
        \west_in_f[DATA][1] , \west_in_f[DATA][0] }), .west_in_b(
        \west_in_b[ACK] ), .resource_in_f({\resource_in_f[REQ] , 
        \resource_in_f[DATA][34] , \resource_in_f[DATA][33] , 
        \resource_in_f[DATA][32] , \resource_in_f[DATA][31] , 
        \resource_in_f[DATA][30] , \resource_in_f[DATA][29] , 
        \resource_in_f[DATA][28] , \resource_in_f[DATA][27] , 
        \resource_in_f[DATA][26] , \resource_in_f[DATA][25] , 
        \resource_in_f[DATA][24] , \resource_in_f[DATA][23] , 
        \resource_in_f[DATA][22] , \resource_in_f[DATA][21] , 
        \resource_in_f[DATA][20] , \resource_in_f[DATA][19] , 
        \resource_in_f[DATA][18] , \resource_in_f[DATA][17] , 
        \resource_in_f[DATA][16] , \resource_in_f[DATA][15] , 
        \resource_in_f[DATA][14] , \resource_in_f[DATA][13] , 
        \resource_in_f[DATA][12] , \resource_in_f[DATA][11] , 
        \resource_in_f[DATA][10] , \resource_in_f[DATA][9] , 
        \resource_in_f[DATA][8] , \resource_in_f[DATA][7] , 
        \resource_in_f[DATA][6] , \resource_in_f[DATA][5] , 
        \resource_in_f[DATA][4] , \resource_in_f[DATA][3] , 
        \resource_in_f[DATA][2] , \resource_in_f[DATA][1] , 
        \resource_in_f[DATA][0] }), .resource_in_b(\resource_in_b[ACK] ), 
    .north_out_f({\north_out_f[REQ] , \north_out_f[DATA][34] , 
        \north_out_f[DATA][33] , \north_out_f[DATA][32] , 
        \north_out_f[DATA][31] , \north_out_f[DATA][30] , 
        \north_out_f[DATA][29] , \north_out_f[DATA][28] , 
        \north_out_f[DATA][27] , \north_out_f[DATA][26] , 
        \north_out_f[DATA][25] , \north_out_f[DATA][24] , 
        \north_out_f[DATA][23] , \north_out_f[DATA][22] , 
        \north_out_f[DATA][21] , \north_out_f[DATA][20] , 
        \north_out_f[DATA][19] , \north_out_f[DATA][18] , 
        \north_out_f[DATA][17] , \north_out_f[DATA][16] , 
        \north_out_f[DATA][15] , \north_out_f[DATA][14] , 
        \north_out_f[DATA][13] , \north_out_f[DATA][12] , 
        \north_out_f[DATA][11] , \north_out_f[DATA][10] , 
        \north_out_f[DATA][9] , \north_out_f[DATA][8] , \north_out_f[DATA][7] , 
        \north_out_f[DATA][6] , \north_out_f[DATA][5] , \north_out_f[DATA][4] , 
        \north_out_f[DATA][3] , \north_out_f[DATA][2] , \north_out_f[DATA][1] , 
        \north_out_f[DATA][0] }), .north_out_b(\north_out_b[ACK] ), 
    .east_out_f({\east_out_f[REQ] , \east_out_f[DATA][34] , 
        \east_out_f[DATA][33] , \east_out_f[DATA][32] , \east_out_f[DATA][31] , 
        \east_out_f[DATA][30] , \east_out_f[DATA][29] , \east_out_f[DATA][28] , 
        \east_out_f[DATA][27] , \east_out_f[DATA][26] , \east_out_f[DATA][25] , 
        \east_out_f[DATA][24] , \east_out_f[DATA][23] , \east_out_f[DATA][22] , 
        \east_out_f[DATA][21] , \east_out_f[DATA][20] , \east_out_f[DATA][19] , 
        \east_out_f[DATA][18] , \east_out_f[DATA][17] , \east_out_f[DATA][16] , 
        \east_out_f[DATA][15] , \east_out_f[DATA][14] , \east_out_f[DATA][13] , 
        \east_out_f[DATA][12] , \east_out_f[DATA][11] , \east_out_f[DATA][10] , 
        \east_out_f[DATA][9] , \east_out_f[DATA][8] , \east_out_f[DATA][7] , 
        \east_out_f[DATA][6] , \east_out_f[DATA][5] , \east_out_f[DATA][4] , 
        \east_out_f[DATA][3] , \east_out_f[DATA][2] , \east_out_f[DATA][1] , 
        \east_out_f[DATA][0] }), .east_out_b(\east_out_b[ACK] ), 
    .south_out_f({\south_out_f[REQ] , \south_out_f[DATA][34] , 
        \south_out_f[DATA][33] , \south_out_f[DATA][32] , 
        \south_out_f[DATA][31] , \south_out_f[DATA][30] , 
        \south_out_f[DATA][29] , \south_out_f[DATA][28] , 
        \south_out_f[DATA][27] , \south_out_f[DATA][26] , 
        \south_out_f[DATA][25] , \south_out_f[DATA][24] , 
        \south_out_f[DATA][23] , \south_out_f[DATA][22] , 
        \south_out_f[DATA][21] , \south_out_f[DATA][20] , 
        \south_out_f[DATA][19] , \south_out_f[DATA][18] , 
        \south_out_f[DATA][17] , \south_out_f[DATA][16] , 
        \south_out_f[DATA][15] , \south_out_f[DATA][14] , 
        \south_out_f[DATA][13] , \south_out_f[DATA][12] , 
        \south_out_f[DATA][11] , \south_out_f[DATA][10] , 
        \south_out_f[DATA][9] , \south_out_f[DATA][8] , \south_out_f[DATA][7] , 
        \south_out_f[DATA][6] , \south_out_f[DATA][5] , \south_out_f[DATA][4] , 
        \south_out_f[DATA][3] , \south_out_f[DATA][2] , \south_out_f[DATA][1] , 
        \south_out_f[DATA][0] }), .south_out_b(\south_out_b[ACK] ), 
    .west_out_f({\west_out_f[REQ] , \west_out_f[DATA][34] , 
        \west_out_f[DATA][33] , \west_out_f[DATA][32] , \west_out_f[DATA][31] , 
        \west_out_f[DATA][30] , \west_out_f[DATA][29] , \west_out_f[DATA][28] , 
        \west_out_f[DATA][27] , \west_out_f[DATA][26] , \west_out_f[DATA][25] , 
        \west_out_f[DATA][24] , \west_out_f[DATA][23] , \west_out_f[DATA][22] , 
        \west_out_f[DATA][21] , \west_out_f[DATA][20] , \west_out_f[DATA][19] , 
        \west_out_f[DATA][18] , \west_out_f[DATA][17] , \west_out_f[DATA][16] , 
        \west_out_f[DATA][15] , \west_out_f[DATA][14] , \west_out_f[DATA][13] , 
        \west_out_f[DATA][12] , \west_out_f[DATA][11] , \west_out_f[DATA][10] , 
        \west_out_f[DATA][9] , \west_out_f[DATA][8] , \west_out_f[DATA][7] , 
        \west_out_f[DATA][6] , \west_out_f[DATA][5] , \west_out_f[DATA][4] , 
        \west_out_f[DATA][3] , \west_out_f[DATA][2] , \west_out_f[DATA][1] , 
        \west_out_f[DATA][0] }), .west_out_b(\west_out_b[ACK] ), 
    .resource_out_f({\resource_out_f[REQ] , \resource_out_f[DATA][34] , 
        \resource_out_f[DATA][33] , \resource_out_f[DATA][32] , 
        \resource_out_f[DATA][31] , \resource_out_f[DATA][30] , 
        \resource_out_f[DATA][29] , \resource_out_f[DATA][28] , 
        \resource_out_f[DATA][27] , \resource_out_f[DATA][26] , 
        \resource_out_f[DATA][25] , \resource_out_f[DATA][24] , 
        \resource_out_f[DATA][23] , \resource_out_f[DATA][22] , 
        \resource_out_f[DATA][21] , \resource_out_f[DATA][20] , 
        \resource_out_f[DATA][19] , \resource_out_f[DATA][18] , 
        \resource_out_f[DATA][17] , \resource_out_f[DATA][16] , 
        \resource_out_f[DATA][15] , \resource_out_f[DATA][14] , 
        \resource_out_f[DATA][13] , \resource_out_f[DATA][12] , 
        \resource_out_f[DATA][11] , \resource_out_f[DATA][10] , 
        \resource_out_f[DATA][9] , \resource_out_f[DATA][8] , 
        \resource_out_f[DATA][7] , \resource_out_f[DATA][6] , 
        \resource_out_f[DATA][5] , \resource_out_f[DATA][4] , 
        \resource_out_f[DATA][3] , \resource_out_f[DATA][2] , 
        \resource_out_f[DATA][1] , \resource_out_f[DATA][0] }), 
    .resource_out_b(\resource_out_b[ACK] ) );
  input preset, \north_in_f[REQ] , \north_in_f[DATA][34] ,
         \north_in_f[DATA][33] , \north_in_f[DATA][32] ,
         \north_in_f[DATA][31] , \north_in_f[DATA][30] ,
         \north_in_f[DATA][29] , \north_in_f[DATA][28] ,
         \north_in_f[DATA][27] , \north_in_f[DATA][26] ,
         \north_in_f[DATA][25] , \north_in_f[DATA][24] ,
         \north_in_f[DATA][23] , \north_in_f[DATA][22] ,
         \north_in_f[DATA][21] , \north_in_f[DATA][20] ,
         \north_in_f[DATA][19] , \north_in_f[DATA][18] ,
         \north_in_f[DATA][17] , \north_in_f[DATA][16] ,
         \north_in_f[DATA][15] , \north_in_f[DATA][14] ,
         \north_in_f[DATA][13] , \north_in_f[DATA][12] ,
         \north_in_f[DATA][11] , \north_in_f[DATA][10] , \north_in_f[DATA][9] ,
         \north_in_f[DATA][8] , \north_in_f[DATA][7] , \north_in_f[DATA][6] ,
         \north_in_f[DATA][5] , \north_in_f[DATA][4] , \north_in_f[DATA][3] ,
         \north_in_f[DATA][2] , \north_in_f[DATA][1] , \north_in_f[DATA][0] ,
         \east_in_f[REQ] , \east_in_f[DATA][34] , \east_in_f[DATA][33] ,
         \east_in_f[DATA][32] , \east_in_f[DATA][31] , \east_in_f[DATA][30] ,
         \east_in_f[DATA][29] , \east_in_f[DATA][28] , \east_in_f[DATA][27] ,
         \east_in_f[DATA][26] , \east_in_f[DATA][25] , \east_in_f[DATA][24] ,
         \east_in_f[DATA][23] , \east_in_f[DATA][22] , \east_in_f[DATA][21] ,
         \east_in_f[DATA][20] , \east_in_f[DATA][19] , \east_in_f[DATA][18] ,
         \east_in_f[DATA][17] , \east_in_f[DATA][16] , \east_in_f[DATA][15] ,
         \east_in_f[DATA][14] , \east_in_f[DATA][13] , \east_in_f[DATA][12] ,
         \east_in_f[DATA][11] , \east_in_f[DATA][10] , \east_in_f[DATA][9] ,
         \east_in_f[DATA][8] , \east_in_f[DATA][7] , \east_in_f[DATA][6] ,
         \east_in_f[DATA][5] , \east_in_f[DATA][4] , \east_in_f[DATA][3] ,
         \east_in_f[DATA][2] , \east_in_f[DATA][1] , \east_in_f[DATA][0] ,
         \south_in_f[REQ] , \south_in_f[DATA][34] , \south_in_f[DATA][33] ,
         \south_in_f[DATA][32] , \south_in_f[DATA][31] ,
         \south_in_f[DATA][30] , \south_in_f[DATA][29] ,
         \south_in_f[DATA][28] , \south_in_f[DATA][27] ,
         \south_in_f[DATA][26] , \south_in_f[DATA][25] ,
         \south_in_f[DATA][24] , \south_in_f[DATA][23] ,
         \south_in_f[DATA][22] , \south_in_f[DATA][21] ,
         \south_in_f[DATA][20] , \south_in_f[DATA][19] ,
         \south_in_f[DATA][18] , \south_in_f[DATA][17] ,
         \south_in_f[DATA][16] , \south_in_f[DATA][15] ,
         \south_in_f[DATA][14] , \south_in_f[DATA][13] ,
         \south_in_f[DATA][12] , \south_in_f[DATA][11] ,
         \south_in_f[DATA][10] , \south_in_f[DATA][9] , \south_in_f[DATA][8] ,
         \south_in_f[DATA][7] , \south_in_f[DATA][6] , \south_in_f[DATA][5] ,
         \south_in_f[DATA][4] , \south_in_f[DATA][3] , \south_in_f[DATA][2] ,
         \south_in_f[DATA][1] , \south_in_f[DATA][0] , \west_in_f[REQ] ,
         \west_in_f[DATA][34] , \west_in_f[DATA][33] , \west_in_f[DATA][32] ,
         \west_in_f[DATA][31] , \west_in_f[DATA][30] , \west_in_f[DATA][29] ,
         \west_in_f[DATA][28] , \west_in_f[DATA][27] , \west_in_f[DATA][26] ,
         \west_in_f[DATA][25] , \west_in_f[DATA][24] , \west_in_f[DATA][23] ,
         \west_in_f[DATA][22] , \west_in_f[DATA][21] , \west_in_f[DATA][20] ,
         \west_in_f[DATA][19] , \west_in_f[DATA][18] , \west_in_f[DATA][17] ,
         \west_in_f[DATA][16] , \west_in_f[DATA][15] , \west_in_f[DATA][14] ,
         \west_in_f[DATA][13] , \west_in_f[DATA][12] , \west_in_f[DATA][11] ,
         \west_in_f[DATA][10] , \west_in_f[DATA][9] , \west_in_f[DATA][8] ,
         \west_in_f[DATA][7] , \west_in_f[DATA][6] , \west_in_f[DATA][5] ,
         \west_in_f[DATA][4] , \west_in_f[DATA][3] , \west_in_f[DATA][2] ,
         \west_in_f[DATA][1] , \west_in_f[DATA][0] , \resource_in_f[REQ] ,
         \resource_in_f[DATA][34] , \resource_in_f[DATA][33] ,
         \resource_in_f[DATA][32] , \resource_in_f[DATA][31] ,
         \resource_in_f[DATA][30] , \resource_in_f[DATA][29] ,
         \resource_in_f[DATA][28] , \resource_in_f[DATA][27] ,
         \resource_in_f[DATA][26] , \resource_in_f[DATA][25] ,
         \resource_in_f[DATA][24] , \resource_in_f[DATA][23] ,
         \resource_in_f[DATA][22] , \resource_in_f[DATA][21] ,
         \resource_in_f[DATA][20] , \resource_in_f[DATA][19] ,
         \resource_in_f[DATA][18] , \resource_in_f[DATA][17] ,
         \resource_in_f[DATA][16] , \resource_in_f[DATA][15] ,
         \resource_in_f[DATA][14] , \resource_in_f[DATA][13] ,
         \resource_in_f[DATA][12] , \resource_in_f[DATA][11] ,
         \resource_in_f[DATA][10] , \resource_in_f[DATA][9] ,
         \resource_in_f[DATA][8] , \resource_in_f[DATA][7] ,
         \resource_in_f[DATA][6] , \resource_in_f[DATA][5] ,
         \resource_in_f[DATA][4] , \resource_in_f[DATA][3] ,
         \resource_in_f[DATA][2] , \resource_in_f[DATA][1] ,
         \resource_in_f[DATA][0] , \north_out_b[ACK] , \east_out_b[ACK] ,
         \south_out_b[ACK] , \west_out_b[ACK] , \resource_out_b[ACK] ;
  output \north_in_b[ACK] , \east_in_b[ACK] , \south_in_b[ACK] ,
         \west_in_b[ACK] , \resource_in_b[ACK] , \north_out_f[REQ] ,
         \north_out_f[DATA][34] , \north_out_f[DATA][33] ,
         \north_out_f[DATA][32] , \north_out_f[DATA][31] ,
         \north_out_f[DATA][30] , \north_out_f[DATA][29] ,
         \north_out_f[DATA][28] , \north_out_f[DATA][27] ,
         \north_out_f[DATA][26] , \north_out_f[DATA][25] ,
         \north_out_f[DATA][24] , \north_out_f[DATA][23] ,
         \north_out_f[DATA][22] , \north_out_f[DATA][21] ,
         \north_out_f[DATA][20] , \north_out_f[DATA][19] ,
         \north_out_f[DATA][18] , \north_out_f[DATA][17] ,
         \north_out_f[DATA][16] , \north_out_f[DATA][15] ,
         \north_out_f[DATA][14] , \north_out_f[DATA][13] ,
         \north_out_f[DATA][12] , \north_out_f[DATA][11] ,
         \north_out_f[DATA][10] , \north_out_f[DATA][9] ,
         \north_out_f[DATA][8] , \north_out_f[DATA][7] ,
         \north_out_f[DATA][6] , \north_out_f[DATA][5] ,
         \north_out_f[DATA][4] , \north_out_f[DATA][3] ,
         \north_out_f[DATA][2] , \north_out_f[DATA][1] ,
         \north_out_f[DATA][0] , \east_out_f[REQ] , \east_out_f[DATA][34] ,
         \east_out_f[DATA][33] , \east_out_f[DATA][32] ,
         \east_out_f[DATA][31] , \east_out_f[DATA][30] ,
         \east_out_f[DATA][29] , \east_out_f[DATA][28] ,
         \east_out_f[DATA][27] , \east_out_f[DATA][26] ,
         \east_out_f[DATA][25] , \east_out_f[DATA][24] ,
         \east_out_f[DATA][23] , \east_out_f[DATA][22] ,
         \east_out_f[DATA][21] , \east_out_f[DATA][20] ,
         \east_out_f[DATA][19] , \east_out_f[DATA][18] ,
         \east_out_f[DATA][17] , \east_out_f[DATA][16] ,
         \east_out_f[DATA][15] , \east_out_f[DATA][14] ,
         \east_out_f[DATA][13] , \east_out_f[DATA][12] ,
         \east_out_f[DATA][11] , \east_out_f[DATA][10] , \east_out_f[DATA][9] ,
         \east_out_f[DATA][8] , \east_out_f[DATA][7] , \east_out_f[DATA][6] ,
         \east_out_f[DATA][5] , \east_out_f[DATA][4] , \east_out_f[DATA][3] ,
         \east_out_f[DATA][2] , \east_out_f[DATA][1] , \east_out_f[DATA][0] ,
         \south_out_f[REQ] , \south_out_f[DATA][34] , \south_out_f[DATA][33] ,
         \south_out_f[DATA][32] , \south_out_f[DATA][31] ,
         \south_out_f[DATA][30] , \south_out_f[DATA][29] ,
         \south_out_f[DATA][28] , \south_out_f[DATA][27] ,
         \south_out_f[DATA][26] , \south_out_f[DATA][25] ,
         \south_out_f[DATA][24] , \south_out_f[DATA][23] ,
         \south_out_f[DATA][22] , \south_out_f[DATA][21] ,
         \south_out_f[DATA][20] , \south_out_f[DATA][19] ,
         \south_out_f[DATA][18] , \south_out_f[DATA][17] ,
         \south_out_f[DATA][16] , \south_out_f[DATA][15] ,
         \south_out_f[DATA][14] , \south_out_f[DATA][13] ,
         \south_out_f[DATA][12] , \south_out_f[DATA][11] ,
         \south_out_f[DATA][10] , \south_out_f[DATA][9] ,
         \south_out_f[DATA][8] , \south_out_f[DATA][7] ,
         \south_out_f[DATA][6] , \south_out_f[DATA][5] ,
         \south_out_f[DATA][4] , \south_out_f[DATA][3] ,
         \south_out_f[DATA][2] , \south_out_f[DATA][1] ,
         \south_out_f[DATA][0] , \west_out_f[REQ] , \west_out_f[DATA][34] ,
         \west_out_f[DATA][33] , \west_out_f[DATA][32] ,
         \west_out_f[DATA][31] , \west_out_f[DATA][30] ,
         \west_out_f[DATA][29] , \west_out_f[DATA][28] ,
         \west_out_f[DATA][27] , \west_out_f[DATA][26] ,
         \west_out_f[DATA][25] , \west_out_f[DATA][24] ,
         \west_out_f[DATA][23] , \west_out_f[DATA][22] ,
         \west_out_f[DATA][21] , \west_out_f[DATA][20] ,
         \west_out_f[DATA][19] , \west_out_f[DATA][18] ,
         \west_out_f[DATA][17] , \west_out_f[DATA][16] ,
         \west_out_f[DATA][15] , \west_out_f[DATA][14] ,
         \west_out_f[DATA][13] , \west_out_f[DATA][12] ,
         \west_out_f[DATA][11] , \west_out_f[DATA][10] , \west_out_f[DATA][9] ,
         \west_out_f[DATA][8] , \west_out_f[DATA][7] , \west_out_f[DATA][6] ,
         \west_out_f[DATA][5] , \west_out_f[DATA][4] , \west_out_f[DATA][3] ,
         \west_out_f[DATA][2] , \west_out_f[DATA][1] , \west_out_f[DATA][0] ,
         \resource_out_f[REQ] , \resource_out_f[DATA][34] ,
         \resource_out_f[DATA][33] , \resource_out_f[DATA][32] ,
         \resource_out_f[DATA][31] , \resource_out_f[DATA][30] ,
         \resource_out_f[DATA][29] , \resource_out_f[DATA][28] ,
         \resource_out_f[DATA][27] , \resource_out_f[DATA][26] ,
         \resource_out_f[DATA][25] , \resource_out_f[DATA][24] ,
         \resource_out_f[DATA][23] , \resource_out_f[DATA][22] ,
         \resource_out_f[DATA][21] , \resource_out_f[DATA][20] ,
         \resource_out_f[DATA][19] , \resource_out_f[DATA][18] ,
         \resource_out_f[DATA][17] , \resource_out_f[DATA][16] ,
         \resource_out_f[DATA][15] , \resource_out_f[DATA][14] ,
         \resource_out_f[DATA][13] , \resource_out_f[DATA][12] ,
         \resource_out_f[DATA][11] , \resource_out_f[DATA][10] ,
         \resource_out_f[DATA][9] , \resource_out_f[DATA][8] ,
         \resource_out_f[DATA][7] , \resource_out_f[DATA][6] ,
         \resource_out_f[DATA][5] , \resource_out_f[DATA][4] ,
         \resource_out_f[DATA][3] , \resource_out_f[DATA][2] ,
         \resource_out_f[DATA][1] , \resource_out_f[DATA][0] ;
  wire   \north_hpu_f[REQ] , \north_hpu_f[DATA][34] , \north_hpu_f[DATA][33] ,
         \north_hpu_f[DATA][32] , \north_hpu_f[DATA][31] ,
         \north_hpu_f[DATA][30] , \north_hpu_f[DATA][29] ,
         \north_hpu_f[DATA][28] , \north_hpu_f[DATA][27] ,
         \north_hpu_f[DATA][26] , \north_hpu_f[DATA][25] ,
         \north_hpu_f[DATA][24] , \north_hpu_f[DATA][23] ,
         \north_hpu_f[DATA][22] , \north_hpu_f[DATA][21] ,
         \north_hpu_f[DATA][20] , \north_hpu_f[DATA][19] ,
         \north_hpu_f[DATA][18] , \north_hpu_f[DATA][17] ,
         \north_hpu_f[DATA][16] , \north_hpu_f[DATA][15] ,
         \north_hpu_f[DATA][14] , \north_hpu_f[DATA][13] ,
         \north_hpu_f[DATA][12] , \north_hpu_f[DATA][11] ,
         \north_hpu_f[DATA][10] , \north_hpu_f[DATA][9] ,
         \north_hpu_f[DATA][8] , \north_hpu_f[DATA][7] ,
         \north_hpu_f[DATA][6] , \north_hpu_f[DATA][5] ,
         \north_hpu_f[DATA][4] , \north_hpu_f[DATA][3] ,
         \north_hpu_f[DATA][2] , \north_hpu_f[DATA][1] ,
         \north_hpu_f[DATA][0] , \north_hpu_b[ACK] , \south_hpu_f[REQ] ,
         \south_hpu_f[DATA][34] , \south_hpu_f[DATA][33] ,
         \south_hpu_f[DATA][32] , \south_hpu_f[DATA][31] ,
         \south_hpu_f[DATA][30] , \south_hpu_f[DATA][29] ,
         \south_hpu_f[DATA][28] , \south_hpu_f[DATA][27] ,
         \south_hpu_f[DATA][26] , \south_hpu_f[DATA][25] ,
         \south_hpu_f[DATA][24] , \south_hpu_f[DATA][23] ,
         \south_hpu_f[DATA][22] , \south_hpu_f[DATA][21] ,
         \south_hpu_f[DATA][20] , \south_hpu_f[DATA][19] ,
         \south_hpu_f[DATA][18] , \south_hpu_f[DATA][17] ,
         \south_hpu_f[DATA][16] , \south_hpu_f[DATA][15] ,
         \south_hpu_f[DATA][14] , \south_hpu_f[DATA][13] ,
         \south_hpu_f[DATA][12] , \south_hpu_f[DATA][11] ,
         \south_hpu_f[DATA][10] , \south_hpu_f[DATA][9] ,
         \south_hpu_f[DATA][8] , \south_hpu_f[DATA][7] ,
         \south_hpu_f[DATA][6] , \south_hpu_f[DATA][5] ,
         \south_hpu_f[DATA][4] , \south_hpu_f[DATA][3] ,
         \south_hpu_f[DATA][2] , \south_hpu_f[DATA][1] ,
         \south_hpu_f[DATA][0] , \south_hpu_b[ACK] , \east_hpu_f[REQ] ,
         \east_hpu_f[DATA][34] , \east_hpu_f[DATA][33] ,
         \east_hpu_f[DATA][32] , \east_hpu_f[DATA][31] ,
         \east_hpu_f[DATA][30] , \east_hpu_f[DATA][29] ,
         \east_hpu_f[DATA][28] , \east_hpu_f[DATA][27] ,
         \east_hpu_f[DATA][26] , \east_hpu_f[DATA][25] ,
         \east_hpu_f[DATA][24] , \east_hpu_f[DATA][23] ,
         \east_hpu_f[DATA][22] , \east_hpu_f[DATA][21] ,
         \east_hpu_f[DATA][20] , \east_hpu_f[DATA][19] ,
         \east_hpu_f[DATA][18] , \east_hpu_f[DATA][17] ,
         \east_hpu_f[DATA][16] , \east_hpu_f[DATA][15] ,
         \east_hpu_f[DATA][14] , \east_hpu_f[DATA][13] ,
         \east_hpu_f[DATA][12] , \east_hpu_f[DATA][11] ,
         \east_hpu_f[DATA][10] , \east_hpu_f[DATA][9] , \east_hpu_f[DATA][8] ,
         \east_hpu_f[DATA][7] , \east_hpu_f[DATA][6] , \east_hpu_f[DATA][5] ,
         \east_hpu_f[DATA][4] , \east_hpu_f[DATA][3] , \east_hpu_f[DATA][2] ,
         \east_hpu_f[DATA][1] , \east_hpu_f[DATA][0] , \east_hpu_b[ACK] ,
         \west_hpu_f[REQ] , \west_hpu_f[DATA][34] , \west_hpu_f[DATA][33] ,
         \west_hpu_f[DATA][32] , \west_hpu_f[DATA][31] ,
         \west_hpu_f[DATA][30] , \west_hpu_f[DATA][29] ,
         \west_hpu_f[DATA][28] , \west_hpu_f[DATA][27] ,
         \west_hpu_f[DATA][26] , \west_hpu_f[DATA][25] ,
         \west_hpu_f[DATA][24] , \west_hpu_f[DATA][23] ,
         \west_hpu_f[DATA][22] , \west_hpu_f[DATA][21] ,
         \west_hpu_f[DATA][20] , \west_hpu_f[DATA][19] ,
         \west_hpu_f[DATA][18] , \west_hpu_f[DATA][17] ,
         \west_hpu_f[DATA][16] , \west_hpu_f[DATA][15] ,
         \west_hpu_f[DATA][14] , \west_hpu_f[DATA][13] ,
         \west_hpu_f[DATA][12] , \west_hpu_f[DATA][11] ,
         \west_hpu_f[DATA][10] , \west_hpu_f[DATA][9] , \west_hpu_f[DATA][8] ,
         \west_hpu_f[DATA][7] , \west_hpu_f[DATA][6] , \west_hpu_f[DATA][5] ,
         \west_hpu_f[DATA][4] , \west_hpu_f[DATA][3] , \west_hpu_f[DATA][2] ,
         \west_hpu_f[DATA][1] , \west_hpu_f[DATA][0] , \west_hpu_b[ACK] ,
         \resource_hpu_f[REQ] , \resource_hpu_f[DATA][34] ,
         \resource_hpu_f[DATA][33] , \resource_hpu_f[DATA][32] ,
         \resource_hpu_f[DATA][31] , \resource_hpu_f[DATA][30] ,
         \resource_hpu_f[DATA][29] , \resource_hpu_f[DATA][28] ,
         \resource_hpu_f[DATA][27] , \resource_hpu_f[DATA][26] ,
         \resource_hpu_f[DATA][25] , \resource_hpu_f[DATA][24] ,
         \resource_hpu_f[DATA][23] , \resource_hpu_f[DATA][22] ,
         \resource_hpu_f[DATA][21] , \resource_hpu_f[DATA][20] ,
         \resource_hpu_f[DATA][19] , \resource_hpu_f[DATA][18] ,
         \resource_hpu_f[DATA][17] , \resource_hpu_f[DATA][16] ,
         \resource_hpu_f[DATA][15] , \resource_hpu_f[DATA][14] ,
         \resource_hpu_f[DATA][13] , \resource_hpu_f[DATA][12] ,
         \resource_hpu_f[DATA][11] , \resource_hpu_f[DATA][10] ,
         \resource_hpu_f[DATA][9] , \resource_hpu_f[DATA][8] ,
         \resource_hpu_f[DATA][7] , \resource_hpu_f[DATA][6] ,
         \resource_hpu_f[DATA][5] , \resource_hpu_f[DATA][4] ,
         \resource_hpu_f[DATA][3] , \resource_hpu_f[DATA][2] ,
         \resource_hpu_f[DATA][1] , \resource_hpu_f[DATA][0] ,
         \resource_hpu_b[ACK] , \chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] ,
         \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] ,
         \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] ,
         \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] ,
         \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] ,
         \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] ,
         \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] ,
         \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] ,
         \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] ,
         \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] ,
         \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] ,
         \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] ,
         \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] ,
         \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] ,
         \chs_in_f[4][DATA][7] , \chs_in_f[4][DATA][6] ,
         \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] ,
         \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] ,
         \chs_in_f[4][DATA][1] , \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] ,
         \chs_in_f[3][DATA][34] , \chs_in_f[3][DATA][33] ,
         \chs_in_f[3][DATA][32] , \chs_in_f[3][DATA][31] ,
         \chs_in_f[3][DATA][30] , \chs_in_f[3][DATA][29] ,
         \chs_in_f[3][DATA][28] , \chs_in_f[3][DATA][27] ,
         \chs_in_f[3][DATA][26] , \chs_in_f[3][DATA][25] ,
         \chs_in_f[3][DATA][24] , \chs_in_f[3][DATA][23] ,
         \chs_in_f[3][DATA][22] , \chs_in_f[3][DATA][21] ,
         \chs_in_f[3][DATA][20] , \chs_in_f[3][DATA][19] ,
         \chs_in_f[3][DATA][18] , \chs_in_f[3][DATA][17] ,
         \chs_in_f[3][DATA][16] , \chs_in_f[3][DATA][15] ,
         \chs_in_f[3][DATA][14] , \chs_in_f[3][DATA][13] ,
         \chs_in_f[3][DATA][12] , \chs_in_f[3][DATA][11] ,
         \chs_in_f[3][DATA][10] , \chs_in_f[3][DATA][9] ,
         \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] ,
         \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] ,
         \chs_in_f[3][DATA][4] , \chs_in_f[3][DATA][3] ,
         \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] ,
         \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] ,
         \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] ,
         \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] ,
         \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] ,
         \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] ,
         \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] ,
         \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] ,
         \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] ,
         \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] ,
         \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] ,
         \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] ,
         \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] ,
         \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] ,
         \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] ,
         \chs_in_f[2][DATA][7] , \chs_in_f[2][DATA][6] ,
         \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] ,
         \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] ,
         \chs_in_f[2][DATA][1] , \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] ,
         \chs_in_f[1][DATA][34] , \chs_in_f[1][DATA][33] ,
         \chs_in_f[1][DATA][32] , \chs_in_f[1][DATA][31] ,
         \chs_in_f[1][DATA][30] , \chs_in_f[1][DATA][29] ,
         \chs_in_f[1][DATA][28] , \chs_in_f[1][DATA][27] ,
         \chs_in_f[1][DATA][26] , \chs_in_f[1][DATA][25] ,
         \chs_in_f[1][DATA][24] , \chs_in_f[1][DATA][23] ,
         \chs_in_f[1][DATA][22] , \chs_in_f[1][DATA][21] ,
         \chs_in_f[1][DATA][20] , \chs_in_f[1][DATA][19] ,
         \chs_in_f[1][DATA][18] , \chs_in_f[1][DATA][17] ,
         \chs_in_f[1][DATA][16] , \chs_in_f[1][DATA][15] ,
         \chs_in_f[1][DATA][14] , \chs_in_f[1][DATA][13] ,
         \chs_in_f[1][DATA][12] , \chs_in_f[1][DATA][11] ,
         \chs_in_f[1][DATA][10] , \chs_in_f[1][DATA][9] ,
         \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] ,
         \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] ,
         \chs_in_f[1][DATA][4] , \chs_in_f[1][DATA][3] ,
         \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] ,
         \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] ,
         \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] ,
         \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] ,
         \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] ,
         \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] ,
         \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] ,
         \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] ,
         \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] ,
         \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] ,
         \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] ,
         \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] ,
         \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] ,
         \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] ,
         \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] ,
         \chs_in_f[0][DATA][7] , \chs_in_f[0][DATA][6] ,
         \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] ,
         \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] ,
         \chs_in_f[0][DATA][1] , \chs_in_f[0][DATA][0] , \chs_in_b[4][ACK] ,
         \chs_in_b[3][ACK] , \chs_in_b[2][ACK] , \chs_in_b[1][ACK] ,
         \chs_in_b[0][ACK] , \switch_sel[4][4] , \switch_sel[4][3] ,
         \switch_sel[4][2] , \switch_sel[4][1] , \switch_sel[4][0] ,
         \switch_sel[3][4] , \switch_sel[3][3] , \switch_sel[3][2] ,
         \switch_sel[3][1] , \switch_sel[3][0] , \switch_sel[2][4] ,
         \switch_sel[2][3] , \switch_sel[2][2] , \switch_sel[2][1] ,
         \switch_sel[2][0] , \switch_sel[1][4] , \switch_sel[1][3] ,
         \switch_sel[1][2] , \switch_sel[1][1] , \switch_sel[1][0] ,
         \switch_sel[0][4] , \switch_sel[0][3] , \switch_sel[0][2] ,
         \switch_sel[0][1] , \switch_sel[0][0] , n2, n3;

  channel_latch_1_xxxxxxxxx_35 north_in_latch ( .preset(n3), .left_in({
        \north_in_f[REQ] , \north_in_f[DATA][34] , \north_in_f[DATA][33] , 
        \north_in_f[DATA][32] , \north_in_f[DATA][31] , \north_in_f[DATA][30] , 
        \north_in_f[DATA][29] , \north_in_f[DATA][28] , \north_in_f[DATA][27] , 
        \north_in_f[DATA][26] , \north_in_f[DATA][25] , \north_in_f[DATA][24] , 
        \north_in_f[DATA][23] , \north_in_f[DATA][22] , \north_in_f[DATA][21] , 
        \north_in_f[DATA][20] , \north_in_f[DATA][19] , \north_in_f[DATA][18] , 
        \north_in_f[DATA][17] , \north_in_f[DATA][16] , \north_in_f[DATA][15] , 
        \north_in_f[DATA][14] , \north_in_f[DATA][13] , \north_in_f[DATA][12] , 
        \north_in_f[DATA][11] , \north_in_f[DATA][10] , \north_in_f[DATA][9] , 
        \north_in_f[DATA][8] , \north_in_f[DATA][7] , \north_in_f[DATA][6] , 
        \north_in_f[DATA][5] , \north_in_f[DATA][4] , \north_in_f[DATA][3] , 
        \north_in_f[DATA][2] , \north_in_f[DATA][1] , \north_in_f[DATA][0] }), 
        .left_out(\north_in_b[ACK] ), .right_out({\north_hpu_f[REQ] , 
        \north_hpu_f[DATA][34] , \north_hpu_f[DATA][33] , 
        \north_hpu_f[DATA][32] , \north_hpu_f[DATA][31] , 
        \north_hpu_f[DATA][30] , \north_hpu_f[DATA][29] , 
        \north_hpu_f[DATA][28] , \north_hpu_f[DATA][27] , 
        \north_hpu_f[DATA][26] , \north_hpu_f[DATA][25] , 
        \north_hpu_f[DATA][24] , \north_hpu_f[DATA][23] , 
        \north_hpu_f[DATA][22] , \north_hpu_f[DATA][21] , 
        \north_hpu_f[DATA][20] , \north_hpu_f[DATA][19] , 
        \north_hpu_f[DATA][18] , \north_hpu_f[DATA][17] , 
        \north_hpu_f[DATA][16] , \north_hpu_f[DATA][15] , 
        \north_hpu_f[DATA][14] , \north_hpu_f[DATA][13] , 
        \north_hpu_f[DATA][12] , \north_hpu_f[DATA][11] , 
        \north_hpu_f[DATA][10] , \north_hpu_f[DATA][9] , 
        \north_hpu_f[DATA][8] , \north_hpu_f[DATA][7] , \north_hpu_f[DATA][6] , 
        \north_hpu_f[DATA][5] , \north_hpu_f[DATA][4] , \north_hpu_f[DATA][3] , 
        \north_hpu_f[DATA][2] , \north_hpu_f[DATA][1] , \north_hpu_f[DATA][0] }), .right_in(\north_hpu_b[ACK] ) );
  channel_latch_1_xxxxxxxxx_34 south_in_latch ( .preset(n3), .left_in({
        \south_in_f[REQ] , \south_in_f[DATA][34] , \south_in_f[DATA][33] , 
        \south_in_f[DATA][32] , \south_in_f[DATA][31] , \south_in_f[DATA][30] , 
        \south_in_f[DATA][29] , \south_in_f[DATA][28] , \south_in_f[DATA][27] , 
        \south_in_f[DATA][26] , \south_in_f[DATA][25] , \south_in_f[DATA][24] , 
        \south_in_f[DATA][23] , \south_in_f[DATA][22] , \south_in_f[DATA][21] , 
        \south_in_f[DATA][20] , \south_in_f[DATA][19] , \south_in_f[DATA][18] , 
        \south_in_f[DATA][17] , \south_in_f[DATA][16] , \south_in_f[DATA][15] , 
        \south_in_f[DATA][14] , \south_in_f[DATA][13] , \south_in_f[DATA][12] , 
        \south_in_f[DATA][11] , \south_in_f[DATA][10] , \south_in_f[DATA][9] , 
        \south_in_f[DATA][8] , \south_in_f[DATA][7] , \south_in_f[DATA][6] , 
        \south_in_f[DATA][5] , \south_in_f[DATA][4] , \south_in_f[DATA][3] , 
        \south_in_f[DATA][2] , \south_in_f[DATA][1] , \south_in_f[DATA][0] }), 
        .left_out(\south_in_b[ACK] ), .right_out({\south_hpu_f[REQ] , 
        \south_hpu_f[DATA][34] , \south_hpu_f[DATA][33] , 
        \south_hpu_f[DATA][32] , \south_hpu_f[DATA][31] , 
        \south_hpu_f[DATA][30] , \south_hpu_f[DATA][29] , 
        \south_hpu_f[DATA][28] , \south_hpu_f[DATA][27] , 
        \south_hpu_f[DATA][26] , \south_hpu_f[DATA][25] , 
        \south_hpu_f[DATA][24] , \south_hpu_f[DATA][23] , 
        \south_hpu_f[DATA][22] , \south_hpu_f[DATA][21] , 
        \south_hpu_f[DATA][20] , \south_hpu_f[DATA][19] , 
        \south_hpu_f[DATA][18] , \south_hpu_f[DATA][17] , 
        \south_hpu_f[DATA][16] , \south_hpu_f[DATA][15] , 
        \south_hpu_f[DATA][14] , \south_hpu_f[DATA][13] , 
        \south_hpu_f[DATA][12] , \south_hpu_f[DATA][11] , 
        \south_hpu_f[DATA][10] , \south_hpu_f[DATA][9] , 
        \south_hpu_f[DATA][8] , \south_hpu_f[DATA][7] , \south_hpu_f[DATA][6] , 
        \south_hpu_f[DATA][5] , \south_hpu_f[DATA][4] , \south_hpu_f[DATA][3] , 
        \south_hpu_f[DATA][2] , \south_hpu_f[DATA][1] , \south_hpu_f[DATA][0] }), .right_in(\south_hpu_b[ACK] ) );
  channel_latch_1_xxxxxxxxx_33 east_in_latch ( .preset(n3), .left_in({
        \east_in_f[REQ] , \east_in_f[DATA][34] , \east_in_f[DATA][33] , 
        \east_in_f[DATA][32] , \east_in_f[DATA][31] , \east_in_f[DATA][30] , 
        \east_in_f[DATA][29] , \east_in_f[DATA][28] , \east_in_f[DATA][27] , 
        \east_in_f[DATA][26] , \east_in_f[DATA][25] , \east_in_f[DATA][24] , 
        \east_in_f[DATA][23] , \east_in_f[DATA][22] , \east_in_f[DATA][21] , 
        \east_in_f[DATA][20] , \east_in_f[DATA][19] , \east_in_f[DATA][18] , 
        \east_in_f[DATA][17] , \east_in_f[DATA][16] , \east_in_f[DATA][15] , 
        \east_in_f[DATA][14] , \east_in_f[DATA][13] , \east_in_f[DATA][12] , 
        \east_in_f[DATA][11] , \east_in_f[DATA][10] , \east_in_f[DATA][9] , 
        \east_in_f[DATA][8] , \east_in_f[DATA][7] , \east_in_f[DATA][6] , 
        \east_in_f[DATA][5] , \east_in_f[DATA][4] , \east_in_f[DATA][3] , 
        \east_in_f[DATA][2] , \east_in_f[DATA][1] , \east_in_f[DATA][0] }), 
        .left_out(\east_in_b[ACK] ), .right_out({\east_hpu_f[REQ] , 
        \east_hpu_f[DATA][34] , \east_hpu_f[DATA][33] , \east_hpu_f[DATA][32] , 
        \east_hpu_f[DATA][31] , \east_hpu_f[DATA][30] , \east_hpu_f[DATA][29] , 
        \east_hpu_f[DATA][28] , \east_hpu_f[DATA][27] , \east_hpu_f[DATA][26] , 
        \east_hpu_f[DATA][25] , \east_hpu_f[DATA][24] , \east_hpu_f[DATA][23] , 
        \east_hpu_f[DATA][22] , \east_hpu_f[DATA][21] , \east_hpu_f[DATA][20] , 
        \east_hpu_f[DATA][19] , \east_hpu_f[DATA][18] , \east_hpu_f[DATA][17] , 
        \east_hpu_f[DATA][16] , \east_hpu_f[DATA][15] , \east_hpu_f[DATA][14] , 
        \east_hpu_f[DATA][13] , \east_hpu_f[DATA][12] , \east_hpu_f[DATA][11] , 
        \east_hpu_f[DATA][10] , \east_hpu_f[DATA][9] , \east_hpu_f[DATA][8] , 
        \east_hpu_f[DATA][7] , \east_hpu_f[DATA][6] , \east_hpu_f[DATA][5] , 
        \east_hpu_f[DATA][4] , \east_hpu_f[DATA][3] , \east_hpu_f[DATA][2] , 
        \east_hpu_f[DATA][1] , \east_hpu_f[DATA][0] }), .right_in(
        \east_hpu_b[ACK] ) );
  channel_latch_1_xxxxxxxxx_32 west_in_latch ( .preset(n3), .left_in({
        \west_in_f[REQ] , \west_in_f[DATA][34] , \west_in_f[DATA][33] , 
        \west_in_f[DATA][32] , \west_in_f[DATA][31] , \west_in_f[DATA][30] , 
        \west_in_f[DATA][29] , \west_in_f[DATA][28] , \west_in_f[DATA][27] , 
        \west_in_f[DATA][26] , \west_in_f[DATA][25] , \west_in_f[DATA][24] , 
        \west_in_f[DATA][23] , \west_in_f[DATA][22] , \west_in_f[DATA][21] , 
        \west_in_f[DATA][20] , \west_in_f[DATA][19] , \west_in_f[DATA][18] , 
        \west_in_f[DATA][17] , \west_in_f[DATA][16] , \west_in_f[DATA][15] , 
        \west_in_f[DATA][14] , \west_in_f[DATA][13] , \west_in_f[DATA][12] , 
        \west_in_f[DATA][11] , \west_in_f[DATA][10] , \west_in_f[DATA][9] , 
        \west_in_f[DATA][8] , \west_in_f[DATA][7] , \west_in_f[DATA][6] , 
        \west_in_f[DATA][5] , \west_in_f[DATA][4] , \west_in_f[DATA][3] , 
        \west_in_f[DATA][2] , \west_in_f[DATA][1] , \west_in_f[DATA][0] }), 
        .left_out(\west_in_b[ACK] ), .right_out({\west_hpu_f[REQ] , 
        \west_hpu_f[DATA][34] , \west_hpu_f[DATA][33] , \west_hpu_f[DATA][32] , 
        \west_hpu_f[DATA][31] , \west_hpu_f[DATA][30] , \west_hpu_f[DATA][29] , 
        \west_hpu_f[DATA][28] , \west_hpu_f[DATA][27] , \west_hpu_f[DATA][26] , 
        \west_hpu_f[DATA][25] , \west_hpu_f[DATA][24] , \west_hpu_f[DATA][23] , 
        \west_hpu_f[DATA][22] , \west_hpu_f[DATA][21] , \west_hpu_f[DATA][20] , 
        \west_hpu_f[DATA][19] , \west_hpu_f[DATA][18] , \west_hpu_f[DATA][17] , 
        \west_hpu_f[DATA][16] , \west_hpu_f[DATA][15] , \west_hpu_f[DATA][14] , 
        \west_hpu_f[DATA][13] , \west_hpu_f[DATA][12] , \west_hpu_f[DATA][11] , 
        \west_hpu_f[DATA][10] , \west_hpu_f[DATA][9] , \west_hpu_f[DATA][8] , 
        \west_hpu_f[DATA][7] , \west_hpu_f[DATA][6] , \west_hpu_f[DATA][5] , 
        \west_hpu_f[DATA][4] , \west_hpu_f[DATA][3] , \west_hpu_f[DATA][2] , 
        \west_hpu_f[DATA][1] , \west_hpu_f[DATA][0] }), .right_in(
        \west_hpu_b[ACK] ) );
  channel_latch_1_xxxxxxxxx_31 resource_in_latch ( .preset(n3), .left_in({
        \resource_in_f[REQ] , \resource_in_f[DATA][34] , 
        \resource_in_f[DATA][33] , \resource_in_f[DATA][32] , 
        \resource_in_f[DATA][31] , \resource_in_f[DATA][30] , 
        \resource_in_f[DATA][29] , \resource_in_f[DATA][28] , 
        \resource_in_f[DATA][27] , \resource_in_f[DATA][26] , 
        \resource_in_f[DATA][25] , \resource_in_f[DATA][24] , 
        \resource_in_f[DATA][23] , \resource_in_f[DATA][22] , 
        \resource_in_f[DATA][21] , \resource_in_f[DATA][20] , 
        \resource_in_f[DATA][19] , \resource_in_f[DATA][18] , 
        \resource_in_f[DATA][17] , \resource_in_f[DATA][16] , 
        \resource_in_f[DATA][15] , \resource_in_f[DATA][14] , 
        \resource_in_f[DATA][13] , \resource_in_f[DATA][12] , 
        \resource_in_f[DATA][11] , \resource_in_f[DATA][10] , 
        \resource_in_f[DATA][9] , \resource_in_f[DATA][8] , 
        \resource_in_f[DATA][7] , \resource_in_f[DATA][6] , 
        \resource_in_f[DATA][5] , \resource_in_f[DATA][4] , 
        \resource_in_f[DATA][3] , \resource_in_f[DATA][2] , 
        \resource_in_f[DATA][1] , \resource_in_f[DATA][0] }), .left_out(
        \resource_in_b[ACK] ), .right_out({\resource_hpu_f[REQ] , 
        \resource_hpu_f[DATA][34] , \resource_hpu_f[DATA][33] , 
        \resource_hpu_f[DATA][32] , \resource_hpu_f[DATA][31] , 
        \resource_hpu_f[DATA][30] , \resource_hpu_f[DATA][29] , 
        \resource_hpu_f[DATA][28] , \resource_hpu_f[DATA][27] , 
        \resource_hpu_f[DATA][26] , \resource_hpu_f[DATA][25] , 
        \resource_hpu_f[DATA][24] , \resource_hpu_f[DATA][23] , 
        \resource_hpu_f[DATA][22] , \resource_hpu_f[DATA][21] , 
        \resource_hpu_f[DATA][20] , \resource_hpu_f[DATA][19] , 
        \resource_hpu_f[DATA][18] , \resource_hpu_f[DATA][17] , 
        \resource_hpu_f[DATA][16] , \resource_hpu_f[DATA][15] , 
        \resource_hpu_f[DATA][14] , \resource_hpu_f[DATA][13] , 
        \resource_hpu_f[DATA][12] , \resource_hpu_f[DATA][11] , 
        \resource_hpu_f[DATA][10] , \resource_hpu_f[DATA][9] , 
        \resource_hpu_f[DATA][8] , \resource_hpu_f[DATA][7] , 
        \resource_hpu_f[DATA][6] , \resource_hpu_f[DATA][5] , 
        \resource_hpu_f[DATA][4] , \resource_hpu_f[DATA][3] , 
        \resource_hpu_f[DATA][2] , \resource_hpu_f[DATA][1] , 
        \resource_hpu_f[DATA][0] }), .right_in(\resource_hpu_b[ACK] ) );
  hpu_0_0_3 north_hpu ( .preset(n2), .chan_in_f({\north_hpu_f[REQ] , 
        \north_hpu_f[DATA][34] , \north_hpu_f[DATA][33] , 
        \north_hpu_f[DATA][32] , \north_hpu_f[DATA][31] , 
        \north_hpu_f[DATA][30] , \north_hpu_f[DATA][29] , 
        \north_hpu_f[DATA][28] , \north_hpu_f[DATA][27] , 
        \north_hpu_f[DATA][26] , \north_hpu_f[DATA][25] , 
        \north_hpu_f[DATA][24] , \north_hpu_f[DATA][23] , 
        \north_hpu_f[DATA][22] , \north_hpu_f[DATA][21] , 
        \north_hpu_f[DATA][20] , \north_hpu_f[DATA][19] , 
        \north_hpu_f[DATA][18] , \north_hpu_f[DATA][17] , 
        \north_hpu_f[DATA][16] , \north_hpu_f[DATA][15] , 
        \north_hpu_f[DATA][14] , \north_hpu_f[DATA][13] , 
        \north_hpu_f[DATA][12] , \north_hpu_f[DATA][11] , 
        \north_hpu_f[DATA][10] , \north_hpu_f[DATA][9] , 
        \north_hpu_f[DATA][8] , \north_hpu_f[DATA][7] , \north_hpu_f[DATA][6] , 
        \north_hpu_f[DATA][5] , \north_hpu_f[DATA][4] , \north_hpu_f[DATA][3] , 
        \north_hpu_f[DATA][2] , \north_hpu_f[DATA][1] , \north_hpu_f[DATA][0] }), .chan_in_b(\north_hpu_b[ACK] ), .chan_out_f({\chs_in_f[0][REQ] , 
        \chs_in_f[0][DATA][34] , \chs_in_f[0][DATA][33] , 
        \chs_in_f[0][DATA][32] , \chs_in_f[0][DATA][31] , 
        \chs_in_f[0][DATA][30] , \chs_in_f[0][DATA][29] , 
        \chs_in_f[0][DATA][28] , \chs_in_f[0][DATA][27] , 
        \chs_in_f[0][DATA][26] , \chs_in_f[0][DATA][25] , 
        \chs_in_f[0][DATA][24] , \chs_in_f[0][DATA][23] , 
        \chs_in_f[0][DATA][22] , \chs_in_f[0][DATA][21] , 
        \chs_in_f[0][DATA][20] , \chs_in_f[0][DATA][19] , 
        \chs_in_f[0][DATA][18] , \chs_in_f[0][DATA][17] , 
        \chs_in_f[0][DATA][16] , \chs_in_f[0][DATA][15] , 
        \chs_in_f[0][DATA][14] , \chs_in_f[0][DATA][13] , 
        \chs_in_f[0][DATA][12] , \chs_in_f[0][DATA][11] , 
        \chs_in_f[0][DATA][10] , \chs_in_f[0][DATA][9] , 
        \chs_in_f[0][DATA][8] , \chs_in_f[0][DATA][7] , \chs_in_f[0][DATA][6] , 
        \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] , \chs_in_f[0][DATA][3] , 
        \chs_in_f[0][DATA][2] , \chs_in_f[0][DATA][1] , \chs_in_f[0][DATA][0] }), .chan_out_b(\chs_in_b[0][ACK] ), .sel({\switch_sel[0][4] , 
        \switch_sel[0][3] , \switch_sel[0][2] , \switch_sel[0][1] , 
        \switch_sel[0][0] }) );
  hpu_0_2_3 south_hpu ( .preset(n2), .chan_in_f({\south_hpu_f[REQ] , 
        \south_hpu_f[DATA][34] , \south_hpu_f[DATA][33] , 
        \south_hpu_f[DATA][32] , \south_hpu_f[DATA][31] , 
        \south_hpu_f[DATA][30] , \south_hpu_f[DATA][29] , 
        \south_hpu_f[DATA][28] , \south_hpu_f[DATA][27] , 
        \south_hpu_f[DATA][26] , \south_hpu_f[DATA][25] , 
        \south_hpu_f[DATA][24] , \south_hpu_f[DATA][23] , 
        \south_hpu_f[DATA][22] , \south_hpu_f[DATA][21] , 
        \south_hpu_f[DATA][20] , \south_hpu_f[DATA][19] , 
        \south_hpu_f[DATA][18] , \south_hpu_f[DATA][17] , 
        \south_hpu_f[DATA][16] , \south_hpu_f[DATA][15] , 
        \south_hpu_f[DATA][14] , \south_hpu_f[DATA][13] , 
        \south_hpu_f[DATA][12] , \south_hpu_f[DATA][11] , 
        \south_hpu_f[DATA][10] , \south_hpu_f[DATA][9] , 
        \south_hpu_f[DATA][8] , \south_hpu_f[DATA][7] , \south_hpu_f[DATA][6] , 
        \south_hpu_f[DATA][5] , \south_hpu_f[DATA][4] , \south_hpu_f[DATA][3] , 
        \south_hpu_f[DATA][2] , \south_hpu_f[DATA][1] , \south_hpu_f[DATA][0] }), .chan_in_b(\south_hpu_b[ACK] ), .chan_out_f({\chs_in_f[2][REQ] , 
        \chs_in_f[2][DATA][34] , \chs_in_f[2][DATA][33] , 
        \chs_in_f[2][DATA][32] , \chs_in_f[2][DATA][31] , 
        \chs_in_f[2][DATA][30] , \chs_in_f[2][DATA][29] , 
        \chs_in_f[2][DATA][28] , \chs_in_f[2][DATA][27] , 
        \chs_in_f[2][DATA][26] , \chs_in_f[2][DATA][25] , 
        \chs_in_f[2][DATA][24] , \chs_in_f[2][DATA][23] , 
        \chs_in_f[2][DATA][22] , \chs_in_f[2][DATA][21] , 
        \chs_in_f[2][DATA][20] , \chs_in_f[2][DATA][19] , 
        \chs_in_f[2][DATA][18] , \chs_in_f[2][DATA][17] , 
        \chs_in_f[2][DATA][16] , \chs_in_f[2][DATA][15] , 
        \chs_in_f[2][DATA][14] , \chs_in_f[2][DATA][13] , 
        \chs_in_f[2][DATA][12] , \chs_in_f[2][DATA][11] , 
        \chs_in_f[2][DATA][10] , \chs_in_f[2][DATA][9] , 
        \chs_in_f[2][DATA][8] , \chs_in_f[2][DATA][7] , \chs_in_f[2][DATA][6] , 
        \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] , \chs_in_f[2][DATA][3] , 
        \chs_in_f[2][DATA][2] , \chs_in_f[2][DATA][1] , \chs_in_f[2][DATA][0] }), .chan_out_b(\chs_in_b[2][ACK] ), .sel({\switch_sel[2][4] , 
        \switch_sel[2][3] , \switch_sel[2][2] , \switch_sel[2][1] , 
        \switch_sel[2][0] }) );
  hpu_0_1_3 east_hpu ( .preset(n2), .chan_in_f({\east_hpu_f[REQ] , 
        \east_hpu_f[DATA][34] , \east_hpu_f[DATA][33] , \east_hpu_f[DATA][32] , 
        \east_hpu_f[DATA][31] , \east_hpu_f[DATA][30] , \east_hpu_f[DATA][29] , 
        \east_hpu_f[DATA][28] , \east_hpu_f[DATA][27] , \east_hpu_f[DATA][26] , 
        \east_hpu_f[DATA][25] , \east_hpu_f[DATA][24] , \east_hpu_f[DATA][23] , 
        \east_hpu_f[DATA][22] , \east_hpu_f[DATA][21] , \east_hpu_f[DATA][20] , 
        \east_hpu_f[DATA][19] , \east_hpu_f[DATA][18] , \east_hpu_f[DATA][17] , 
        \east_hpu_f[DATA][16] , \east_hpu_f[DATA][15] , \east_hpu_f[DATA][14] , 
        \east_hpu_f[DATA][13] , \east_hpu_f[DATA][12] , \east_hpu_f[DATA][11] , 
        \east_hpu_f[DATA][10] , \east_hpu_f[DATA][9] , \east_hpu_f[DATA][8] , 
        \east_hpu_f[DATA][7] , \east_hpu_f[DATA][6] , \east_hpu_f[DATA][5] , 
        \east_hpu_f[DATA][4] , \east_hpu_f[DATA][3] , \east_hpu_f[DATA][2] , 
        \east_hpu_f[DATA][1] , \east_hpu_f[DATA][0] }), .chan_in_b(
        \east_hpu_b[ACK] ), .chan_out_f({\chs_in_f[1][REQ] , 
        \chs_in_f[1][DATA][34] , \chs_in_f[1][DATA][33] , 
        \chs_in_f[1][DATA][32] , \chs_in_f[1][DATA][31] , 
        \chs_in_f[1][DATA][30] , \chs_in_f[1][DATA][29] , 
        \chs_in_f[1][DATA][28] , \chs_in_f[1][DATA][27] , 
        \chs_in_f[1][DATA][26] , \chs_in_f[1][DATA][25] , 
        \chs_in_f[1][DATA][24] , \chs_in_f[1][DATA][23] , 
        \chs_in_f[1][DATA][22] , \chs_in_f[1][DATA][21] , 
        \chs_in_f[1][DATA][20] , \chs_in_f[1][DATA][19] , 
        \chs_in_f[1][DATA][18] , \chs_in_f[1][DATA][17] , 
        \chs_in_f[1][DATA][16] , \chs_in_f[1][DATA][15] , 
        \chs_in_f[1][DATA][14] , \chs_in_f[1][DATA][13] , 
        \chs_in_f[1][DATA][12] , \chs_in_f[1][DATA][11] , 
        \chs_in_f[1][DATA][10] , \chs_in_f[1][DATA][9] , 
        \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] , \chs_in_f[1][DATA][6] , 
        \chs_in_f[1][DATA][5] , \chs_in_f[1][DATA][4] , \chs_in_f[1][DATA][3] , 
        \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] , \chs_in_f[1][DATA][0] }), .chan_out_b(\chs_in_b[1][ACK] ), .sel({\switch_sel[1][4] , 
        \switch_sel[1][3] , \switch_sel[1][2] , \switch_sel[1][1] , 
        \switch_sel[1][0] }) );
  hpu_0_3_3 west_hpu ( .preset(n2), .chan_in_f({\west_hpu_f[REQ] , 
        \west_hpu_f[DATA][34] , \west_hpu_f[DATA][33] , \west_hpu_f[DATA][32] , 
        \west_hpu_f[DATA][31] , \west_hpu_f[DATA][30] , \west_hpu_f[DATA][29] , 
        \west_hpu_f[DATA][28] , \west_hpu_f[DATA][27] , \west_hpu_f[DATA][26] , 
        \west_hpu_f[DATA][25] , \west_hpu_f[DATA][24] , \west_hpu_f[DATA][23] , 
        \west_hpu_f[DATA][22] , \west_hpu_f[DATA][21] , \west_hpu_f[DATA][20] , 
        \west_hpu_f[DATA][19] , \west_hpu_f[DATA][18] , \west_hpu_f[DATA][17] , 
        \west_hpu_f[DATA][16] , \west_hpu_f[DATA][15] , \west_hpu_f[DATA][14] , 
        \west_hpu_f[DATA][13] , \west_hpu_f[DATA][12] , \west_hpu_f[DATA][11] , 
        \west_hpu_f[DATA][10] , \west_hpu_f[DATA][9] , \west_hpu_f[DATA][8] , 
        \west_hpu_f[DATA][7] , \west_hpu_f[DATA][6] , \west_hpu_f[DATA][5] , 
        \west_hpu_f[DATA][4] , \west_hpu_f[DATA][3] , \west_hpu_f[DATA][2] , 
        \west_hpu_f[DATA][1] , \west_hpu_f[DATA][0] }), .chan_in_b(
        \west_hpu_b[ACK] ), .chan_out_f({\chs_in_f[3][REQ] , 
        \chs_in_f[3][DATA][34] , \chs_in_f[3][DATA][33] , 
        \chs_in_f[3][DATA][32] , \chs_in_f[3][DATA][31] , 
        \chs_in_f[3][DATA][30] , \chs_in_f[3][DATA][29] , 
        \chs_in_f[3][DATA][28] , \chs_in_f[3][DATA][27] , 
        \chs_in_f[3][DATA][26] , \chs_in_f[3][DATA][25] , 
        \chs_in_f[3][DATA][24] , \chs_in_f[3][DATA][23] , 
        \chs_in_f[3][DATA][22] , \chs_in_f[3][DATA][21] , 
        \chs_in_f[3][DATA][20] , \chs_in_f[3][DATA][19] , 
        \chs_in_f[3][DATA][18] , \chs_in_f[3][DATA][17] , 
        \chs_in_f[3][DATA][16] , \chs_in_f[3][DATA][15] , 
        \chs_in_f[3][DATA][14] , \chs_in_f[3][DATA][13] , 
        \chs_in_f[3][DATA][12] , \chs_in_f[3][DATA][11] , 
        \chs_in_f[3][DATA][10] , \chs_in_f[3][DATA][9] , 
        \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] , \chs_in_f[3][DATA][6] , 
        \chs_in_f[3][DATA][5] , \chs_in_f[3][DATA][4] , \chs_in_f[3][DATA][3] , 
        \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] , \chs_in_f[3][DATA][0] }), .chan_out_b(\chs_in_b[3][ACK] ), .sel({\switch_sel[3][4] , 
        \switch_sel[3][3] , \switch_sel[3][2] , \switch_sel[3][1] , 
        \switch_sel[3][0] }) );
  hpu_1_x_3 resource_hpu ( .preset(n2), .chan_in_f({\resource_hpu_f[REQ] , 
        \resource_hpu_f[DATA][34] , \resource_hpu_f[DATA][33] , 
        \resource_hpu_f[DATA][32] , \resource_hpu_f[DATA][31] , 
        \resource_hpu_f[DATA][30] , \resource_hpu_f[DATA][29] , 
        \resource_hpu_f[DATA][28] , \resource_hpu_f[DATA][27] , 
        \resource_hpu_f[DATA][26] , \resource_hpu_f[DATA][25] , 
        \resource_hpu_f[DATA][24] , \resource_hpu_f[DATA][23] , 
        \resource_hpu_f[DATA][22] , \resource_hpu_f[DATA][21] , 
        \resource_hpu_f[DATA][20] , \resource_hpu_f[DATA][19] , 
        \resource_hpu_f[DATA][18] , \resource_hpu_f[DATA][17] , 
        \resource_hpu_f[DATA][16] , \resource_hpu_f[DATA][15] , 
        \resource_hpu_f[DATA][14] , \resource_hpu_f[DATA][13] , 
        \resource_hpu_f[DATA][12] , \resource_hpu_f[DATA][11] , 
        \resource_hpu_f[DATA][10] , \resource_hpu_f[DATA][9] , 
        \resource_hpu_f[DATA][8] , \resource_hpu_f[DATA][7] , 
        \resource_hpu_f[DATA][6] , \resource_hpu_f[DATA][5] , 
        \resource_hpu_f[DATA][4] , \resource_hpu_f[DATA][3] , 
        \resource_hpu_f[DATA][2] , \resource_hpu_f[DATA][1] , 
        \resource_hpu_f[DATA][0] }), .chan_in_b(\resource_hpu_b[ACK] ), 
        .chan_out_f({\chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] , 
        \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] , 
        \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] , 
        \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] , 
        \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] , 
        \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] , 
        \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] , 
        \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] , 
        \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] , 
        \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] , 
        \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] , 
        \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] , 
        \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] , 
        \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] , \chs_in_f[4][DATA][7] , 
        \chs_in_f[4][DATA][6] , \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] , 
        \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] , \chs_in_f[4][DATA][1] , 
        \chs_in_f[4][DATA][0] }), .chan_out_b(\chs_in_b[4][ACK] ), .sel({
        \switch_sel[4][4] , \switch_sel[4][3] , \switch_sel[4][2] , 
        \switch_sel[4][1] , \switch_sel[4][0] }) );
  crossbar_stage_3 xbar_with_latches ( .preset(n3), .switch_sel({1'b0, 
        \switch_sel[4][3] , \switch_sel[4][2] , \switch_sel[4][1] , 
        \switch_sel[4][0] , \switch_sel[3][4] , 1'b0, \switch_sel[3][2] , 
        \switch_sel[3][1] , \switch_sel[3][0] , \switch_sel[2][4] , 
        \switch_sel[2][3] , 1'b0, \switch_sel[2][1] , \switch_sel[2][0] , 
        \switch_sel[1][4] , \switch_sel[1][3] , \switch_sel[1][2] , 1'b0, 
        \switch_sel[1][0] , \switch_sel[0][4] , \switch_sel[0][3] , 
        \switch_sel[0][2] , \switch_sel[0][1] , 1'b0}), .chs_in_f({
        \chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] , \chs_in_f[4][DATA][33] , 
        \chs_in_f[4][DATA][32] , \chs_in_f[4][DATA][31] , 
        \chs_in_f[4][DATA][30] , \chs_in_f[4][DATA][29] , 
        \chs_in_f[4][DATA][28] , \chs_in_f[4][DATA][27] , 
        \chs_in_f[4][DATA][26] , \chs_in_f[4][DATA][25] , 
        \chs_in_f[4][DATA][24] , \chs_in_f[4][DATA][23] , 
        \chs_in_f[4][DATA][22] , \chs_in_f[4][DATA][21] , 
        \chs_in_f[4][DATA][20] , \chs_in_f[4][DATA][19] , 
        \chs_in_f[4][DATA][18] , \chs_in_f[4][DATA][17] , 
        \chs_in_f[4][DATA][16] , \chs_in_f[4][DATA][15] , 
        \chs_in_f[4][DATA][14] , \chs_in_f[4][DATA][13] , 
        \chs_in_f[4][DATA][12] , \chs_in_f[4][DATA][11] , 
        \chs_in_f[4][DATA][10] , \chs_in_f[4][DATA][9] , 
        \chs_in_f[4][DATA][8] , \chs_in_f[4][DATA][7] , \chs_in_f[4][DATA][6] , 
        \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] , \chs_in_f[4][DATA][3] , 
        \chs_in_f[4][DATA][2] , \chs_in_f[4][DATA][1] , \chs_in_f[4][DATA][0] , 
        \chs_in_f[3][REQ] , \chs_in_f[3][DATA][34] , \chs_in_f[3][DATA][33] , 
        \chs_in_f[3][DATA][32] , \chs_in_f[3][DATA][31] , 
        \chs_in_f[3][DATA][30] , \chs_in_f[3][DATA][29] , 
        \chs_in_f[3][DATA][28] , \chs_in_f[3][DATA][27] , 
        \chs_in_f[3][DATA][26] , \chs_in_f[3][DATA][25] , 
        \chs_in_f[3][DATA][24] , \chs_in_f[3][DATA][23] , 
        \chs_in_f[3][DATA][22] , \chs_in_f[3][DATA][21] , 
        \chs_in_f[3][DATA][20] , \chs_in_f[3][DATA][19] , 
        \chs_in_f[3][DATA][18] , \chs_in_f[3][DATA][17] , 
        \chs_in_f[3][DATA][16] , \chs_in_f[3][DATA][15] , 
        \chs_in_f[3][DATA][14] , \chs_in_f[3][DATA][13] , 
        \chs_in_f[3][DATA][12] , \chs_in_f[3][DATA][11] , 
        \chs_in_f[3][DATA][10] , \chs_in_f[3][DATA][9] , 
        \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] , \chs_in_f[3][DATA][6] , 
        \chs_in_f[3][DATA][5] , \chs_in_f[3][DATA][4] , \chs_in_f[3][DATA][3] , 
        \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] , \chs_in_f[3][DATA][0] , 
        \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] , \chs_in_f[2][DATA][33] , 
        \chs_in_f[2][DATA][32] , \chs_in_f[2][DATA][31] , 
        \chs_in_f[2][DATA][30] , \chs_in_f[2][DATA][29] , 
        \chs_in_f[2][DATA][28] , \chs_in_f[2][DATA][27] , 
        \chs_in_f[2][DATA][26] , \chs_in_f[2][DATA][25] , 
        \chs_in_f[2][DATA][24] , \chs_in_f[2][DATA][23] , 
        \chs_in_f[2][DATA][22] , \chs_in_f[2][DATA][21] , 
        \chs_in_f[2][DATA][20] , \chs_in_f[2][DATA][19] , 
        \chs_in_f[2][DATA][18] , \chs_in_f[2][DATA][17] , 
        \chs_in_f[2][DATA][16] , \chs_in_f[2][DATA][15] , 
        \chs_in_f[2][DATA][14] , \chs_in_f[2][DATA][13] , 
        \chs_in_f[2][DATA][12] , \chs_in_f[2][DATA][11] , 
        \chs_in_f[2][DATA][10] , \chs_in_f[2][DATA][9] , 
        \chs_in_f[2][DATA][8] , \chs_in_f[2][DATA][7] , \chs_in_f[2][DATA][6] , 
        \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] , \chs_in_f[2][DATA][3] , 
        \chs_in_f[2][DATA][2] , \chs_in_f[2][DATA][1] , \chs_in_f[2][DATA][0] , 
        \chs_in_f[1][REQ] , \chs_in_f[1][DATA][34] , \chs_in_f[1][DATA][33] , 
        \chs_in_f[1][DATA][32] , \chs_in_f[1][DATA][31] , 
        \chs_in_f[1][DATA][30] , \chs_in_f[1][DATA][29] , 
        \chs_in_f[1][DATA][28] , \chs_in_f[1][DATA][27] , 
        \chs_in_f[1][DATA][26] , \chs_in_f[1][DATA][25] , 
        \chs_in_f[1][DATA][24] , \chs_in_f[1][DATA][23] , 
        \chs_in_f[1][DATA][22] , \chs_in_f[1][DATA][21] , 
        \chs_in_f[1][DATA][20] , \chs_in_f[1][DATA][19] , 
        \chs_in_f[1][DATA][18] , \chs_in_f[1][DATA][17] , 
        \chs_in_f[1][DATA][16] , \chs_in_f[1][DATA][15] , 
        \chs_in_f[1][DATA][14] , \chs_in_f[1][DATA][13] , 
        \chs_in_f[1][DATA][12] , \chs_in_f[1][DATA][11] , 
        \chs_in_f[1][DATA][10] , \chs_in_f[1][DATA][9] , 
        \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] , \chs_in_f[1][DATA][6] , 
        \chs_in_f[1][DATA][5] , \chs_in_f[1][DATA][4] , \chs_in_f[1][DATA][3] , 
        \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] , \chs_in_f[1][DATA][0] , 
        \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] , \chs_in_f[0][DATA][33] , 
        \chs_in_f[0][DATA][32] , \chs_in_f[0][DATA][31] , 
        \chs_in_f[0][DATA][30] , \chs_in_f[0][DATA][29] , 
        \chs_in_f[0][DATA][28] , \chs_in_f[0][DATA][27] , 
        \chs_in_f[0][DATA][26] , \chs_in_f[0][DATA][25] , 
        \chs_in_f[0][DATA][24] , \chs_in_f[0][DATA][23] , 
        \chs_in_f[0][DATA][22] , \chs_in_f[0][DATA][21] , 
        \chs_in_f[0][DATA][20] , \chs_in_f[0][DATA][19] , 
        \chs_in_f[0][DATA][18] , \chs_in_f[0][DATA][17] , 
        \chs_in_f[0][DATA][16] , \chs_in_f[0][DATA][15] , 
        \chs_in_f[0][DATA][14] , \chs_in_f[0][DATA][13] , 
        \chs_in_f[0][DATA][12] , \chs_in_f[0][DATA][11] , 
        \chs_in_f[0][DATA][10] , \chs_in_f[0][DATA][9] , 
        \chs_in_f[0][DATA][8] , \chs_in_f[0][DATA][7] , \chs_in_f[0][DATA][6] , 
        \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] , \chs_in_f[0][DATA][3] , 
        \chs_in_f[0][DATA][2] , \chs_in_f[0][DATA][1] , \chs_in_f[0][DATA][0] }), .chs_in_b({\chs_in_b[4][ACK] , \chs_in_b[3][ACK] , \chs_in_b[2][ACK] , 
        \chs_in_b[1][ACK] , \chs_in_b[0][ACK] }), .latches_out_f({
        \resource_out_f[REQ] , \resource_out_f[DATA][34] , 
        \resource_out_f[DATA][33] , \resource_out_f[DATA][32] , 
        \resource_out_f[DATA][31] , \resource_out_f[DATA][30] , 
        \resource_out_f[DATA][29] , \resource_out_f[DATA][28] , 
        \resource_out_f[DATA][27] , \resource_out_f[DATA][26] , 
        \resource_out_f[DATA][25] , \resource_out_f[DATA][24] , 
        \resource_out_f[DATA][23] , \resource_out_f[DATA][22] , 
        \resource_out_f[DATA][21] , \resource_out_f[DATA][20] , 
        \resource_out_f[DATA][19] , \resource_out_f[DATA][18] , 
        \resource_out_f[DATA][17] , \resource_out_f[DATA][16] , 
        \resource_out_f[DATA][15] , \resource_out_f[DATA][14] , 
        \resource_out_f[DATA][13] , \resource_out_f[DATA][12] , 
        \resource_out_f[DATA][11] , \resource_out_f[DATA][10] , 
        \resource_out_f[DATA][9] , \resource_out_f[DATA][8] , 
        \resource_out_f[DATA][7] , \resource_out_f[DATA][6] , 
        \resource_out_f[DATA][5] , \resource_out_f[DATA][4] , 
        \resource_out_f[DATA][3] , \resource_out_f[DATA][2] , 
        \resource_out_f[DATA][1] , \resource_out_f[DATA][0] , 
        \west_out_f[REQ] , \west_out_f[DATA][34] , \west_out_f[DATA][33] , 
        \west_out_f[DATA][32] , \west_out_f[DATA][31] , \west_out_f[DATA][30] , 
        \west_out_f[DATA][29] , \west_out_f[DATA][28] , \west_out_f[DATA][27] , 
        \west_out_f[DATA][26] , \west_out_f[DATA][25] , \west_out_f[DATA][24] , 
        \west_out_f[DATA][23] , \west_out_f[DATA][22] , \west_out_f[DATA][21] , 
        \west_out_f[DATA][20] , \west_out_f[DATA][19] , \west_out_f[DATA][18] , 
        \west_out_f[DATA][17] , \west_out_f[DATA][16] , \west_out_f[DATA][15] , 
        \west_out_f[DATA][14] , \west_out_f[DATA][13] , \west_out_f[DATA][12] , 
        \west_out_f[DATA][11] , \west_out_f[DATA][10] , \west_out_f[DATA][9] , 
        \west_out_f[DATA][8] , \west_out_f[DATA][7] , \west_out_f[DATA][6] , 
        \west_out_f[DATA][5] , \west_out_f[DATA][4] , \west_out_f[DATA][3] , 
        \west_out_f[DATA][2] , \west_out_f[DATA][1] , \west_out_f[DATA][0] , 
        \south_out_f[REQ] , \south_out_f[DATA][34] , \south_out_f[DATA][33] , 
        \south_out_f[DATA][32] , \south_out_f[DATA][31] , 
        \south_out_f[DATA][30] , \south_out_f[DATA][29] , 
        \south_out_f[DATA][28] , \south_out_f[DATA][27] , 
        \south_out_f[DATA][26] , \south_out_f[DATA][25] , 
        \south_out_f[DATA][24] , \south_out_f[DATA][23] , 
        \south_out_f[DATA][22] , \south_out_f[DATA][21] , 
        \south_out_f[DATA][20] , \south_out_f[DATA][19] , 
        \south_out_f[DATA][18] , \south_out_f[DATA][17] , 
        \south_out_f[DATA][16] , \south_out_f[DATA][15] , 
        \south_out_f[DATA][14] , \south_out_f[DATA][13] , 
        \south_out_f[DATA][12] , \south_out_f[DATA][11] , 
        \south_out_f[DATA][10] , \south_out_f[DATA][9] , 
        \south_out_f[DATA][8] , \south_out_f[DATA][7] , \south_out_f[DATA][6] , 
        \south_out_f[DATA][5] , \south_out_f[DATA][4] , \south_out_f[DATA][3] , 
        \south_out_f[DATA][2] , \south_out_f[DATA][1] , \south_out_f[DATA][0] , 
        \east_out_f[REQ] , \east_out_f[DATA][34] , \east_out_f[DATA][33] , 
        \east_out_f[DATA][32] , \east_out_f[DATA][31] , \east_out_f[DATA][30] , 
        \east_out_f[DATA][29] , \east_out_f[DATA][28] , \east_out_f[DATA][27] , 
        \east_out_f[DATA][26] , \east_out_f[DATA][25] , \east_out_f[DATA][24] , 
        \east_out_f[DATA][23] , \east_out_f[DATA][22] , \east_out_f[DATA][21] , 
        \east_out_f[DATA][20] , \east_out_f[DATA][19] , \east_out_f[DATA][18] , 
        \east_out_f[DATA][17] , \east_out_f[DATA][16] , \east_out_f[DATA][15] , 
        \east_out_f[DATA][14] , \east_out_f[DATA][13] , \east_out_f[DATA][12] , 
        \east_out_f[DATA][11] , \east_out_f[DATA][10] , \east_out_f[DATA][9] , 
        \east_out_f[DATA][8] , \east_out_f[DATA][7] , \east_out_f[DATA][6] , 
        \east_out_f[DATA][5] , \east_out_f[DATA][4] , \east_out_f[DATA][3] , 
        \east_out_f[DATA][2] , \east_out_f[DATA][1] , \east_out_f[DATA][0] , 
        \north_out_f[REQ] , \north_out_f[DATA][34] , \north_out_f[DATA][33] , 
        \north_out_f[DATA][32] , \north_out_f[DATA][31] , 
        \north_out_f[DATA][30] , \north_out_f[DATA][29] , 
        \north_out_f[DATA][28] , \north_out_f[DATA][27] , 
        \north_out_f[DATA][26] , \north_out_f[DATA][25] , 
        \north_out_f[DATA][24] , \north_out_f[DATA][23] , 
        \north_out_f[DATA][22] , \north_out_f[DATA][21] , 
        \north_out_f[DATA][20] , \north_out_f[DATA][19] , 
        \north_out_f[DATA][18] , \north_out_f[DATA][17] , 
        \north_out_f[DATA][16] , \north_out_f[DATA][15] , 
        \north_out_f[DATA][14] , \north_out_f[DATA][13] , 
        \north_out_f[DATA][12] , \north_out_f[DATA][11] , 
        \north_out_f[DATA][10] , \north_out_f[DATA][9] , 
        \north_out_f[DATA][8] , \north_out_f[DATA][7] , \north_out_f[DATA][6] , 
        \north_out_f[DATA][5] , \north_out_f[DATA][4] , \north_out_f[DATA][3] , 
        \north_out_f[DATA][2] , \north_out_f[DATA][1] , \north_out_f[DATA][0] }), .latches_out_b({\resource_out_b[ACK] , \west_out_b[ACK] , 
        \south_out_b[ACK] , \east_out_b[ACK] , \north_out_b[ACK] }) );
  HS65_LS_BFX9 U1 ( .A(preset), .Z(n3) );
  HS65_LS_BFX9 U2 ( .A(preset), .Z(n2) );
endmodule


module noc_node_3 ( p_clk, n_clk, reset, .proc_in({\proc_in[MCMD][1] , 
        \proc_in[MCMD][0] , \proc_in[MADDR][31] , \proc_in[MADDR][30] , 
        \proc_in[MADDR][29] , \proc_in[MADDR][28] , \proc_in[MADDR][27] , 
        \proc_in[MADDR][26] , \proc_in[MADDR][25] , \proc_in[MADDR][24] , 
        \proc_in[MADDR][23] , \proc_in[MADDR][22] , \proc_in[MADDR][21] , 
        \proc_in[MADDR][20] , \proc_in[MADDR][19] , \proc_in[MADDR][18] , 
        \proc_in[MADDR][17] , \proc_in[MADDR][16] , \proc_in[MADDR][15] , 
        \proc_in[MADDR][14] , \proc_in[MADDR][13] , \proc_in[MADDR][12] , 
        \proc_in[MADDR][11] , \proc_in[MADDR][10] , \proc_in[MADDR][9] , 
        \proc_in[MADDR][8] , \proc_in[MADDR][7] , \proc_in[MADDR][6] , 
        \proc_in[MADDR][5] , \proc_in[MADDR][4] , \proc_in[MADDR][3] , 
        \proc_in[MADDR][2] , \proc_in[MADDR][1] , \proc_in[MADDR][0] , 
        \proc_in[MDATA][31] , \proc_in[MDATA][30] , \proc_in[MDATA][29] , 
        \proc_in[MDATA][28] , \proc_in[MDATA][27] , \proc_in[MDATA][26] , 
        \proc_in[MDATA][25] , \proc_in[MDATA][24] , \proc_in[MDATA][23] , 
        \proc_in[MDATA][22] , \proc_in[MDATA][21] , \proc_in[MDATA][20] , 
        \proc_in[MDATA][19] , \proc_in[MDATA][18] , \proc_in[MDATA][17] , 
        \proc_in[MDATA][16] , \proc_in[MDATA][15] , \proc_in[MDATA][14] , 
        \proc_in[MDATA][13] , \proc_in[MDATA][12] , \proc_in[MDATA][11] , 
        \proc_in[MDATA][10] , \proc_in[MDATA][9] , \proc_in[MDATA][8] , 
        \proc_in[MDATA][7] , \proc_in[MDATA][6] , \proc_in[MDATA][5] , 
        \proc_in[MDATA][4] , \proc_in[MDATA][3] , \proc_in[MDATA][2] , 
        \proc_in[MDATA][1] , \proc_in[MDATA][0] }), .proc_out({
        \proc_out[SCMDACCEPT] , \proc_out[SRESP] , \proc_out[SDATA][31] , 
        \proc_out[SDATA][30] , \proc_out[SDATA][29] , \proc_out[SDATA][28] , 
        \proc_out[SDATA][27] , \proc_out[SDATA][26] , \proc_out[SDATA][25] , 
        \proc_out[SDATA][24] , \proc_out[SDATA][23] , \proc_out[SDATA][22] , 
        \proc_out[SDATA][21] , \proc_out[SDATA][20] , \proc_out[SDATA][19] , 
        \proc_out[SDATA][18] , \proc_out[SDATA][17] , \proc_out[SDATA][16] , 
        \proc_out[SDATA][15] , \proc_out[SDATA][14] , \proc_out[SDATA][13] , 
        \proc_out[SDATA][12] , \proc_out[SDATA][11] , \proc_out[SDATA][10] , 
        \proc_out[SDATA][9] , \proc_out[SDATA][8] , \proc_out[SDATA][7] , 
        \proc_out[SDATA][6] , \proc_out[SDATA][5] , \proc_out[SDATA][4] , 
        \proc_out[SDATA][3] , \proc_out[SDATA][2] , \proc_out[SDATA][1] , 
        \proc_out[SDATA][0] }), .spm_in({\spm_in[SCMDACCEPT] , \spm_in[SRESP] , 
        \spm_in[SDATA][63] , \spm_in[SDATA][62] , \spm_in[SDATA][61] , 
        \spm_in[SDATA][60] , \spm_in[SDATA][59] , \spm_in[SDATA][58] , 
        \spm_in[SDATA][57] , \spm_in[SDATA][56] , \spm_in[SDATA][55] , 
        \spm_in[SDATA][54] , \spm_in[SDATA][53] , \spm_in[SDATA][52] , 
        \spm_in[SDATA][51] , \spm_in[SDATA][50] , \spm_in[SDATA][49] , 
        \spm_in[SDATA][48] , \spm_in[SDATA][47] , \spm_in[SDATA][46] , 
        \spm_in[SDATA][45] , \spm_in[SDATA][44] , \spm_in[SDATA][43] , 
        \spm_in[SDATA][42] , \spm_in[SDATA][41] , \spm_in[SDATA][40] , 
        \spm_in[SDATA][39] , \spm_in[SDATA][38] , \spm_in[SDATA][37] , 
        \spm_in[SDATA][36] , \spm_in[SDATA][35] , \spm_in[SDATA][34] , 
        \spm_in[SDATA][33] , \spm_in[SDATA][32] , \spm_in[SDATA][31] , 
        \spm_in[SDATA][30] , \spm_in[SDATA][29] , \spm_in[SDATA][28] , 
        \spm_in[SDATA][27] , \spm_in[SDATA][26] , \spm_in[SDATA][25] , 
        \spm_in[SDATA][24] , \spm_in[SDATA][23] , \spm_in[SDATA][22] , 
        \spm_in[SDATA][21] , \spm_in[SDATA][20] , \spm_in[SDATA][19] , 
        \spm_in[SDATA][18] , \spm_in[SDATA][17] , \spm_in[SDATA][16] , 
        \spm_in[SDATA][15] , \spm_in[SDATA][14] , \spm_in[SDATA][13] , 
        \spm_in[SDATA][12] , \spm_in[SDATA][11] , \spm_in[SDATA][10] , 
        \spm_in[SDATA][9] , \spm_in[SDATA][8] , \spm_in[SDATA][7] , 
        \spm_in[SDATA][6] , \spm_in[SDATA][5] , \spm_in[SDATA][4] , 
        \spm_in[SDATA][3] , \spm_in[SDATA][2] , \spm_in[SDATA][1] , 
        \spm_in[SDATA][0] }), .spm_out({\spm_out[MCMD][1] , \spm_out[MCMD][0] , 
        \spm_out[MADDR][31] , \spm_out[MADDR][30] , \spm_out[MADDR][29] , 
        \spm_out[MADDR][28] , \spm_out[MADDR][27] , \spm_out[MADDR][26] , 
        \spm_out[MADDR][25] , \spm_out[MADDR][24] , \spm_out[MADDR][23] , 
        \spm_out[MADDR][22] , \spm_out[MADDR][21] , \spm_out[MADDR][20] , 
        \spm_out[MADDR][19] , \spm_out[MADDR][18] , \spm_out[MADDR][17] , 
        \spm_out[MADDR][16] , \spm_out[MADDR][15] , \spm_out[MADDR][14] , 
        \spm_out[MADDR][13] , \spm_out[MADDR][12] , \spm_out[MADDR][11] , 
        \spm_out[MADDR][10] , \spm_out[MADDR][9] , \spm_out[MADDR][8] , 
        \spm_out[MADDR][7] , \spm_out[MADDR][6] , \spm_out[MADDR][5] , 
        \spm_out[MADDR][4] , \spm_out[MADDR][3] , \spm_out[MADDR][2] , 
        \spm_out[MADDR][1] , \spm_out[MADDR][0] , \spm_out[MDATA][63] , 
        \spm_out[MDATA][62] , \spm_out[MDATA][61] , \spm_out[MDATA][60] , 
        \spm_out[MDATA][59] , \spm_out[MDATA][58] , \spm_out[MDATA][57] , 
        \spm_out[MDATA][56] , \spm_out[MDATA][55] , \spm_out[MDATA][54] , 
        \spm_out[MDATA][53] , \spm_out[MDATA][52] , \spm_out[MDATA][51] , 
        \spm_out[MDATA][50] , \spm_out[MDATA][49] , \spm_out[MDATA][48] , 
        \spm_out[MDATA][47] , \spm_out[MDATA][46] , \spm_out[MDATA][45] , 
        \spm_out[MDATA][44] , \spm_out[MDATA][43] , \spm_out[MDATA][42] , 
        \spm_out[MDATA][41] , \spm_out[MDATA][40] , \spm_out[MDATA][39] , 
        \spm_out[MDATA][38] , \spm_out[MDATA][37] , \spm_out[MDATA][36] , 
        \spm_out[MDATA][35] , \spm_out[MDATA][34] , \spm_out[MDATA][33] , 
        \spm_out[MDATA][32] , \spm_out[MDATA][31] , \spm_out[MDATA][30] , 
        \spm_out[MDATA][29] , \spm_out[MDATA][28] , \spm_out[MDATA][27] , 
        \spm_out[MDATA][26] , \spm_out[MDATA][25] , \spm_out[MDATA][24] , 
        \spm_out[MDATA][23] , \spm_out[MDATA][22] , \spm_out[MDATA][21] , 
        \spm_out[MDATA][20] , \spm_out[MDATA][19] , \spm_out[MDATA][18] , 
        \spm_out[MDATA][17] , \spm_out[MDATA][16] , \spm_out[MDATA][15] , 
        \spm_out[MDATA][14] , \spm_out[MDATA][13] , \spm_out[MDATA][12] , 
        \spm_out[MDATA][11] , \spm_out[MDATA][10] , \spm_out[MDATA][9] , 
        \spm_out[MDATA][8] , \spm_out[MDATA][7] , \spm_out[MDATA][6] , 
        \spm_out[MDATA][5] , \spm_out[MDATA][4] , \spm_out[MDATA][3] , 
        \spm_out[MDATA][2] , \spm_out[MDATA][1] , \spm_out[MDATA][0] }), 
    .north_in_f({\north_in_f[REQ] , \north_in_f[DATA][34] , 
        \north_in_f[DATA][33] , \north_in_f[DATA][32] , \north_in_f[DATA][31] , 
        \north_in_f[DATA][30] , \north_in_f[DATA][29] , \north_in_f[DATA][28] , 
        \north_in_f[DATA][27] , \north_in_f[DATA][26] , \north_in_f[DATA][25] , 
        \north_in_f[DATA][24] , \north_in_f[DATA][23] , \north_in_f[DATA][22] , 
        \north_in_f[DATA][21] , \north_in_f[DATA][20] , \north_in_f[DATA][19] , 
        \north_in_f[DATA][18] , \north_in_f[DATA][17] , \north_in_f[DATA][16] , 
        \north_in_f[DATA][15] , \north_in_f[DATA][14] , \north_in_f[DATA][13] , 
        \north_in_f[DATA][12] , \north_in_f[DATA][11] , \north_in_f[DATA][10] , 
        \north_in_f[DATA][9] , \north_in_f[DATA][8] , \north_in_f[DATA][7] , 
        \north_in_f[DATA][6] , \north_in_f[DATA][5] , \north_in_f[DATA][4] , 
        \north_in_f[DATA][3] , \north_in_f[DATA][2] , \north_in_f[DATA][1] , 
        \north_in_f[DATA][0] }), .north_in_b(\north_in_b[ACK] ), .east_in_f({
        \east_in_f[REQ] , \east_in_f[DATA][34] , \east_in_f[DATA][33] , 
        \east_in_f[DATA][32] , \east_in_f[DATA][31] , \east_in_f[DATA][30] , 
        \east_in_f[DATA][29] , \east_in_f[DATA][28] , \east_in_f[DATA][27] , 
        \east_in_f[DATA][26] , \east_in_f[DATA][25] , \east_in_f[DATA][24] , 
        \east_in_f[DATA][23] , \east_in_f[DATA][22] , \east_in_f[DATA][21] , 
        \east_in_f[DATA][20] , \east_in_f[DATA][19] , \east_in_f[DATA][18] , 
        \east_in_f[DATA][17] , \east_in_f[DATA][16] , \east_in_f[DATA][15] , 
        \east_in_f[DATA][14] , \east_in_f[DATA][13] , \east_in_f[DATA][12] , 
        \east_in_f[DATA][11] , \east_in_f[DATA][10] , \east_in_f[DATA][9] , 
        \east_in_f[DATA][8] , \east_in_f[DATA][7] , \east_in_f[DATA][6] , 
        \east_in_f[DATA][5] , \east_in_f[DATA][4] , \east_in_f[DATA][3] , 
        \east_in_f[DATA][2] , \east_in_f[DATA][1] , \east_in_f[DATA][0] }), 
    .east_in_b(\east_in_b[ACK] ), .south_in_f({\south_in_f[REQ] , 
        \south_in_f[DATA][34] , \south_in_f[DATA][33] , \south_in_f[DATA][32] , 
        \south_in_f[DATA][31] , \south_in_f[DATA][30] , \south_in_f[DATA][29] , 
        \south_in_f[DATA][28] , \south_in_f[DATA][27] , \south_in_f[DATA][26] , 
        \south_in_f[DATA][25] , \south_in_f[DATA][24] , \south_in_f[DATA][23] , 
        \south_in_f[DATA][22] , \south_in_f[DATA][21] , \south_in_f[DATA][20] , 
        \south_in_f[DATA][19] , \south_in_f[DATA][18] , \south_in_f[DATA][17] , 
        \south_in_f[DATA][16] , \south_in_f[DATA][15] , \south_in_f[DATA][14] , 
        \south_in_f[DATA][13] , \south_in_f[DATA][12] , \south_in_f[DATA][11] , 
        \south_in_f[DATA][10] , \south_in_f[DATA][9] , \south_in_f[DATA][8] , 
        \south_in_f[DATA][7] , \south_in_f[DATA][6] , \south_in_f[DATA][5] , 
        \south_in_f[DATA][4] , \south_in_f[DATA][3] , \south_in_f[DATA][2] , 
        \south_in_f[DATA][1] , \south_in_f[DATA][0] }), .south_in_b(
        \south_in_b[ACK] ), .west_in_f({\west_in_f[REQ] , 
        \west_in_f[DATA][34] , \west_in_f[DATA][33] , \west_in_f[DATA][32] , 
        \west_in_f[DATA][31] , \west_in_f[DATA][30] , \west_in_f[DATA][29] , 
        \west_in_f[DATA][28] , \west_in_f[DATA][27] , \west_in_f[DATA][26] , 
        \west_in_f[DATA][25] , \west_in_f[DATA][24] , \west_in_f[DATA][23] , 
        \west_in_f[DATA][22] , \west_in_f[DATA][21] , \west_in_f[DATA][20] , 
        \west_in_f[DATA][19] , \west_in_f[DATA][18] , \west_in_f[DATA][17] , 
        \west_in_f[DATA][16] , \west_in_f[DATA][15] , \west_in_f[DATA][14] , 
        \west_in_f[DATA][13] , \west_in_f[DATA][12] , \west_in_f[DATA][11] , 
        \west_in_f[DATA][10] , \west_in_f[DATA][9] , \west_in_f[DATA][8] , 
        \west_in_f[DATA][7] , \west_in_f[DATA][6] , \west_in_f[DATA][5] , 
        \west_in_f[DATA][4] , \west_in_f[DATA][3] , \west_in_f[DATA][2] , 
        \west_in_f[DATA][1] , \west_in_f[DATA][0] }), .west_in_b(
        \west_in_b[ACK] ), .north_out_f({\north_out_f[REQ] , 
        \north_out_f[DATA][34] , \north_out_f[DATA][33] , 
        \north_out_f[DATA][32] , \north_out_f[DATA][31] , 
        \north_out_f[DATA][30] , \north_out_f[DATA][29] , 
        \north_out_f[DATA][28] , \north_out_f[DATA][27] , 
        \north_out_f[DATA][26] , \north_out_f[DATA][25] , 
        \north_out_f[DATA][24] , \north_out_f[DATA][23] , 
        \north_out_f[DATA][22] , \north_out_f[DATA][21] , 
        \north_out_f[DATA][20] , \north_out_f[DATA][19] , 
        \north_out_f[DATA][18] , \north_out_f[DATA][17] , 
        \north_out_f[DATA][16] , \north_out_f[DATA][15] , 
        \north_out_f[DATA][14] , \north_out_f[DATA][13] , 
        \north_out_f[DATA][12] , \north_out_f[DATA][11] , 
        \north_out_f[DATA][10] , \north_out_f[DATA][9] , 
        \north_out_f[DATA][8] , \north_out_f[DATA][7] , \north_out_f[DATA][6] , 
        \north_out_f[DATA][5] , \north_out_f[DATA][4] , \north_out_f[DATA][3] , 
        \north_out_f[DATA][2] , \north_out_f[DATA][1] , \north_out_f[DATA][0] 
        }), .north_out_b(\north_out_b[ACK] ), .east_out_f({\east_out_f[REQ] , 
        \east_out_f[DATA][34] , \east_out_f[DATA][33] , \east_out_f[DATA][32] , 
        \east_out_f[DATA][31] , \east_out_f[DATA][30] , \east_out_f[DATA][29] , 
        \east_out_f[DATA][28] , \east_out_f[DATA][27] , \east_out_f[DATA][26] , 
        \east_out_f[DATA][25] , \east_out_f[DATA][24] , \east_out_f[DATA][23] , 
        \east_out_f[DATA][22] , \east_out_f[DATA][21] , \east_out_f[DATA][20] , 
        \east_out_f[DATA][19] , \east_out_f[DATA][18] , \east_out_f[DATA][17] , 
        \east_out_f[DATA][16] , \east_out_f[DATA][15] , \east_out_f[DATA][14] , 
        \east_out_f[DATA][13] , \east_out_f[DATA][12] , \east_out_f[DATA][11] , 
        \east_out_f[DATA][10] , \east_out_f[DATA][9] , \east_out_f[DATA][8] , 
        \east_out_f[DATA][7] , \east_out_f[DATA][6] , \east_out_f[DATA][5] , 
        \east_out_f[DATA][4] , \east_out_f[DATA][3] , \east_out_f[DATA][2] , 
        \east_out_f[DATA][1] , \east_out_f[DATA][0] }), .east_out_b(
        \east_out_b[ACK] ), .south_out_f({\south_out_f[REQ] , 
        \south_out_f[DATA][34] , \south_out_f[DATA][33] , 
        \south_out_f[DATA][32] , \south_out_f[DATA][31] , 
        \south_out_f[DATA][30] , \south_out_f[DATA][29] , 
        \south_out_f[DATA][28] , \south_out_f[DATA][27] , 
        \south_out_f[DATA][26] , \south_out_f[DATA][25] , 
        \south_out_f[DATA][24] , \south_out_f[DATA][23] , 
        \south_out_f[DATA][22] , \south_out_f[DATA][21] , 
        \south_out_f[DATA][20] , \south_out_f[DATA][19] , 
        \south_out_f[DATA][18] , \south_out_f[DATA][17] , 
        \south_out_f[DATA][16] , \south_out_f[DATA][15] , 
        \south_out_f[DATA][14] , \south_out_f[DATA][13] , 
        \south_out_f[DATA][12] , \south_out_f[DATA][11] , 
        \south_out_f[DATA][10] , \south_out_f[DATA][9] , 
        \south_out_f[DATA][8] , \south_out_f[DATA][7] , \south_out_f[DATA][6] , 
        \south_out_f[DATA][5] , \south_out_f[DATA][4] , \south_out_f[DATA][3] , 
        \south_out_f[DATA][2] , \south_out_f[DATA][1] , \south_out_f[DATA][0] 
        }), .south_out_b(\south_out_b[ACK] ), .west_out_f({\west_out_f[REQ] , 
        \west_out_f[DATA][34] , \west_out_f[DATA][33] , \west_out_f[DATA][32] , 
        \west_out_f[DATA][31] , \west_out_f[DATA][30] , \west_out_f[DATA][29] , 
        \west_out_f[DATA][28] , \west_out_f[DATA][27] , \west_out_f[DATA][26] , 
        \west_out_f[DATA][25] , \west_out_f[DATA][24] , \west_out_f[DATA][23] , 
        \west_out_f[DATA][22] , \west_out_f[DATA][21] , \west_out_f[DATA][20] , 
        \west_out_f[DATA][19] , \west_out_f[DATA][18] , \west_out_f[DATA][17] , 
        \west_out_f[DATA][16] , \west_out_f[DATA][15] , \west_out_f[DATA][14] , 
        \west_out_f[DATA][13] , \west_out_f[DATA][12] , \west_out_f[DATA][11] , 
        \west_out_f[DATA][10] , \west_out_f[DATA][9] , \west_out_f[DATA][8] , 
        \west_out_f[DATA][7] , \west_out_f[DATA][6] , \west_out_f[DATA][5] , 
        \west_out_f[DATA][4] , \west_out_f[DATA][3] , \west_out_f[DATA][2] , 
        \west_out_f[DATA][1] , \west_out_f[DATA][0] }), .west_out_b(
        \west_out_b[ACK] ) );
  input p_clk, n_clk, reset, \proc_in[MCMD][1] , \proc_in[MCMD][0] ,
         \proc_in[MADDR][31] , \proc_in[MADDR][30] , \proc_in[MADDR][29] ,
         \proc_in[MADDR][28] , \proc_in[MADDR][27] , \proc_in[MADDR][26] ,
         \proc_in[MADDR][25] , \proc_in[MADDR][24] , \proc_in[MADDR][23] ,
         \proc_in[MADDR][22] , \proc_in[MADDR][21] , \proc_in[MADDR][20] ,
         \proc_in[MADDR][19] , \proc_in[MADDR][18] , \proc_in[MADDR][17] ,
         \proc_in[MADDR][16] , \proc_in[MADDR][15] , \proc_in[MADDR][14] ,
         \proc_in[MADDR][13] , \proc_in[MADDR][12] , \proc_in[MADDR][11] ,
         \proc_in[MADDR][10] , \proc_in[MADDR][9] , \proc_in[MADDR][8] ,
         \proc_in[MADDR][7] , \proc_in[MADDR][6] , \proc_in[MADDR][5] ,
         \proc_in[MADDR][4] , \proc_in[MADDR][3] , \proc_in[MADDR][2] ,
         \proc_in[MADDR][1] , \proc_in[MADDR][0] , \proc_in[MDATA][31] ,
         \proc_in[MDATA][30] , \proc_in[MDATA][29] , \proc_in[MDATA][28] ,
         \proc_in[MDATA][27] , \proc_in[MDATA][26] , \proc_in[MDATA][25] ,
         \proc_in[MDATA][24] , \proc_in[MDATA][23] , \proc_in[MDATA][22] ,
         \proc_in[MDATA][21] , \proc_in[MDATA][20] , \proc_in[MDATA][19] ,
         \proc_in[MDATA][18] , \proc_in[MDATA][17] , \proc_in[MDATA][16] ,
         \proc_in[MDATA][15] , \proc_in[MDATA][14] , \proc_in[MDATA][13] ,
         \proc_in[MDATA][12] , \proc_in[MDATA][11] , \proc_in[MDATA][10] ,
         \proc_in[MDATA][9] , \proc_in[MDATA][8] , \proc_in[MDATA][7] ,
         \proc_in[MDATA][6] , \proc_in[MDATA][5] , \proc_in[MDATA][4] ,
         \proc_in[MDATA][3] , \proc_in[MDATA][2] , \proc_in[MDATA][1] ,
         \proc_in[MDATA][0] , \spm_in[SCMDACCEPT] , \spm_in[SRESP] ,
         \spm_in[SDATA][63] , \spm_in[SDATA][62] , \spm_in[SDATA][61] ,
         \spm_in[SDATA][60] , \spm_in[SDATA][59] , \spm_in[SDATA][58] ,
         \spm_in[SDATA][57] , \spm_in[SDATA][56] , \spm_in[SDATA][55] ,
         \spm_in[SDATA][54] , \spm_in[SDATA][53] , \spm_in[SDATA][52] ,
         \spm_in[SDATA][51] , \spm_in[SDATA][50] , \spm_in[SDATA][49] ,
         \spm_in[SDATA][48] , \spm_in[SDATA][47] , \spm_in[SDATA][46] ,
         \spm_in[SDATA][45] , \spm_in[SDATA][44] , \spm_in[SDATA][43] ,
         \spm_in[SDATA][42] , \spm_in[SDATA][41] , \spm_in[SDATA][40] ,
         \spm_in[SDATA][39] , \spm_in[SDATA][38] , \spm_in[SDATA][37] ,
         \spm_in[SDATA][36] , \spm_in[SDATA][35] , \spm_in[SDATA][34] ,
         \spm_in[SDATA][33] , \spm_in[SDATA][32] , \spm_in[SDATA][31] ,
         \spm_in[SDATA][30] , \spm_in[SDATA][29] , \spm_in[SDATA][28] ,
         \spm_in[SDATA][27] , \spm_in[SDATA][26] , \spm_in[SDATA][25] ,
         \spm_in[SDATA][24] , \spm_in[SDATA][23] , \spm_in[SDATA][22] ,
         \spm_in[SDATA][21] , \spm_in[SDATA][20] , \spm_in[SDATA][19] ,
         \spm_in[SDATA][18] , \spm_in[SDATA][17] , \spm_in[SDATA][16] ,
         \spm_in[SDATA][15] , \spm_in[SDATA][14] , \spm_in[SDATA][13] ,
         \spm_in[SDATA][12] , \spm_in[SDATA][11] , \spm_in[SDATA][10] ,
         \spm_in[SDATA][9] , \spm_in[SDATA][8] , \spm_in[SDATA][7] ,
         \spm_in[SDATA][6] , \spm_in[SDATA][5] , \spm_in[SDATA][4] ,
         \spm_in[SDATA][3] , \spm_in[SDATA][2] , \spm_in[SDATA][1] ,
         \spm_in[SDATA][0] , \north_in_f[REQ] , \north_in_f[DATA][34] ,
         \north_in_f[DATA][33] , \north_in_f[DATA][32] ,
         \north_in_f[DATA][31] , \north_in_f[DATA][30] ,
         \north_in_f[DATA][29] , \north_in_f[DATA][28] ,
         \north_in_f[DATA][27] , \north_in_f[DATA][26] ,
         \north_in_f[DATA][25] , \north_in_f[DATA][24] ,
         \north_in_f[DATA][23] , \north_in_f[DATA][22] ,
         \north_in_f[DATA][21] , \north_in_f[DATA][20] ,
         \north_in_f[DATA][19] , \north_in_f[DATA][18] ,
         \north_in_f[DATA][17] , \north_in_f[DATA][16] ,
         \north_in_f[DATA][15] , \north_in_f[DATA][14] ,
         \north_in_f[DATA][13] , \north_in_f[DATA][12] ,
         \north_in_f[DATA][11] , \north_in_f[DATA][10] , \north_in_f[DATA][9] ,
         \north_in_f[DATA][8] , \north_in_f[DATA][7] , \north_in_f[DATA][6] ,
         \north_in_f[DATA][5] , \north_in_f[DATA][4] , \north_in_f[DATA][3] ,
         \north_in_f[DATA][2] , \north_in_f[DATA][1] , \north_in_f[DATA][0] ,
         \east_in_f[REQ] , \east_in_f[DATA][34] , \east_in_f[DATA][33] ,
         \east_in_f[DATA][32] , \east_in_f[DATA][31] , \east_in_f[DATA][30] ,
         \east_in_f[DATA][29] , \east_in_f[DATA][28] , \east_in_f[DATA][27] ,
         \east_in_f[DATA][26] , \east_in_f[DATA][25] , \east_in_f[DATA][24] ,
         \east_in_f[DATA][23] , \east_in_f[DATA][22] , \east_in_f[DATA][21] ,
         \east_in_f[DATA][20] , \east_in_f[DATA][19] , \east_in_f[DATA][18] ,
         \east_in_f[DATA][17] , \east_in_f[DATA][16] , \east_in_f[DATA][15] ,
         \east_in_f[DATA][14] , \east_in_f[DATA][13] , \east_in_f[DATA][12] ,
         \east_in_f[DATA][11] , \east_in_f[DATA][10] , \east_in_f[DATA][9] ,
         \east_in_f[DATA][8] , \east_in_f[DATA][7] , \east_in_f[DATA][6] ,
         \east_in_f[DATA][5] , \east_in_f[DATA][4] , \east_in_f[DATA][3] ,
         \east_in_f[DATA][2] , \east_in_f[DATA][1] , \east_in_f[DATA][0] ,
         \south_in_f[REQ] , \south_in_f[DATA][34] , \south_in_f[DATA][33] ,
         \south_in_f[DATA][32] , \south_in_f[DATA][31] ,
         \south_in_f[DATA][30] , \south_in_f[DATA][29] ,
         \south_in_f[DATA][28] , \south_in_f[DATA][27] ,
         \south_in_f[DATA][26] , \south_in_f[DATA][25] ,
         \south_in_f[DATA][24] , \south_in_f[DATA][23] ,
         \south_in_f[DATA][22] , \south_in_f[DATA][21] ,
         \south_in_f[DATA][20] , \south_in_f[DATA][19] ,
         \south_in_f[DATA][18] , \south_in_f[DATA][17] ,
         \south_in_f[DATA][16] , \south_in_f[DATA][15] ,
         \south_in_f[DATA][14] , \south_in_f[DATA][13] ,
         \south_in_f[DATA][12] , \south_in_f[DATA][11] ,
         \south_in_f[DATA][10] , \south_in_f[DATA][9] , \south_in_f[DATA][8] ,
         \south_in_f[DATA][7] , \south_in_f[DATA][6] , \south_in_f[DATA][5] ,
         \south_in_f[DATA][4] , \south_in_f[DATA][3] , \south_in_f[DATA][2] ,
         \south_in_f[DATA][1] , \south_in_f[DATA][0] , \west_in_f[REQ] ,
         \west_in_f[DATA][34] , \west_in_f[DATA][33] , \west_in_f[DATA][32] ,
         \west_in_f[DATA][31] , \west_in_f[DATA][30] , \west_in_f[DATA][29] ,
         \west_in_f[DATA][28] , \west_in_f[DATA][27] , \west_in_f[DATA][26] ,
         \west_in_f[DATA][25] , \west_in_f[DATA][24] , \west_in_f[DATA][23] ,
         \west_in_f[DATA][22] , \west_in_f[DATA][21] , \west_in_f[DATA][20] ,
         \west_in_f[DATA][19] , \west_in_f[DATA][18] , \west_in_f[DATA][17] ,
         \west_in_f[DATA][16] , \west_in_f[DATA][15] , \west_in_f[DATA][14] ,
         \west_in_f[DATA][13] , \west_in_f[DATA][12] , \west_in_f[DATA][11] ,
         \west_in_f[DATA][10] , \west_in_f[DATA][9] , \west_in_f[DATA][8] ,
         \west_in_f[DATA][7] , \west_in_f[DATA][6] , \west_in_f[DATA][5] ,
         \west_in_f[DATA][4] , \west_in_f[DATA][3] , \west_in_f[DATA][2] ,
         \west_in_f[DATA][1] , \west_in_f[DATA][0] , \north_out_b[ACK] ,
         \east_out_b[ACK] , \south_out_b[ACK] , \west_out_b[ACK] ;
  output \proc_out[SCMDACCEPT] , \proc_out[SRESP] , \proc_out[SDATA][31] ,
         \proc_out[SDATA][30] , \proc_out[SDATA][29] , \proc_out[SDATA][28] ,
         \proc_out[SDATA][27] , \proc_out[SDATA][26] , \proc_out[SDATA][25] ,
         \proc_out[SDATA][24] , \proc_out[SDATA][23] , \proc_out[SDATA][22] ,
         \proc_out[SDATA][21] , \proc_out[SDATA][20] , \proc_out[SDATA][19] ,
         \proc_out[SDATA][18] , \proc_out[SDATA][17] , \proc_out[SDATA][16] ,
         \proc_out[SDATA][15] , \proc_out[SDATA][14] , \proc_out[SDATA][13] ,
         \proc_out[SDATA][12] , \proc_out[SDATA][11] , \proc_out[SDATA][10] ,
         \proc_out[SDATA][9] , \proc_out[SDATA][8] , \proc_out[SDATA][7] ,
         \proc_out[SDATA][6] , \proc_out[SDATA][5] , \proc_out[SDATA][4] ,
         \proc_out[SDATA][3] , \proc_out[SDATA][2] , \proc_out[SDATA][1] ,
         \proc_out[SDATA][0] , \spm_out[MCMD][1] , \spm_out[MCMD][0] ,
         \spm_out[MADDR][31] , \spm_out[MADDR][30] , \spm_out[MADDR][29] ,
         \spm_out[MADDR][28] , \spm_out[MADDR][27] , \spm_out[MADDR][26] ,
         \spm_out[MADDR][25] , \spm_out[MADDR][24] , \spm_out[MADDR][23] ,
         \spm_out[MADDR][22] , \spm_out[MADDR][21] , \spm_out[MADDR][20] ,
         \spm_out[MADDR][19] , \spm_out[MADDR][18] , \spm_out[MADDR][17] ,
         \spm_out[MADDR][16] , \spm_out[MADDR][15] , \spm_out[MADDR][14] ,
         \spm_out[MADDR][13] , \spm_out[MADDR][12] , \spm_out[MADDR][11] ,
         \spm_out[MADDR][10] , \spm_out[MADDR][9] , \spm_out[MADDR][8] ,
         \spm_out[MADDR][7] , \spm_out[MADDR][6] , \spm_out[MADDR][5] ,
         \spm_out[MADDR][4] , \spm_out[MADDR][3] , \spm_out[MADDR][2] ,
         \spm_out[MADDR][1] , \spm_out[MADDR][0] , \spm_out[MDATA][63] ,
         \spm_out[MDATA][62] , \spm_out[MDATA][61] , \spm_out[MDATA][60] ,
         \spm_out[MDATA][59] , \spm_out[MDATA][58] , \spm_out[MDATA][57] ,
         \spm_out[MDATA][56] , \spm_out[MDATA][55] , \spm_out[MDATA][54] ,
         \spm_out[MDATA][53] , \spm_out[MDATA][52] , \spm_out[MDATA][51] ,
         \spm_out[MDATA][50] , \spm_out[MDATA][49] , \spm_out[MDATA][48] ,
         \spm_out[MDATA][47] , \spm_out[MDATA][46] , \spm_out[MDATA][45] ,
         \spm_out[MDATA][44] , \spm_out[MDATA][43] , \spm_out[MDATA][42] ,
         \spm_out[MDATA][41] , \spm_out[MDATA][40] , \spm_out[MDATA][39] ,
         \spm_out[MDATA][38] , \spm_out[MDATA][37] , \spm_out[MDATA][36] ,
         \spm_out[MDATA][35] , \spm_out[MDATA][34] , \spm_out[MDATA][33] ,
         \spm_out[MDATA][32] , \spm_out[MDATA][31] , \spm_out[MDATA][30] ,
         \spm_out[MDATA][29] , \spm_out[MDATA][28] , \spm_out[MDATA][27] ,
         \spm_out[MDATA][26] , \spm_out[MDATA][25] , \spm_out[MDATA][24] ,
         \spm_out[MDATA][23] , \spm_out[MDATA][22] , \spm_out[MDATA][21] ,
         \spm_out[MDATA][20] , \spm_out[MDATA][19] , \spm_out[MDATA][18] ,
         \spm_out[MDATA][17] , \spm_out[MDATA][16] , \spm_out[MDATA][15] ,
         \spm_out[MDATA][14] , \spm_out[MDATA][13] , \spm_out[MDATA][12] ,
         \spm_out[MDATA][11] , \spm_out[MDATA][10] , \spm_out[MDATA][9] ,
         \spm_out[MDATA][8] , \spm_out[MDATA][7] , \spm_out[MDATA][6] ,
         \spm_out[MDATA][5] , \spm_out[MDATA][4] , \spm_out[MDATA][3] ,
         \spm_out[MDATA][2] , \spm_out[MDATA][1] , \spm_out[MDATA][0] ,
         \north_in_b[ACK] , \east_in_b[ACK] , \south_in_b[ACK] ,
         \west_in_b[ACK] , \north_out_f[REQ] , \north_out_f[DATA][34] ,
         \north_out_f[DATA][33] , \north_out_f[DATA][32] ,
         \north_out_f[DATA][31] , \north_out_f[DATA][30] ,
         \north_out_f[DATA][29] , \north_out_f[DATA][28] ,
         \north_out_f[DATA][27] , \north_out_f[DATA][26] ,
         \north_out_f[DATA][25] , \north_out_f[DATA][24] ,
         \north_out_f[DATA][23] , \north_out_f[DATA][22] ,
         \north_out_f[DATA][21] , \north_out_f[DATA][20] ,
         \north_out_f[DATA][19] , \north_out_f[DATA][18] ,
         \north_out_f[DATA][17] , \north_out_f[DATA][16] ,
         \north_out_f[DATA][15] , \north_out_f[DATA][14] ,
         \north_out_f[DATA][13] , \north_out_f[DATA][12] ,
         \north_out_f[DATA][11] , \north_out_f[DATA][10] ,
         \north_out_f[DATA][9] , \north_out_f[DATA][8] ,
         \north_out_f[DATA][7] , \north_out_f[DATA][6] ,
         \north_out_f[DATA][5] , \north_out_f[DATA][4] ,
         \north_out_f[DATA][3] , \north_out_f[DATA][2] ,
         \north_out_f[DATA][1] , \north_out_f[DATA][0] , \east_out_f[REQ] ,
         \east_out_f[DATA][34] , \east_out_f[DATA][33] ,
         \east_out_f[DATA][32] , \east_out_f[DATA][31] ,
         \east_out_f[DATA][30] , \east_out_f[DATA][29] ,
         \east_out_f[DATA][28] , \east_out_f[DATA][27] ,
         \east_out_f[DATA][26] , \east_out_f[DATA][25] ,
         \east_out_f[DATA][24] , \east_out_f[DATA][23] ,
         \east_out_f[DATA][22] , \east_out_f[DATA][21] ,
         \east_out_f[DATA][20] , \east_out_f[DATA][19] ,
         \east_out_f[DATA][18] , \east_out_f[DATA][17] ,
         \east_out_f[DATA][16] , \east_out_f[DATA][15] ,
         \east_out_f[DATA][14] , \east_out_f[DATA][13] ,
         \east_out_f[DATA][12] , \east_out_f[DATA][11] ,
         \east_out_f[DATA][10] , \east_out_f[DATA][9] , \east_out_f[DATA][8] ,
         \east_out_f[DATA][7] , \east_out_f[DATA][6] , \east_out_f[DATA][5] ,
         \east_out_f[DATA][4] , \east_out_f[DATA][3] , \east_out_f[DATA][2] ,
         \east_out_f[DATA][1] , \east_out_f[DATA][0] , \south_out_f[REQ] ,
         \south_out_f[DATA][34] , \south_out_f[DATA][33] ,
         \south_out_f[DATA][32] , \south_out_f[DATA][31] ,
         \south_out_f[DATA][30] , \south_out_f[DATA][29] ,
         \south_out_f[DATA][28] , \south_out_f[DATA][27] ,
         \south_out_f[DATA][26] , \south_out_f[DATA][25] ,
         \south_out_f[DATA][24] , \south_out_f[DATA][23] ,
         \south_out_f[DATA][22] , \south_out_f[DATA][21] ,
         \south_out_f[DATA][20] , \south_out_f[DATA][19] ,
         \south_out_f[DATA][18] , \south_out_f[DATA][17] ,
         \south_out_f[DATA][16] , \south_out_f[DATA][15] ,
         \south_out_f[DATA][14] , \south_out_f[DATA][13] ,
         \south_out_f[DATA][12] , \south_out_f[DATA][11] ,
         \south_out_f[DATA][10] , \south_out_f[DATA][9] ,
         \south_out_f[DATA][8] , \south_out_f[DATA][7] ,
         \south_out_f[DATA][6] , \south_out_f[DATA][5] ,
         \south_out_f[DATA][4] , \south_out_f[DATA][3] ,
         \south_out_f[DATA][2] , \south_out_f[DATA][1] ,
         \south_out_f[DATA][0] , \west_out_f[REQ] , \west_out_f[DATA][34] ,
         \west_out_f[DATA][33] , \west_out_f[DATA][32] ,
         \west_out_f[DATA][31] , \west_out_f[DATA][30] ,
         \west_out_f[DATA][29] , \west_out_f[DATA][28] ,
         \west_out_f[DATA][27] , \west_out_f[DATA][26] ,
         \west_out_f[DATA][25] , \west_out_f[DATA][24] ,
         \west_out_f[DATA][23] , \west_out_f[DATA][22] ,
         \west_out_f[DATA][21] , \west_out_f[DATA][20] ,
         \west_out_f[DATA][19] , \west_out_f[DATA][18] ,
         \west_out_f[DATA][17] , \west_out_f[DATA][16] ,
         \west_out_f[DATA][15] , \west_out_f[DATA][14] ,
         \west_out_f[DATA][13] , \west_out_f[DATA][12] ,
         \west_out_f[DATA][11] , \west_out_f[DATA][10] , \west_out_f[DATA][9] ,
         \west_out_f[DATA][8] , \west_out_f[DATA][7] , \west_out_f[DATA][6] ,
         \west_out_f[DATA][5] , \west_out_f[DATA][4] , \west_out_f[DATA][3] ,
         \west_out_f[DATA][2] , \west_out_f[DATA][1] , \west_out_f[DATA][0] ;
  wire   del_half_clk0, \ip_to_net_f[REQ] , n1, n3, n4, n5, n6, n7, n8, n9,
         n10, n11;
  wire   [34:0] net_to_ip;
  wire   [34:0] ip_to_net;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17;
  assign \spm_out[MADDR][31]  = 1'b0;
  assign \spm_out[MADDR][30]  = 1'b0;
  assign \spm_out[MADDR][29]  = 1'b0;
  assign \spm_out[MADDR][28]  = 1'b0;
  assign \spm_out[MADDR][27]  = 1'b0;
  assign \spm_out[MADDR][26]  = 1'b0;
  assign \spm_out[MADDR][25]  = 1'b0;
  assign \spm_out[MADDR][24]  = 1'b0;
  assign \spm_out[MADDR][23]  = 1'b0;
  assign \spm_out[MADDR][22]  = 1'b0;
  assign \spm_out[MADDR][21]  = 1'b0;
  assign \spm_out[MADDR][20]  = 1'b0;
  assign \spm_out[MADDR][19]  = 1'b0;
  assign \spm_out[MADDR][18]  = 1'b0;
  assign \spm_out[MADDR][17]  = 1'b0;
  assign \spm_out[MADDR][16]  = 1'b0;
  assign \spm_out[MADDR][15]  = 1'b0;

  nAdapter_3 na ( .na_clk(n_clk), .na_reset(reset), .proc_in({
        \proc_in[MCMD][1] , \proc_in[MCMD][0] , \proc_in[MADDR][31] , 
        \proc_in[MADDR][30] , \proc_in[MADDR][29] , \proc_in[MADDR][28] , 
        \proc_in[MADDR][27] , \proc_in[MADDR][26] , \proc_in[MADDR][25] , 
        \proc_in[MADDR][24] , \proc_in[MADDR][23] , \proc_in[MADDR][22] , 
        \proc_in[MADDR][21] , \proc_in[MADDR][20] , \proc_in[MADDR][19] , 
        \proc_in[MADDR][18] , \proc_in[MADDR][17] , \proc_in[MADDR][16] , 
        \proc_in[MADDR][15] , \proc_in[MADDR][14] , \proc_in[MADDR][13] , 
        \proc_in[MADDR][12] , \proc_in[MADDR][11] , \proc_in[MADDR][10] , 
        \proc_in[MADDR][9] , \proc_in[MADDR][8] , \proc_in[MADDR][7] , 
        \proc_in[MADDR][6] , \proc_in[MADDR][5] , \proc_in[MADDR][4] , 
        \proc_in[MADDR][3] , \proc_in[MADDR][2] , \proc_in[MADDR][1] , 
        \proc_in[MADDR][0] , \proc_in[MDATA][31] , \proc_in[MDATA][30] , 
        \proc_in[MDATA][29] , \proc_in[MDATA][28] , \proc_in[MDATA][27] , 
        \proc_in[MDATA][26] , \proc_in[MDATA][25] , \proc_in[MDATA][24] , 
        \proc_in[MDATA][23] , \proc_in[MDATA][22] , \proc_in[MDATA][21] , 
        \proc_in[MDATA][20] , \proc_in[MDATA][19] , \proc_in[MDATA][18] , 
        \proc_in[MDATA][17] , \proc_in[MDATA][16] , \proc_in[MDATA][15] , 
        \proc_in[MDATA][14] , \proc_in[MDATA][13] , \proc_in[MDATA][12] , 
        \proc_in[MDATA][11] , \proc_in[MDATA][10] , \proc_in[MDATA][9] , 
        \proc_in[MDATA][8] , \proc_in[MDATA][7] , \proc_in[MDATA][6] , 
        \proc_in[MDATA][5] , \proc_in[MDATA][4] , \proc_in[MDATA][3] , 
        \proc_in[MDATA][2] , \proc_in[MDATA][1] , \proc_in[MDATA][0] }), 
        .proc_out({\proc_out[SCMDACCEPT] , \proc_out[SRESP] , 
        \proc_out[SDATA][31] , \proc_out[SDATA][30] , \proc_out[SDATA][29] , 
        \proc_out[SDATA][28] , \proc_out[SDATA][27] , \proc_out[SDATA][26] , 
        \proc_out[SDATA][25] , \proc_out[SDATA][24] , \proc_out[SDATA][23] , 
        \proc_out[SDATA][22] , \proc_out[SDATA][21] , \proc_out[SDATA][20] , 
        \proc_out[SDATA][19] , \proc_out[SDATA][18] , \proc_out[SDATA][17] , 
        \proc_out[SDATA][16] , \proc_out[SDATA][15] , \proc_out[SDATA][14] , 
        \proc_out[SDATA][13] , \proc_out[SDATA][12] , \proc_out[SDATA][11] , 
        \proc_out[SDATA][10] , \proc_out[SDATA][9] , \proc_out[SDATA][8] , 
        \proc_out[SDATA][7] , \proc_out[SDATA][6] , \proc_out[SDATA][5] , 
        \proc_out[SDATA][4] , \proc_out[SDATA][3] , \proc_out[SDATA][2] , 
        \proc_out[SDATA][1] , \proc_out[SDATA][0] }), .spm_in({
        \spm_in[SCMDACCEPT] , \spm_in[SRESP] , \spm_in[SDATA][63] , 
        \spm_in[SDATA][62] , \spm_in[SDATA][61] , \spm_in[SDATA][60] , 
        \spm_in[SDATA][59] , \spm_in[SDATA][58] , \spm_in[SDATA][57] , 
        \spm_in[SDATA][56] , \spm_in[SDATA][55] , \spm_in[SDATA][54] , 
        \spm_in[SDATA][53] , \spm_in[SDATA][52] , \spm_in[SDATA][51] , 
        \spm_in[SDATA][50] , \spm_in[SDATA][49] , \spm_in[SDATA][48] , 
        \spm_in[SDATA][47] , \spm_in[SDATA][46] , \spm_in[SDATA][45] , 
        \spm_in[SDATA][44] , \spm_in[SDATA][43] , \spm_in[SDATA][42] , 
        \spm_in[SDATA][41] , \spm_in[SDATA][40] , \spm_in[SDATA][39] , 
        \spm_in[SDATA][38] , \spm_in[SDATA][37] , \spm_in[SDATA][36] , 
        \spm_in[SDATA][35] , \spm_in[SDATA][34] , \spm_in[SDATA][33] , 
        \spm_in[SDATA][32] , \spm_in[SDATA][31] , \spm_in[SDATA][30] , 
        \spm_in[SDATA][29] , \spm_in[SDATA][28] , \spm_in[SDATA][27] , 
        \spm_in[SDATA][26] , \spm_in[SDATA][25] , \spm_in[SDATA][24] , 
        \spm_in[SDATA][23] , \spm_in[SDATA][22] , \spm_in[SDATA][21] , 
        \spm_in[SDATA][20] , \spm_in[SDATA][19] , \spm_in[SDATA][18] , 
        \spm_in[SDATA][17] , \spm_in[SDATA][16] , \spm_in[SDATA][15] , 
        \spm_in[SDATA][14] , \spm_in[SDATA][13] , \spm_in[SDATA][12] , 
        \spm_in[SDATA][11] , \spm_in[SDATA][10] , \spm_in[SDATA][9] , 
        \spm_in[SDATA][8] , \spm_in[SDATA][7] , \spm_in[SDATA][6] , 
        \spm_in[SDATA][5] , \spm_in[SDATA][4] , \spm_in[SDATA][3] , 
        \spm_in[SDATA][2] , \spm_in[SDATA][1] , \spm_in[SDATA][0] }), 
        .spm_out({\spm_out[MCMD][1] , \spm_out[MCMD][0] , 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, \spm_out[MADDR][14] , \spm_out[MADDR][13] , 
        \spm_out[MADDR][12] , \spm_out[MADDR][11] , \spm_out[MADDR][10] , 
        \spm_out[MADDR][9] , \spm_out[MADDR][8] , \spm_out[MADDR][7] , 
        \spm_out[MADDR][6] , \spm_out[MADDR][5] , \spm_out[MADDR][4] , 
        \spm_out[MADDR][3] , \spm_out[MADDR][2] , \spm_out[MADDR][1] , 
        \spm_out[MADDR][0] , \spm_out[MDATA][63] , \spm_out[MDATA][62] , 
        \spm_out[MDATA][61] , \spm_out[MDATA][60] , \spm_out[MDATA][59] , 
        \spm_out[MDATA][58] , \spm_out[MDATA][57] , \spm_out[MDATA][56] , 
        \spm_out[MDATA][55] , \spm_out[MDATA][54] , \spm_out[MDATA][53] , 
        \spm_out[MDATA][52] , \spm_out[MDATA][51] , \spm_out[MDATA][50] , 
        \spm_out[MDATA][49] , \spm_out[MDATA][48] , \spm_out[MDATA][47] , 
        \spm_out[MDATA][46] , \spm_out[MDATA][45] , \spm_out[MDATA][44] , 
        \spm_out[MDATA][43] , \spm_out[MDATA][42] , \spm_out[MDATA][41] , 
        \spm_out[MDATA][40] , \spm_out[MDATA][39] , \spm_out[MDATA][38] , 
        \spm_out[MDATA][37] , \spm_out[MDATA][36] , \spm_out[MDATA][35] , 
        \spm_out[MDATA][34] , \spm_out[MDATA][33] , \spm_out[MDATA][32] , 
        \spm_out[MDATA][31] , \spm_out[MDATA][30] , \spm_out[MDATA][29] , 
        \spm_out[MDATA][28] , \spm_out[MDATA][27] , \spm_out[MDATA][26] , 
        \spm_out[MDATA][25] , \spm_out[MDATA][24] , \spm_out[MDATA][23] , 
        \spm_out[MDATA][22] , \spm_out[MDATA][21] , \spm_out[MDATA][20] , 
        \spm_out[MDATA][19] , \spm_out[MDATA][18] , \spm_out[MDATA][17] , 
        \spm_out[MDATA][16] , \spm_out[MDATA][15] , \spm_out[MDATA][14] , 
        \spm_out[MDATA][13] , \spm_out[MDATA][12] , \spm_out[MDATA][11] , 
        \spm_out[MDATA][10] , \spm_out[MDATA][9] , \spm_out[MDATA][8] , 
        \spm_out[MDATA][7] , \spm_out[MDATA][6] , \spm_out[MDATA][5] , 
        \spm_out[MDATA][4] , \spm_out[MDATA][3] , \spm_out[MDATA][2] , 
        \spm_out[MDATA][1] , \spm_out[MDATA][0] }), .pkt_in(net_to_ip), 
        .pkt_out(ip_to_net) );
  noc_switch_3 r ( .preset(reset), .north_in_f({\north_in_f[REQ] , 
        \north_in_f[DATA][34] , \north_in_f[DATA][33] , \north_in_f[DATA][32] , 
        \north_in_f[DATA][31] , \north_in_f[DATA][30] , \north_in_f[DATA][29] , 
        \north_in_f[DATA][28] , \north_in_f[DATA][27] , \north_in_f[DATA][26] , 
        \north_in_f[DATA][25] , \north_in_f[DATA][24] , \north_in_f[DATA][23] , 
        \north_in_f[DATA][22] , \north_in_f[DATA][21] , \north_in_f[DATA][20] , 
        \north_in_f[DATA][19] , \north_in_f[DATA][18] , \north_in_f[DATA][17] , 
        \north_in_f[DATA][16] , \north_in_f[DATA][15] , \north_in_f[DATA][14] , 
        \north_in_f[DATA][13] , \north_in_f[DATA][12] , \north_in_f[DATA][11] , 
        \north_in_f[DATA][10] , \north_in_f[DATA][9] , \north_in_f[DATA][8] , 
        \north_in_f[DATA][7] , \north_in_f[DATA][6] , \north_in_f[DATA][5] , 
        \north_in_f[DATA][4] , \north_in_f[DATA][3] , \north_in_f[DATA][2] , 
        \north_in_f[DATA][1] , \north_in_f[DATA][0] }), .north_in_b(
        \north_in_b[ACK] ), .east_in_f({\east_in_f[REQ] , 
        \east_in_f[DATA][34] , \east_in_f[DATA][33] , \east_in_f[DATA][32] , 
        \east_in_f[DATA][31] , \east_in_f[DATA][30] , \east_in_f[DATA][29] , 
        \east_in_f[DATA][28] , \east_in_f[DATA][27] , \east_in_f[DATA][26] , 
        \east_in_f[DATA][25] , \east_in_f[DATA][24] , \east_in_f[DATA][23] , 
        \east_in_f[DATA][22] , \east_in_f[DATA][21] , \east_in_f[DATA][20] , 
        \east_in_f[DATA][19] , \east_in_f[DATA][18] , \east_in_f[DATA][17] , 
        \east_in_f[DATA][16] , \east_in_f[DATA][15] , \east_in_f[DATA][14] , 
        \east_in_f[DATA][13] , \east_in_f[DATA][12] , \east_in_f[DATA][11] , 
        \east_in_f[DATA][10] , \east_in_f[DATA][9] , \east_in_f[DATA][8] , 
        \east_in_f[DATA][7] , \east_in_f[DATA][6] , \east_in_f[DATA][5] , 
        \east_in_f[DATA][4] , \east_in_f[DATA][3] , \east_in_f[DATA][2] , 
        \east_in_f[DATA][1] , \east_in_f[DATA][0] }), .east_in_b(
        \east_in_b[ACK] ), .south_in_f({\south_in_f[REQ] , 
        \south_in_f[DATA][34] , \south_in_f[DATA][33] , \south_in_f[DATA][32] , 
        \south_in_f[DATA][31] , \south_in_f[DATA][30] , \south_in_f[DATA][29] , 
        \south_in_f[DATA][28] , \south_in_f[DATA][27] , \south_in_f[DATA][26] , 
        \south_in_f[DATA][25] , \south_in_f[DATA][24] , \south_in_f[DATA][23] , 
        \south_in_f[DATA][22] , \south_in_f[DATA][21] , \south_in_f[DATA][20] , 
        \south_in_f[DATA][19] , \south_in_f[DATA][18] , \south_in_f[DATA][17] , 
        \south_in_f[DATA][16] , \south_in_f[DATA][15] , \south_in_f[DATA][14] , 
        \south_in_f[DATA][13] , \south_in_f[DATA][12] , \south_in_f[DATA][11] , 
        \south_in_f[DATA][10] , \south_in_f[DATA][9] , \south_in_f[DATA][8] , 
        \south_in_f[DATA][7] , \south_in_f[DATA][6] , \south_in_f[DATA][5] , 
        \south_in_f[DATA][4] , \south_in_f[DATA][3] , \south_in_f[DATA][2] , 
        \south_in_f[DATA][1] , \south_in_f[DATA][0] }), .south_in_b(
        \south_in_b[ACK] ), .west_in_f({\west_in_f[REQ] , 
        \west_in_f[DATA][34] , \west_in_f[DATA][33] , \west_in_f[DATA][32] , 
        \west_in_f[DATA][31] , \west_in_f[DATA][30] , \west_in_f[DATA][29] , 
        \west_in_f[DATA][28] , \west_in_f[DATA][27] , \west_in_f[DATA][26] , 
        \west_in_f[DATA][25] , \west_in_f[DATA][24] , \west_in_f[DATA][23] , 
        \west_in_f[DATA][22] , \west_in_f[DATA][21] , \west_in_f[DATA][20] , 
        \west_in_f[DATA][19] , \west_in_f[DATA][18] , \west_in_f[DATA][17] , 
        \west_in_f[DATA][16] , \west_in_f[DATA][15] , \west_in_f[DATA][14] , 
        \west_in_f[DATA][13] , \west_in_f[DATA][12] , \west_in_f[DATA][11] , 
        \west_in_f[DATA][10] , \west_in_f[DATA][9] , \west_in_f[DATA][8] , 
        \west_in_f[DATA][7] , \west_in_f[DATA][6] , \west_in_f[DATA][5] , 
        \west_in_f[DATA][4] , \west_in_f[DATA][3] , \west_in_f[DATA][2] , 
        \west_in_f[DATA][1] , \west_in_f[DATA][0] }), .west_in_b(
        \west_in_b[ACK] ), .resource_in_f({\ip_to_net_f[REQ] , ip_to_net}), 
        .north_out_f({\north_out_f[REQ] , \north_out_f[DATA][34] , 
        \north_out_f[DATA][33] , \north_out_f[DATA][32] , 
        \north_out_f[DATA][31] , \north_out_f[DATA][30] , 
        \north_out_f[DATA][29] , \north_out_f[DATA][28] , 
        \north_out_f[DATA][27] , \north_out_f[DATA][26] , 
        \north_out_f[DATA][25] , \north_out_f[DATA][24] , 
        \north_out_f[DATA][23] , \north_out_f[DATA][22] , 
        \north_out_f[DATA][21] , \north_out_f[DATA][20] , 
        \north_out_f[DATA][19] , \north_out_f[DATA][18] , 
        \north_out_f[DATA][17] , \north_out_f[DATA][16] , 
        \north_out_f[DATA][15] , \north_out_f[DATA][14] , 
        \north_out_f[DATA][13] , \north_out_f[DATA][12] , 
        \north_out_f[DATA][11] , \north_out_f[DATA][10] , 
        \north_out_f[DATA][9] , \north_out_f[DATA][8] , \north_out_f[DATA][7] , 
        \north_out_f[DATA][6] , \north_out_f[DATA][5] , \north_out_f[DATA][4] , 
        \north_out_f[DATA][3] , \north_out_f[DATA][2] , \north_out_f[DATA][1] , 
        \north_out_f[DATA][0] }), .north_out_b(\north_out_b[ACK] ), 
        .east_out_f({\east_out_f[REQ] , \east_out_f[DATA][34] , 
        \east_out_f[DATA][33] , \east_out_f[DATA][32] , \east_out_f[DATA][31] , 
        \east_out_f[DATA][30] , \east_out_f[DATA][29] , \east_out_f[DATA][28] , 
        \east_out_f[DATA][27] , \east_out_f[DATA][26] , \east_out_f[DATA][25] , 
        \east_out_f[DATA][24] , \east_out_f[DATA][23] , \east_out_f[DATA][22] , 
        \east_out_f[DATA][21] , \east_out_f[DATA][20] , \east_out_f[DATA][19] , 
        \east_out_f[DATA][18] , \east_out_f[DATA][17] , \east_out_f[DATA][16] , 
        \east_out_f[DATA][15] , \east_out_f[DATA][14] , \east_out_f[DATA][13] , 
        \east_out_f[DATA][12] , \east_out_f[DATA][11] , \east_out_f[DATA][10] , 
        \east_out_f[DATA][9] , \east_out_f[DATA][8] , \east_out_f[DATA][7] , 
        \east_out_f[DATA][6] , \east_out_f[DATA][5] , \east_out_f[DATA][4] , 
        \east_out_f[DATA][3] , \east_out_f[DATA][2] , \east_out_f[DATA][1] , 
        \east_out_f[DATA][0] }), .east_out_b(\east_out_b[ACK] ), .south_out_f(
        {\south_out_f[REQ] , \south_out_f[DATA][34] , \south_out_f[DATA][33] , 
        \south_out_f[DATA][32] , \south_out_f[DATA][31] , 
        \south_out_f[DATA][30] , \south_out_f[DATA][29] , 
        \south_out_f[DATA][28] , \south_out_f[DATA][27] , 
        \south_out_f[DATA][26] , \south_out_f[DATA][25] , 
        \south_out_f[DATA][24] , \south_out_f[DATA][23] , 
        \south_out_f[DATA][22] , \south_out_f[DATA][21] , 
        \south_out_f[DATA][20] , \south_out_f[DATA][19] , 
        \south_out_f[DATA][18] , \south_out_f[DATA][17] , 
        \south_out_f[DATA][16] , \south_out_f[DATA][15] , 
        \south_out_f[DATA][14] , \south_out_f[DATA][13] , 
        \south_out_f[DATA][12] , \south_out_f[DATA][11] , 
        \south_out_f[DATA][10] , \south_out_f[DATA][9] , 
        \south_out_f[DATA][8] , \south_out_f[DATA][7] , \south_out_f[DATA][6] , 
        \south_out_f[DATA][5] , \south_out_f[DATA][4] , \south_out_f[DATA][3] , 
        \south_out_f[DATA][2] , \south_out_f[DATA][1] , \south_out_f[DATA][0] }), .south_out_b(\south_out_b[ACK] ), .west_out_f({\west_out_f[REQ] , 
        \west_out_f[DATA][34] , \west_out_f[DATA][33] , \west_out_f[DATA][32] , 
        \west_out_f[DATA][31] , \west_out_f[DATA][30] , \west_out_f[DATA][29] , 
        \west_out_f[DATA][28] , \west_out_f[DATA][27] , \west_out_f[DATA][26] , 
        \west_out_f[DATA][25] , \west_out_f[DATA][24] , \west_out_f[DATA][23] , 
        \west_out_f[DATA][22] , \west_out_f[DATA][21] , \west_out_f[DATA][20] , 
        \west_out_f[DATA][19] , \west_out_f[DATA][18] , \west_out_f[DATA][17] , 
        \west_out_f[DATA][16] , \west_out_f[DATA][15] , \west_out_f[DATA][14] , 
        \west_out_f[DATA][13] , \west_out_f[DATA][12] , \west_out_f[DATA][11] , 
        \west_out_f[DATA][10] , \west_out_f[DATA][9] , \west_out_f[DATA][8] , 
        \west_out_f[DATA][7] , \west_out_f[DATA][6] , \west_out_f[DATA][5] , 
        \west_out_f[DATA][4] , \west_out_f[DATA][3] , \west_out_f[DATA][2] , 
        \west_out_f[DATA][1] , \west_out_f[DATA][0] }), .west_out_b(
        \west_out_b[ACK] ), .resource_out_f({SYNOPSYS_UNCONNECTED__17, 
        net_to_ip}), .resource_out_b(n9) );
  HS65_LS_DFPRQNX9 half_clk_reg ( .D(n11), .CP(n_clk), .RN(n8), .QN(n11) );
  HS65_LS_IVX9 I_2 ( .A(n4), .Z(\ip_to_net_f[REQ] ) );
  HS65_LH_IVX2 I_1 ( .A(n10), .Z(del_half_clk0) );
  HS65_LS_IVX9 U3 ( .A(n11), .Z(n10) );
  HS65_LH_IVX2 U4 ( .A(n1), .Z(n3) );
  HS65_LS_IVX106 U5 ( .A(del_half_clk0), .Z(n1) );
  HS65_LS_BFX9 U6 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U7 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U8 ( .A(n7), .Z(n6) );
  HS65_LS_BFX9 U9 ( .A(n3), .Z(n7) );
  HS65_LS_IVX9 U10 ( .A(reset), .Z(n8) );
  HS65_LS_IVX9 U11 ( .A(del_half_clk0), .Z(n9) );
endmodule


module counter_WIDTH3_2 ( clk, reset, enable, cnt );
  output [2:0] cnt;
  input clk, reset, enable;
  wire   n1, n2, n3, n4, n5, n8, n9, n10, n11;

  HS65_LS_DFPRQX9 \reg_reg[0]  ( .D(n5), .CP(clk), .RN(n1), .Q(cnt[0]) );
  HS65_LS_DFPRQX9 \reg_reg[2]  ( .D(n8), .CP(clk), .RN(n1), .Q(cnt[2]) );
  HS65_LS_DFPRQX9 \reg_reg[1]  ( .D(n9), .CP(clk), .RN(n1), .Q(cnt[1]) );
  HS65_LS_IVX9 U3 ( .A(reset), .Z(n1) );
  HS65_LS_OAI32X5 U4 ( .A(n4), .B(n11), .C(n2), .D(enable), .E(n3), .Z(n8) );
  HS65_LS_NAND2X7 U5 ( .A(enable), .B(n3), .Z(n11) );
  HS65_LS_OAI32X5 U6 ( .A(n2), .B(cnt[1]), .C(n11), .D(n10), .E(n4), .Z(n9) );
  HS65_LS_OA12X9 U7 ( .A(cnt[0]), .B(cnt[2]), .C(enable), .Z(n10) );
  HS65_LS_OAI22X6 U8 ( .A(enable), .B(n2), .C(cnt[0]), .D(n11), .Z(n5) );
  HS65_LS_IVX9 U9 ( .A(cnt[0]), .Z(n2) );
  HS65_LS_IVX9 U10 ( .A(cnt[1]), .Z(n4) );
  HS65_LS_IVX9 U11 ( .A(cnt[2]), .Z(n3) );
endmodule


module bram_DATA16_ADDR2_4 ( clk, reset, rd_addr, wr_addr, wr_data, wr_ena, 
        rd_data );
  input [1:0] rd_addr;
  input [1:0] wr_addr;
  input [15:0] wr_data;
  output [15:0] rd_data;
  input clk, reset, wr_ena;
  wire   \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] ,
         \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][15] , \mem[1][14] , \mem[1][13] ,
         \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] , \mem[1][8] ,
         \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] ,
         \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][15] , \mem[0][14] ,
         \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] ,
         \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] ,
         \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, n1,
         n2, n3, n4, n5, n6, n7, n8, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162;

  HS65_LS_DFPRQX9 \mem_reg[3][15]  ( .D(n91), .CP(clk), .RN(n1), .Q(
        \mem[3][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][14]  ( .D(n92), .CP(clk), .RN(n1), .Q(
        \mem[3][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][13]  ( .D(n93), .CP(clk), .RN(n1), .Q(
        \mem[3][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][12]  ( .D(n94), .CP(clk), .RN(n1), .Q(
        \mem[3][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][11]  ( .D(n95), .CP(clk), .RN(n1), .Q(
        \mem[3][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][10]  ( .D(n96), .CP(clk), .RN(n1), .Q(
        \mem[3][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][9]  ( .D(n97), .CP(clk), .RN(n1), .Q(\mem[3][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][8]  ( .D(n98), .CP(clk), .RN(n1), .Q(\mem[3][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][7]  ( .D(n99), .CP(clk), .RN(n1), .Q(\mem[3][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][6]  ( .D(n100), .CP(clk), .RN(n1), .Q(
        \mem[3][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][5]  ( .D(n101), .CP(clk), .RN(n1), .Q(
        \mem[3][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][4]  ( .D(n102), .CP(clk), .RN(n1), .Q(
        \mem[3][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][3]  ( .D(n103), .CP(clk), .RN(n1), .Q(
        \mem[3][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][2]  ( .D(n104), .CP(clk), .RN(n2), .Q(
        \mem[3][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][1]  ( .D(n105), .CP(clk), .RN(n2), .Q(
        \mem[3][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][0]  ( .D(n106), .CP(clk), .RN(n2), .Q(
        \mem[3][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][15]  ( .D(n107), .CP(clk), .RN(n2), .Q(
        \mem[2][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][14]  ( .D(n108), .CP(clk), .RN(n2), .Q(
        \mem[2][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][13]  ( .D(n109), .CP(clk), .RN(n2), .Q(
        \mem[2][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][12]  ( .D(n110), .CP(clk), .RN(n2), .Q(
        \mem[2][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][11]  ( .D(n111), .CP(clk), .RN(n2), .Q(
        \mem[2][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][10]  ( .D(n112), .CP(clk), .RN(n2), .Q(
        \mem[2][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][9]  ( .D(n113), .CP(clk), .RN(n2), .Q(
        \mem[2][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][8]  ( .D(n114), .CP(clk), .RN(n2), .Q(
        \mem[2][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][7]  ( .D(n115), .CP(clk), .RN(n2), .Q(
        \mem[2][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][6]  ( .D(n116), .CP(clk), .RN(n2), .Q(
        \mem[2][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][5]  ( .D(n117), .CP(clk), .RN(n3), .Q(
        \mem[2][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][4]  ( .D(n118), .CP(clk), .RN(n3), .Q(
        \mem[2][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][3]  ( .D(n119), .CP(clk), .RN(n3), .Q(
        \mem[2][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][2]  ( .D(n120), .CP(clk), .RN(n3), .Q(
        \mem[2][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][1]  ( .D(n121), .CP(clk), .RN(n3), .Q(
        \mem[2][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][0]  ( .D(n122), .CP(clk), .RN(n3), .Q(
        \mem[2][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][15]  ( .D(n123), .CP(clk), .RN(n3), .Q(
        \mem[1][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][14]  ( .D(n124), .CP(clk), .RN(n3), .Q(
        \mem[1][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][13]  ( .D(n125), .CP(clk), .RN(n3), .Q(
        \mem[1][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][12]  ( .D(n126), .CP(clk), .RN(n3), .Q(
        \mem[1][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][11]  ( .D(n127), .CP(clk), .RN(n3), .Q(
        \mem[1][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][10]  ( .D(n128), .CP(clk), .RN(n3), .Q(
        \mem[1][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][9]  ( .D(n129), .CP(clk), .RN(n3), .Q(
        \mem[1][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][8]  ( .D(n130), .CP(clk), .RN(n4), .Q(
        \mem[1][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][7]  ( .D(n131), .CP(clk), .RN(n4), .Q(
        \mem[1][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][6]  ( .D(n132), .CP(clk), .RN(n4), .Q(
        \mem[1][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][5]  ( .D(n133), .CP(clk), .RN(n4), .Q(
        \mem[1][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][4]  ( .D(n134), .CP(clk), .RN(n4), .Q(
        \mem[1][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][3]  ( .D(n135), .CP(clk), .RN(n4), .Q(
        \mem[1][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][2]  ( .D(n136), .CP(clk), .RN(n4), .Q(
        \mem[1][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][1]  ( .D(n137), .CP(clk), .RN(n4), .Q(
        \mem[1][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][0]  ( .D(n138), .CP(clk), .RN(n4), .Q(
        \mem[1][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][15]  ( .D(n139), .CP(clk), .RN(n4), .Q(
        \mem[0][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][14]  ( .D(n140), .CP(clk), .RN(n4), .Q(
        \mem[0][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][13]  ( .D(n141), .CP(clk), .RN(n4), .Q(
        \mem[0][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][12]  ( .D(n142), .CP(clk), .RN(n4), .Q(
        \mem[0][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][11]  ( .D(n143), .CP(clk), .RN(n5), .Q(
        \mem[0][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][10]  ( .D(n144), .CP(clk), .RN(n5), .Q(
        \mem[0][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][9]  ( .D(n145), .CP(clk), .RN(n5), .Q(
        \mem[0][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][8]  ( .D(n146), .CP(clk), .RN(n5), .Q(
        \mem[0][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][7]  ( .D(n147), .CP(clk), .RN(n5), .Q(
        \mem[0][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][6]  ( .D(n148), .CP(clk), .RN(n5), .Q(
        \mem[0][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][5]  ( .D(n149), .CP(clk), .RN(n5), .Q(
        \mem[0][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][4]  ( .D(n150), .CP(clk), .RN(n5), .Q(
        \mem[0][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][3]  ( .D(n151), .CP(clk), .RN(n5), .Q(
        \mem[0][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][2]  ( .D(n152), .CP(clk), .RN(n5), .Q(
        \mem[0][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][1]  ( .D(n153), .CP(clk), .RN(n5), .Q(
        \mem[0][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][0]  ( .D(n154), .CP(clk), .RN(n5), .Q(
        \mem[0][0] ) );
  HS65_LS_DFPRQX9 \rd_data_reg[15]  ( .D(N17), .CP(clk), .RN(n5), .Q(
        rd_data[15]) );
  HS65_LS_DFPRQX9 \rd_data_reg[14]  ( .D(N18), .CP(clk), .RN(n6), .Q(
        rd_data[14]) );
  HS65_LS_DFPRQX9 \rd_data_reg[13]  ( .D(N19), .CP(clk), .RN(n6), .Q(
        rd_data[13]) );
  HS65_LS_DFPRQX9 \rd_data_reg[12]  ( .D(N20), .CP(clk), .RN(n6), .Q(
        rd_data[12]) );
  HS65_LS_DFPRQX9 \rd_data_reg[11]  ( .D(N21), .CP(clk), .RN(n6), .Q(
        rd_data[11]) );
  HS65_LS_DFPRQX9 \rd_data_reg[10]  ( .D(N22), .CP(clk), .RN(n6), .Q(
        rd_data[10]) );
  HS65_LS_DFPRQX9 \rd_data_reg[9]  ( .D(N23), .CP(clk), .RN(n6), .Q(rd_data[9]) );
  HS65_LS_DFPRQX9 \rd_data_reg[8]  ( .D(N24), .CP(clk), .RN(n6), .Q(rd_data[8]) );
  HS65_LS_DFPRQX9 \rd_data_reg[7]  ( .D(N25), .CP(clk), .RN(n6), .Q(rd_data[7]) );
  HS65_LS_DFPRQX9 \rd_data_reg[6]  ( .D(N26), .CP(clk), .RN(n6), .Q(rd_data[6]) );
  HS65_LS_DFPRQX9 \rd_data_reg[5]  ( .D(N27), .CP(clk), .RN(n6), .Q(rd_data[5]) );
  HS65_LS_DFPRQX9 \rd_data_reg[4]  ( .D(N28), .CP(clk), .RN(n6), .Q(rd_data[4]) );
  HS65_LS_DFPRQX9 \rd_data_reg[3]  ( .D(N29), .CP(clk), .RN(n6), .Q(rd_data[3]) );
  HS65_LS_DFPRQX9 \rd_data_reg[2]  ( .D(N30), .CP(clk), .RN(n6), .Q(rd_data[2]) );
  HS65_LS_DFPRQX9 \rd_data_reg[1]  ( .D(N31), .CP(clk), .RN(n7), .Q(rd_data[1]) );
  HS65_LS_DFPRQX9 \rd_data_reg[0]  ( .D(N32), .CP(clk), .RN(n7), .Q(rd_data[0]) );
  HS65_LS_BFX9 U3 ( .A(n81), .Z(n4) );
  HS65_LS_BFX9 U4 ( .A(n81), .Z(n3) );
  HS65_LS_BFX9 U5 ( .A(n81), .Z(n2) );
  HS65_LS_BFX9 U6 ( .A(n83), .Z(n81) );
  HS65_LS_BFX9 U7 ( .A(n8), .Z(n6) );
  HS65_LS_BFX9 U8 ( .A(n8), .Z(n5) );
  HS65_LS_BFX9 U9 ( .A(n82), .Z(n1) );
  HS65_LS_BFX9 U10 ( .A(n83), .Z(n82) );
  HS65_LS_BFX9 U11 ( .A(n8), .Z(n7) );
  HS65_LS_BFX9 U12 ( .A(n83), .Z(n8) );
  HS65_LS_IVX9 U13 ( .A(reset), .Z(n83) );
  HS65_LS_IVX9 U14 ( .A(n161), .Z(n86) );
  HS65_LS_IVX9 U15 ( .A(n162), .Z(n87) );
  HS65_LS_NAND3X5 U16 ( .A(wr_ena), .B(n88), .C(wr_addr[0]), .Z(n161) );
  HS65_LS_IVX9 U17 ( .A(wr_addr[0]), .Z(n89) );
  HS65_LS_NAND3X5 U18 ( .A(n89), .B(n88), .C(wr_ena), .Z(n162) );
  HS65_LS_IVX9 U19 ( .A(n160), .Z(n85) );
  HS65_LS_IVX9 U20 ( .A(n159), .Z(n84) );
  HS65_LS_NAND3X5 U21 ( .A(wr_ena), .B(n89), .C(wr_addr[1]), .Z(n160) );
  HS65_LS_NOR2X6 U22 ( .A(n90), .B(rd_addr[1]), .Z(n157) );
  HS65_LS_NOR2X6 U23 ( .A(rd_addr[0]), .B(rd_addr[1]), .Z(n158) );
  HS65_LS_IVX9 U24 ( .A(wr_addr[1]), .Z(n88) );
  HS65_LS_NAND3X5 U25 ( .A(wr_addr[0]), .B(wr_ena), .C(wr_addr[1]), .Z(n159)
         );
  HS65_LS_AND2X4 U26 ( .A(rd_addr[1]), .B(n90), .Z(n156) );
  HS65_LS_IVX9 U27 ( .A(rd_addr[0]), .Z(n90) );
  HS65_LS_AND2X4 U28 ( .A(rd_addr[1]), .B(rd_addr[0]), .Z(n155) );
  HS65_LS_MX41X7 U29 ( .D0(n158), .S0(\mem[0][0] ), .D1(n157), .S1(\mem[1][0] ), .D2(n156), .S2(\mem[2][0] ), .D3(n155), .S3(\mem[3][0] ), .Z(N32) );
  HS65_LS_MX41X7 U30 ( .D0(n158), .S0(\mem[0][1] ), .D1(n157), .S1(\mem[1][1] ), .D2(n156), .S2(\mem[2][1] ), .D3(n155), .S3(\mem[3][1] ), .Z(N31) );
  HS65_LS_MX41X7 U31 ( .D0(n158), .S0(\mem[0][2] ), .D1(n157), .S1(\mem[1][2] ), .D2(n156), .S2(\mem[2][2] ), .D3(n155), .S3(\mem[3][2] ), .Z(N30) );
  HS65_LS_MX41X7 U32 ( .D0(n158), .S0(\mem[0][3] ), .D1(n157), .S1(\mem[1][3] ), .D2(n156), .S2(\mem[2][3] ), .D3(n155), .S3(\mem[3][3] ), .Z(N29) );
  HS65_LS_MX41X7 U33 ( .D0(n158), .S0(\mem[0][4] ), .D1(n157), .S1(\mem[1][4] ), .D2(n156), .S2(\mem[2][4] ), .D3(n155), .S3(\mem[3][4] ), .Z(N28) );
  HS65_LS_MX41X7 U34 ( .D0(n158), .S0(\mem[0][5] ), .D1(n157), .S1(\mem[1][5] ), .D2(n156), .S2(\mem[2][5] ), .D3(n155), .S3(\mem[3][5] ), .Z(N27) );
  HS65_LS_MX41X7 U35 ( .D0(n158), .S0(\mem[0][6] ), .D1(n157), .S1(\mem[1][6] ), .D2(n156), .S2(\mem[2][6] ), .D3(n155), .S3(\mem[3][6] ), .Z(N26) );
  HS65_LS_MX41X7 U36 ( .D0(n158), .S0(\mem[0][7] ), .D1(n157), .S1(\mem[1][7] ), .D2(n156), .S2(\mem[2][7] ), .D3(n155), .S3(\mem[3][7] ), .Z(N25) );
  HS65_LS_MX41X7 U37 ( .D0(n158), .S0(\mem[0][8] ), .D1(n157), .S1(\mem[1][8] ), .D2(n156), .S2(\mem[2][8] ), .D3(n155), .S3(\mem[3][8] ), .Z(N24) );
  HS65_LS_MX41X7 U38 ( .D0(n158), .S0(\mem[0][9] ), .D1(n157), .S1(\mem[1][9] ), .D2(n156), .S2(\mem[2][9] ), .D3(n155), .S3(\mem[3][9] ), .Z(N23) );
  HS65_LS_MX41X7 U39 ( .D0(n158), .S0(\mem[0][10] ), .D1(n157), .S1(
        \mem[1][10] ), .D2(n156), .S2(\mem[2][10] ), .D3(n155), .S3(
        \mem[3][10] ), .Z(N22) );
  HS65_LS_MX41X7 U40 ( .D0(n158), .S0(\mem[0][11] ), .D1(n157), .S1(
        \mem[1][11] ), .D2(n156), .S2(\mem[2][11] ), .D3(n155), .S3(
        \mem[3][11] ), .Z(N21) );
  HS65_LS_MX41X7 U41 ( .D0(n158), .S0(\mem[0][12] ), .D1(n157), .S1(
        \mem[1][12] ), .D2(n156), .S2(\mem[2][12] ), .D3(n155), .S3(
        \mem[3][12] ), .Z(N20) );
  HS65_LS_MX41X7 U42 ( .D0(n158), .S0(\mem[0][13] ), .D1(n157), .S1(
        \mem[1][13] ), .D2(n156), .S2(\mem[2][13] ), .D3(n155), .S3(
        \mem[3][13] ), .Z(N19) );
  HS65_LS_MX41X7 U43 ( .D0(n158), .S0(\mem[0][14] ), .D1(n157), .S1(
        \mem[1][14] ), .D2(n156), .S2(\mem[2][14] ), .D3(n155), .S3(
        \mem[3][14] ), .Z(N18) );
  HS65_LS_MX41X7 U44 ( .D0(n158), .S0(\mem[0][15] ), .D1(n157), .S1(
        \mem[1][15] ), .D2(n156), .S2(\mem[2][15] ), .D3(n155), .S3(
        \mem[3][15] ), .Z(N17) );
  HS65_LS_AO22X9 U45 ( .A(wr_data[0]), .B(n86), .C(n161), .D(\mem[1][0] ), .Z(
        n138) );
  HS65_LS_AO22X9 U46 ( .A(wr_data[1]), .B(n86), .C(n161), .D(\mem[1][1] ), .Z(
        n137) );
  HS65_LS_AO22X9 U47 ( .A(wr_data[2]), .B(n86), .C(n161), .D(\mem[1][2] ), .Z(
        n136) );
  HS65_LS_AO22X9 U48 ( .A(wr_data[3]), .B(n86), .C(n161), .D(\mem[1][3] ), .Z(
        n135) );
  HS65_LS_AO22X9 U49 ( .A(wr_data[4]), .B(n86), .C(n161), .D(\mem[1][4] ), .Z(
        n134) );
  HS65_LS_AO22X9 U50 ( .A(wr_data[5]), .B(n86), .C(n161), .D(\mem[1][5] ), .Z(
        n133) );
  HS65_LS_AO22X9 U51 ( .A(wr_data[6]), .B(n86), .C(n161), .D(\mem[1][6] ), .Z(
        n132) );
  HS65_LS_AO22X9 U52 ( .A(wr_data[7]), .B(n86), .C(n161), .D(\mem[1][7] ), .Z(
        n131) );
  HS65_LS_AO22X9 U53 ( .A(wr_data[8]), .B(n86), .C(n161), .D(\mem[1][8] ), .Z(
        n130) );
  HS65_LS_AO22X9 U54 ( .A(wr_data[9]), .B(n86), .C(n161), .D(\mem[1][9] ), .Z(
        n129) );
  HS65_LS_AO22X9 U55 ( .A(wr_data[10]), .B(n86), .C(n161), .D(\mem[1][10] ), 
        .Z(n128) );
  HS65_LS_AO22X9 U56 ( .A(wr_data[11]), .B(n86), .C(n161), .D(\mem[1][11] ), 
        .Z(n127) );
  HS65_LS_AO22X9 U57 ( .A(wr_data[12]), .B(n86), .C(n161), .D(\mem[1][12] ), 
        .Z(n126) );
  HS65_LS_AO22X9 U58 ( .A(wr_data[13]), .B(n86), .C(n161), .D(\mem[1][13] ), 
        .Z(n125) );
  HS65_LS_AO22X9 U59 ( .A(wr_data[14]), .B(n86), .C(n161), .D(\mem[1][14] ), 
        .Z(n124) );
  HS65_LS_AO22X9 U60 ( .A(wr_data[15]), .B(n86), .C(n161), .D(\mem[1][15] ), 
        .Z(n123) );
  HS65_LS_AO22X9 U61 ( .A(wr_data[0]), .B(n85), .C(n160), .D(\mem[2][0] ), .Z(
        n122) );
  HS65_LS_AO22X9 U62 ( .A(wr_data[1]), .B(n85), .C(n160), .D(\mem[2][1] ), .Z(
        n121) );
  HS65_LS_AO22X9 U63 ( .A(wr_data[2]), .B(n85), .C(n160), .D(\mem[2][2] ), .Z(
        n120) );
  HS65_LS_AO22X9 U64 ( .A(wr_data[3]), .B(n85), .C(n160), .D(\mem[2][3] ), .Z(
        n119) );
  HS65_LS_AO22X9 U65 ( .A(wr_data[4]), .B(n85), .C(n160), .D(\mem[2][4] ), .Z(
        n118) );
  HS65_LS_AO22X9 U66 ( .A(wr_data[5]), .B(n85), .C(n160), .D(\mem[2][5] ), .Z(
        n117) );
  HS65_LS_AO22X9 U67 ( .A(wr_data[6]), .B(n85), .C(n160), .D(\mem[2][6] ), .Z(
        n116) );
  HS65_LS_AO22X9 U68 ( .A(wr_data[7]), .B(n85), .C(n160), .D(\mem[2][7] ), .Z(
        n115) );
  HS65_LS_AO22X9 U69 ( .A(wr_data[8]), .B(n85), .C(n160), .D(\mem[2][8] ), .Z(
        n114) );
  HS65_LS_AO22X9 U70 ( .A(wr_data[9]), .B(n85), .C(n160), .D(\mem[2][9] ), .Z(
        n113) );
  HS65_LS_AO22X9 U71 ( .A(wr_data[10]), .B(n85), .C(n160), .D(\mem[2][10] ), 
        .Z(n112) );
  HS65_LS_AO22X9 U72 ( .A(wr_data[11]), .B(n85), .C(n160), .D(\mem[2][11] ), 
        .Z(n111) );
  HS65_LS_AO22X9 U73 ( .A(wr_data[12]), .B(n85), .C(n160), .D(\mem[2][12] ), 
        .Z(n110) );
  HS65_LS_AO22X9 U74 ( .A(wr_data[13]), .B(n85), .C(n160), .D(\mem[2][13] ), 
        .Z(n109) );
  HS65_LS_AO22X9 U75 ( .A(wr_data[14]), .B(n85), .C(n160), .D(\mem[2][14] ), 
        .Z(n108) );
  HS65_LS_AO22X9 U76 ( .A(wr_data[15]), .B(n85), .C(n160), .D(\mem[2][15] ), 
        .Z(n107) );
  HS65_LS_AO22X9 U77 ( .A(n87), .B(wr_data[0]), .C(n162), .D(\mem[0][0] ), .Z(
        n154) );
  HS65_LS_AO22X9 U78 ( .A(n87), .B(wr_data[1]), .C(n162), .D(\mem[0][1] ), .Z(
        n153) );
  HS65_LS_AO22X9 U79 ( .A(n87), .B(wr_data[2]), .C(n162), .D(\mem[0][2] ), .Z(
        n152) );
  HS65_LS_AO22X9 U80 ( .A(n87), .B(wr_data[3]), .C(n162), .D(\mem[0][3] ), .Z(
        n151) );
  HS65_LS_AO22X9 U81 ( .A(n87), .B(wr_data[4]), .C(n162), .D(\mem[0][4] ), .Z(
        n150) );
  HS65_LS_AO22X9 U82 ( .A(n87), .B(wr_data[5]), .C(n162), .D(\mem[0][5] ), .Z(
        n149) );
  HS65_LS_AO22X9 U83 ( .A(n87), .B(wr_data[6]), .C(n162), .D(\mem[0][6] ), .Z(
        n148) );
  HS65_LS_AO22X9 U84 ( .A(n87), .B(wr_data[7]), .C(n162), .D(\mem[0][7] ), .Z(
        n147) );
  HS65_LS_AO22X9 U85 ( .A(n87), .B(wr_data[8]), .C(n162), .D(\mem[0][8] ), .Z(
        n146) );
  HS65_LS_AO22X9 U86 ( .A(n87), .B(wr_data[9]), .C(n162), .D(\mem[0][9] ), .Z(
        n145) );
  HS65_LS_AO22X9 U87 ( .A(n87), .B(wr_data[10]), .C(n162), .D(\mem[0][10] ), 
        .Z(n144) );
  HS65_LS_AO22X9 U88 ( .A(n87), .B(wr_data[11]), .C(n162), .D(\mem[0][11] ), 
        .Z(n143) );
  HS65_LS_AO22X9 U89 ( .A(n87), .B(wr_data[12]), .C(n162), .D(\mem[0][12] ), 
        .Z(n142) );
  HS65_LS_AO22X9 U90 ( .A(n87), .B(wr_data[13]), .C(n162), .D(\mem[0][13] ), 
        .Z(n141) );
  HS65_LS_AO22X9 U91 ( .A(n87), .B(wr_data[14]), .C(n162), .D(\mem[0][14] ), 
        .Z(n140) );
  HS65_LS_AO22X9 U92 ( .A(n87), .B(wr_data[15]), .C(n162), .D(\mem[0][15] ), 
        .Z(n139) );
  HS65_LS_AO22X9 U93 ( .A(wr_data[0]), .B(n84), .C(n159), .D(\mem[3][0] ), .Z(
        n106) );
  HS65_LS_AO22X9 U94 ( .A(wr_data[1]), .B(n84), .C(n159), .D(\mem[3][1] ), .Z(
        n105) );
  HS65_LS_AO22X9 U95 ( .A(wr_data[2]), .B(n84), .C(n159), .D(\mem[3][2] ), .Z(
        n104) );
  HS65_LS_AO22X9 U96 ( .A(wr_data[3]), .B(n84), .C(n159), .D(\mem[3][3] ), .Z(
        n103) );
  HS65_LS_AO22X9 U97 ( .A(wr_data[4]), .B(n84), .C(n159), .D(\mem[3][4] ), .Z(
        n102) );
  HS65_LS_AO22X9 U98 ( .A(wr_data[5]), .B(n84), .C(n159), .D(\mem[3][5] ), .Z(
        n101) );
  HS65_LS_AO22X9 U99 ( .A(wr_data[6]), .B(n84), .C(n159), .D(\mem[3][6] ), .Z(
        n100) );
  HS65_LS_AO22X9 U100 ( .A(wr_data[7]), .B(n84), .C(n159), .D(\mem[3][7] ), 
        .Z(n99) );
  HS65_LS_AO22X9 U101 ( .A(wr_data[8]), .B(n84), .C(n159), .D(\mem[3][8] ), 
        .Z(n98) );
  HS65_LS_AO22X9 U102 ( .A(wr_data[9]), .B(n84), .C(n159), .D(\mem[3][9] ), 
        .Z(n97) );
  HS65_LS_AO22X9 U103 ( .A(wr_data[10]), .B(n84), .C(n159), .D(\mem[3][10] ), 
        .Z(n96) );
  HS65_LS_AO22X9 U104 ( .A(wr_data[11]), .B(n84), .C(n159), .D(\mem[3][11] ), 
        .Z(n95) );
  HS65_LS_AO22X9 U105 ( .A(wr_data[12]), .B(n84), .C(n159), .D(\mem[3][12] ), 
        .Z(n94) );
  HS65_LS_AO22X9 U106 ( .A(wr_data[13]), .B(n84), .C(n159), .D(\mem[3][13] ), 
        .Z(n93) );
  HS65_LS_AO22X9 U107 ( .A(wr_data[14]), .B(n84), .C(n159), .D(\mem[3][14] ), 
        .Z(n92) );
  HS65_LS_AO22X9 U108 ( .A(wr_data[15]), .B(n84), .C(n159), .D(\mem[3][15] ), 
        .Z(n91) );
endmodule


module bram_DATA32_ADDR2_2 ( clk, reset, rd_addr, wr_addr, wr_data, wr_ena, 
        rd_data );
  input [1:0] rd_addr;
  input [1:0] wr_addr;
  input [31:0] wr_data;
  output [31:0] rd_data;
  input clk, reset, wr_ena;
  wire   \mem[3][31] , \mem[3][30] , \mem[3][29] , \mem[3][28] , \mem[3][27] ,
         \mem[3][26] , \mem[3][25] , \mem[3][24] , \mem[3][23] , \mem[3][22] ,
         \mem[3][21] , \mem[3][20] , \mem[3][19] , \mem[3][18] , \mem[3][17] ,
         \mem[3][16] , \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] ,
         \mem[3][11] , \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] ,
         \mem[3][6] , \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] ,
         \mem[3][1] , \mem[3][0] , \mem[2][31] , \mem[2][30] , \mem[2][29] ,
         \mem[2][28] , \mem[2][27] , \mem[2][26] , \mem[2][25] , \mem[2][24] ,
         \mem[2][23] , \mem[2][22] , \mem[2][21] , \mem[2][20] , \mem[2][19] ,
         \mem[2][18] , \mem[2][17] , \mem[2][16] , \mem[2][15] , \mem[2][14] ,
         \mem[2][13] , \mem[2][12] , \mem[2][11] , \mem[2][10] , \mem[2][9] ,
         \mem[2][8] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][31] ,
         \mem[1][30] , \mem[1][29] , \mem[1][28] , \mem[1][27] , \mem[1][26] ,
         \mem[1][25] , \mem[1][24] , \mem[1][23] , \mem[1][22] , \mem[1][21] ,
         \mem[1][20] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][31] , \mem[0][30] , \mem[0][29] , \mem[0][28] ,
         \mem[0][27] , \mem[0][26] , \mem[0][25] , \mem[0][24] , \mem[0][23] ,
         \mem[0][22] , \mem[0][21] , \mem[0][20] , \mem[0][19] , \mem[0][18] ,
         \mem[0][17] , \mem[0][16] , \mem[0][15] , \mem[0][14] , \mem[0][13] ,
         \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] , \mem[0][8] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N17, N18, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36,
         N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327;

  HS65_LS_DFPRQX9 \mem_reg[3][31]  ( .D(n193), .CP(clk), .RN(n171), .Q(
        \mem[3][31] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][30]  ( .D(n194), .CP(clk), .RN(n171), .Q(
        \mem[3][30] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][29]  ( .D(n195), .CP(clk), .RN(n171), .Q(
        \mem[3][29] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][28]  ( .D(n196), .CP(clk), .RN(n171), .Q(
        \mem[3][28] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][27]  ( .D(n197), .CP(clk), .RN(n171), .Q(
        \mem[3][27] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][26]  ( .D(n198), .CP(clk), .RN(n171), .Q(
        \mem[3][26] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][25]  ( .D(n199), .CP(clk), .RN(n171), .Q(
        \mem[3][25] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][24]  ( .D(n200), .CP(clk), .RN(n171), .Q(
        \mem[3][24] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][23]  ( .D(n201), .CP(clk), .RN(n171), .Q(
        \mem[3][23] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][22]  ( .D(n202), .CP(clk), .RN(n171), .Q(
        \mem[3][22] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][21]  ( .D(n203), .CP(clk), .RN(n171), .Q(
        \mem[3][21] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][20]  ( .D(n204), .CP(clk), .RN(n171), .Q(
        \mem[3][20] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][19]  ( .D(n205), .CP(clk), .RN(n171), .Q(
        \mem[3][19] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][18]  ( .D(n206), .CP(clk), .RN(n172), .Q(
        \mem[3][18] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][17]  ( .D(n207), .CP(clk), .RN(n172), .Q(
        \mem[3][17] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][16]  ( .D(n208), .CP(clk), .RN(n172), .Q(
        \mem[3][16] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][15]  ( .D(n209), .CP(clk), .RN(n172), .Q(
        \mem[3][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][14]  ( .D(n210), .CP(clk), .RN(n172), .Q(
        \mem[3][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][13]  ( .D(n211), .CP(clk), .RN(n172), .Q(
        \mem[3][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][12]  ( .D(n212), .CP(clk), .RN(n172), .Q(
        \mem[3][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][11]  ( .D(n213), .CP(clk), .RN(n172), .Q(
        \mem[3][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][10]  ( .D(n214), .CP(clk), .RN(n172), .Q(
        \mem[3][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][9]  ( .D(n215), .CP(clk), .RN(n172), .Q(
        \mem[3][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][8]  ( .D(n216), .CP(clk), .RN(n172), .Q(
        \mem[3][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][7]  ( .D(n217), .CP(clk), .RN(n172), .Q(
        \mem[3][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][6]  ( .D(n218), .CP(clk), .RN(n172), .Q(
        \mem[3][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][5]  ( .D(n219), .CP(clk), .RN(n173), .Q(
        \mem[3][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][4]  ( .D(n220), .CP(clk), .RN(n173), .Q(
        \mem[3][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][3]  ( .D(n221), .CP(clk), .RN(n173), .Q(
        \mem[3][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][2]  ( .D(n222), .CP(clk), .RN(n173), .Q(
        \mem[3][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][1]  ( .D(n223), .CP(clk), .RN(n173), .Q(
        \mem[3][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][0]  ( .D(n224), .CP(clk), .RN(n173), .Q(
        \mem[3][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][31]  ( .D(n225), .CP(clk), .RN(n173), .Q(
        \mem[2][31] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][30]  ( .D(n226), .CP(clk), .RN(n173), .Q(
        \mem[2][30] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][29]  ( .D(n227), .CP(clk), .RN(n173), .Q(
        \mem[2][29] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][28]  ( .D(n228), .CP(clk), .RN(n173), .Q(
        \mem[2][28] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][27]  ( .D(n229), .CP(clk), .RN(n173), .Q(
        \mem[2][27] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][26]  ( .D(n230), .CP(clk), .RN(n173), .Q(
        \mem[2][26] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][25]  ( .D(n231), .CP(clk), .RN(n173), .Q(
        \mem[2][25] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][24]  ( .D(n232), .CP(clk), .RN(n174), .Q(
        \mem[2][24] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][23]  ( .D(n233), .CP(clk), .RN(n174), .Q(
        \mem[2][23] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][22]  ( .D(n234), .CP(clk), .RN(n174), .Q(
        \mem[2][22] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][21]  ( .D(n235), .CP(clk), .RN(n174), .Q(
        \mem[2][21] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][20]  ( .D(n236), .CP(clk), .RN(n174), .Q(
        \mem[2][20] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][19]  ( .D(n237), .CP(clk), .RN(n174), .Q(
        \mem[2][19] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][18]  ( .D(n238), .CP(clk), .RN(n174), .Q(
        \mem[2][18] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][17]  ( .D(n239), .CP(clk), .RN(n174), .Q(
        \mem[2][17] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][16]  ( .D(n240), .CP(clk), .RN(n174), .Q(
        \mem[2][16] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][15]  ( .D(n241), .CP(clk), .RN(n174), .Q(
        \mem[2][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][14]  ( .D(n242), .CP(clk), .RN(n174), .Q(
        \mem[2][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][13]  ( .D(n243), .CP(clk), .RN(n174), .Q(
        \mem[2][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][12]  ( .D(n244), .CP(clk), .RN(n174), .Q(
        \mem[2][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][11]  ( .D(n245), .CP(clk), .RN(n175), .Q(
        \mem[2][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][10]  ( .D(n246), .CP(clk), .RN(n175), .Q(
        \mem[2][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][9]  ( .D(n247), .CP(clk), .RN(n175), .Q(
        \mem[2][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][8]  ( .D(n248), .CP(clk), .RN(n175), .Q(
        \mem[2][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][7]  ( .D(n249), .CP(clk), .RN(n175), .Q(
        \mem[2][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][6]  ( .D(n250), .CP(clk), .RN(n175), .Q(
        \mem[2][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][5]  ( .D(n251), .CP(clk), .RN(n175), .Q(
        \mem[2][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][4]  ( .D(n252), .CP(clk), .RN(n175), .Q(
        \mem[2][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][3]  ( .D(n253), .CP(clk), .RN(n175), .Q(
        \mem[2][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][2]  ( .D(n254), .CP(clk), .RN(n175), .Q(
        \mem[2][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][1]  ( .D(n255), .CP(clk), .RN(n175), .Q(
        \mem[2][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][0]  ( .D(n256), .CP(clk), .RN(n175), .Q(
        \mem[2][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][31]  ( .D(n257), .CP(clk), .RN(n175), .Q(
        \mem[1][31] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][30]  ( .D(n258), .CP(clk), .RN(n176), .Q(
        \mem[1][30] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][29]  ( .D(n259), .CP(clk), .RN(n176), .Q(
        \mem[1][29] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][28]  ( .D(n260), .CP(clk), .RN(n176), .Q(
        \mem[1][28] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][27]  ( .D(n261), .CP(clk), .RN(n176), .Q(
        \mem[1][27] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][26]  ( .D(n262), .CP(clk), .RN(n176), .Q(
        \mem[1][26] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][25]  ( .D(n263), .CP(clk), .RN(n176), .Q(
        \mem[1][25] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][24]  ( .D(n264), .CP(clk), .RN(n176), .Q(
        \mem[1][24] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][23]  ( .D(n265), .CP(clk), .RN(n176), .Q(
        \mem[1][23] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][22]  ( .D(n266), .CP(clk), .RN(n176), .Q(
        \mem[1][22] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][21]  ( .D(n267), .CP(clk), .RN(n176), .Q(
        \mem[1][21] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][20]  ( .D(n268), .CP(clk), .RN(n176), .Q(
        \mem[1][20] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][19]  ( .D(n269), .CP(clk), .RN(n176), .Q(
        \mem[1][19] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][18]  ( .D(n270), .CP(clk), .RN(n176), .Q(
        \mem[1][18] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][17]  ( .D(n271), .CP(clk), .RN(n177), .Q(
        \mem[1][17] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][16]  ( .D(n272), .CP(clk), .RN(n177), .Q(
        \mem[1][16] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][15]  ( .D(n273), .CP(clk), .RN(n177), .Q(
        \mem[1][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][14]  ( .D(n274), .CP(clk), .RN(n177), .Q(
        \mem[1][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][13]  ( .D(n275), .CP(clk), .RN(n177), .Q(
        \mem[1][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][12]  ( .D(n276), .CP(clk), .RN(n177), .Q(
        \mem[1][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][11]  ( .D(n277), .CP(clk), .RN(n177), .Q(
        \mem[1][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][10]  ( .D(n278), .CP(clk), .RN(n177), .Q(
        \mem[1][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][9]  ( .D(n279), .CP(clk), .RN(n177), .Q(
        \mem[1][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][8]  ( .D(n280), .CP(clk), .RN(n177), .Q(
        \mem[1][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][7]  ( .D(n281), .CP(clk), .RN(n177), .Q(
        \mem[1][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][6]  ( .D(n282), .CP(clk), .RN(n177), .Q(
        \mem[1][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][5]  ( .D(n283), .CP(clk), .RN(n177), .Q(
        \mem[1][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][4]  ( .D(n284), .CP(clk), .RN(n178), .Q(
        \mem[1][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][3]  ( .D(n285), .CP(clk), .RN(n178), .Q(
        \mem[1][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][2]  ( .D(n286), .CP(clk), .RN(n178), .Q(
        \mem[1][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][1]  ( .D(n287), .CP(clk), .RN(n178), .Q(
        \mem[1][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][0]  ( .D(n288), .CP(clk), .RN(n178), .Q(
        \mem[1][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][31]  ( .D(n289), .CP(clk), .RN(n178), .Q(
        \mem[0][31] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][30]  ( .D(n290), .CP(clk), .RN(n178), .Q(
        \mem[0][30] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][29]  ( .D(n291), .CP(clk), .RN(n178), .Q(
        \mem[0][29] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][28]  ( .D(n292), .CP(clk), .RN(n178), .Q(
        \mem[0][28] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][27]  ( .D(n293), .CP(clk), .RN(n178), .Q(
        \mem[0][27] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][26]  ( .D(n294), .CP(clk), .RN(n178), .Q(
        \mem[0][26] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][25]  ( .D(n295), .CP(clk), .RN(n178), .Q(
        \mem[0][25] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][24]  ( .D(n296), .CP(clk), .RN(n178), .Q(
        \mem[0][24] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][23]  ( .D(n297), .CP(clk), .RN(n179), .Q(
        \mem[0][23] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][22]  ( .D(n298), .CP(clk), .RN(n179), .Q(
        \mem[0][22] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][21]  ( .D(n299), .CP(clk), .RN(n179), .Q(
        \mem[0][21] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][20]  ( .D(n300), .CP(clk), .RN(n179), .Q(
        \mem[0][20] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][19]  ( .D(n301), .CP(clk), .RN(n179), .Q(
        \mem[0][19] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][18]  ( .D(n302), .CP(clk), .RN(n179), .Q(
        \mem[0][18] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][17]  ( .D(n303), .CP(clk), .RN(n179), .Q(
        \mem[0][17] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][16]  ( .D(n304), .CP(clk), .RN(n179), .Q(
        \mem[0][16] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][15]  ( .D(n305), .CP(clk), .RN(n179), .Q(
        \mem[0][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][14]  ( .D(n306), .CP(clk), .RN(n179), .Q(
        \mem[0][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][13]  ( .D(n307), .CP(clk), .RN(n179), .Q(
        \mem[0][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][12]  ( .D(n308), .CP(clk), .RN(n179), .Q(
        \mem[0][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][11]  ( .D(n309), .CP(clk), .RN(n179), .Q(
        \mem[0][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][10]  ( .D(n310), .CP(clk), .RN(n180), .Q(
        \mem[0][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][9]  ( .D(n311), .CP(clk), .RN(n180), .Q(
        \mem[0][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][8]  ( .D(n312), .CP(clk), .RN(n180), .Q(
        \mem[0][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][7]  ( .D(n313), .CP(clk), .RN(n180), .Q(
        \mem[0][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][6]  ( .D(n314), .CP(clk), .RN(n180), .Q(
        \mem[0][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][5]  ( .D(n315), .CP(clk), .RN(n180), .Q(
        \mem[0][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][4]  ( .D(n316), .CP(clk), .RN(n180), .Q(
        \mem[0][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][3]  ( .D(n317), .CP(clk), .RN(n180), .Q(
        \mem[0][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][2]  ( .D(n318), .CP(clk), .RN(n180), .Q(
        \mem[0][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][1]  ( .D(n319), .CP(clk), .RN(n180), .Q(
        \mem[0][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][0]  ( .D(n320), .CP(clk), .RN(n180), .Q(
        \mem[0][0] ) );
  HS65_LS_DFPRQX9 \rd_data_reg[31]  ( .D(N17), .CP(clk), .RN(n180), .Q(
        rd_data[31]) );
  HS65_LS_DFPRQX9 \rd_data_reg[30]  ( .D(N18), .CP(clk), .RN(n180), .Q(
        rd_data[30]) );
  HS65_LS_DFPRQX9 \rd_data_reg[29]  ( .D(N19), .CP(clk), .RN(n181), .Q(
        rd_data[29]) );
  HS65_LS_DFPRQX9 \rd_data_reg[28]  ( .D(N20), .CP(clk), .RN(n181), .Q(
        rd_data[28]) );
  HS65_LS_DFPRQX9 \rd_data_reg[27]  ( .D(N21), .CP(clk), .RN(n181), .Q(
        rd_data[27]) );
  HS65_LS_DFPRQX9 \rd_data_reg[26]  ( .D(N22), .CP(clk), .RN(n181), .Q(
        rd_data[26]) );
  HS65_LS_DFPRQX9 \rd_data_reg[25]  ( .D(N23), .CP(clk), .RN(n181), .Q(
        rd_data[25]) );
  HS65_LS_DFPRQX9 \rd_data_reg[24]  ( .D(N24), .CP(clk), .RN(n181), .Q(
        rd_data[24]) );
  HS65_LS_DFPRQX9 \rd_data_reg[23]  ( .D(N25), .CP(clk), .RN(n181), .Q(
        rd_data[23]) );
  HS65_LS_DFPRQX9 \rd_data_reg[22]  ( .D(N26), .CP(clk), .RN(n181), .Q(
        rd_data[22]) );
  HS65_LS_DFPRQX9 \rd_data_reg[21]  ( .D(N27), .CP(clk), .RN(n181), .Q(
        rd_data[21]) );
  HS65_LS_DFPRQX9 \rd_data_reg[20]  ( .D(N28), .CP(clk), .RN(n181), .Q(
        rd_data[20]) );
  HS65_LS_DFPRQX9 \rd_data_reg[19]  ( .D(N29), .CP(clk), .RN(n181), .Q(
        rd_data[19]) );
  HS65_LS_DFPRQX9 \rd_data_reg[18]  ( .D(N30), .CP(clk), .RN(n181), .Q(
        rd_data[18]) );
  HS65_LS_DFPRQX9 \rd_data_reg[17]  ( .D(N31), .CP(clk), .RN(n181), .Q(
        rd_data[17]) );
  HS65_LS_DFPRQX9 \rd_data_reg[16]  ( .D(N32), .CP(clk), .RN(n182), .Q(
        rd_data[16]) );
  HS65_LS_DFPRQX9 \rd_data_reg[15]  ( .D(N33), .CP(clk), .RN(n182), .Q(
        rd_data[15]) );
  HS65_LS_DFPRQX9 \rd_data_reg[14]  ( .D(N34), .CP(clk), .RN(n182), .Q(
        rd_data[14]) );
  HS65_LS_DFPRQX9 \rd_data_reg[13]  ( .D(N35), .CP(clk), .RN(n182), .Q(
        rd_data[13]) );
  HS65_LS_DFPRQX9 \rd_data_reg[12]  ( .D(N36), .CP(clk), .RN(n182), .Q(
        rd_data[12]) );
  HS65_LS_DFPRQX9 \rd_data_reg[11]  ( .D(N37), .CP(clk), .RN(n182), .Q(
        rd_data[11]) );
  HS65_LS_DFPRQX9 \rd_data_reg[10]  ( .D(N38), .CP(clk), .RN(n182), .Q(
        rd_data[10]) );
  HS65_LS_DFPRQX9 \rd_data_reg[9]  ( .D(N39), .CP(clk), .RN(n182), .Q(
        rd_data[9]) );
  HS65_LS_DFPRQX9 \rd_data_reg[8]  ( .D(N40), .CP(clk), .RN(n182), .Q(
        rd_data[8]) );
  HS65_LS_DFPRQX9 \rd_data_reg[7]  ( .D(N41), .CP(clk), .RN(n182), .Q(
        rd_data[7]) );
  HS65_LS_DFPRQX9 \rd_data_reg[6]  ( .D(N42), .CP(clk), .RN(n182), .Q(
        rd_data[6]) );
  HS65_LS_DFPRQX9 \rd_data_reg[5]  ( .D(N43), .CP(clk), .RN(n182), .Q(
        rd_data[5]) );
  HS65_LS_DFPRQX9 \rd_data_reg[4]  ( .D(N44), .CP(clk), .RN(n182), .Q(
        rd_data[4]) );
  HS65_LS_DFPRQX9 \rd_data_reg[3]  ( .D(N45), .CP(clk), .RN(n183), .Q(
        rd_data[3]) );
  HS65_LS_DFPRQX9 \rd_data_reg[2]  ( .D(N46), .CP(clk), .RN(n183), .Q(
        rd_data[2]) );
  HS65_LS_DFPRQX9 \rd_data_reg[1]  ( .D(N47), .CP(clk), .RN(n183), .Q(
        rd_data[1]) );
  HS65_LS_DFPRQX9 \rd_data_reg[0]  ( .D(N48), .CP(clk), .RN(n183), .Q(
        rd_data[0]) );
  HS65_LS_AND3X9 U3 ( .A(n191), .B(n190), .C(wr_ena), .Z(n1) );
  HS65_LS_BFX9 U4 ( .A(n165), .Z(n162) );
  HS65_LS_BFX9 U5 ( .A(n1), .Z(n168) );
  HS65_LS_BFX9 U6 ( .A(n155), .Z(n152) );
  HS65_LS_BFX9 U7 ( .A(n160), .Z(n157) );
  HS65_LS_AND2X4 U8 ( .A(rd_addr[1]), .B(rd_addr[0]), .Z(n321) );
  HS65_LS_AND2X4 U9 ( .A(rd_addr[1]), .B(n192), .Z(n322) );
  HS65_LS_BFX9 U10 ( .A(n185), .Z(n180) );
  HS65_LS_BFX9 U11 ( .A(n185), .Z(n179) );
  HS65_LS_BFX9 U12 ( .A(n185), .Z(n178) );
  HS65_LS_BFX9 U13 ( .A(n186), .Z(n177) );
  HS65_LS_BFX9 U14 ( .A(n186), .Z(n176) );
  HS65_LS_BFX9 U15 ( .A(n186), .Z(n175) );
  HS65_LS_BFX9 U16 ( .A(n187), .Z(n174) );
  HS65_LS_BFX9 U17 ( .A(n187), .Z(n173) );
  HS65_LS_BFX9 U18 ( .A(n187), .Z(n172) );
  HS65_LS_BFX9 U19 ( .A(n188), .Z(n185) );
  HS65_LS_BFX9 U20 ( .A(n188), .Z(n186) );
  HS65_LS_BFX9 U21 ( .A(n189), .Z(n187) );
  HS65_LS_BFX9 U22 ( .A(n184), .Z(n182) );
  HS65_LS_BFX9 U23 ( .A(n184), .Z(n181) );
  HS65_LS_BFX9 U24 ( .A(n188), .Z(n171) );
  HS65_LS_BFX9 U25 ( .A(n189), .Z(n188) );
  HS65_LS_BFX9 U26 ( .A(n184), .Z(n183) );
  HS65_LS_BFX9 U27 ( .A(n189), .Z(n184) );
  HS65_LS_IVX9 U28 ( .A(reset), .Z(n189) );
  HS65_LS_IVX9 U29 ( .A(n168), .Z(n167) );
  HS65_LS_IVX9 U30 ( .A(n168), .Z(n166) );
  HS65_LS_IVX9 U31 ( .A(n162), .Z(n161) );
  HS65_LS_BFX9 U32 ( .A(n1), .Z(n169) );
  HS65_LS_BFX9 U33 ( .A(n165), .Z(n163) );
  HS65_LS_BFX9 U34 ( .A(n1), .Z(n170) );
  HS65_LS_BFX9 U35 ( .A(n162), .Z(n164) );
  HS65_LS_IVX9 U36 ( .A(n157), .Z(n156) );
  HS65_LS_IVX9 U37 ( .A(n152), .Z(n151) );
  HS65_LS_BFX9 U38 ( .A(n160), .Z(n158) );
  HS65_LS_BFX9 U39 ( .A(n155), .Z(n153) );
  HS65_LS_BFX9 U40 ( .A(n157), .Z(n159) );
  HS65_LS_BFX9 U41 ( .A(n152), .Z(n154) );
  HS65_LS_IVX9 U42 ( .A(n327), .Z(n165) );
  HS65_LS_IVX9 U43 ( .A(wr_addr[0]), .Z(n191) );
  HS65_LS_NAND3X5 U44 ( .A(wr_ena), .B(n190), .C(wr_addr[0]), .Z(n327) );
  HS65_LS_BFX9 U45 ( .A(n322), .Z(n6) );
  HS65_LS_BFX9 U46 ( .A(n322), .Z(n5) );
  HS65_LS_BFX9 U47 ( .A(n321), .Z(n3) );
  HS65_LS_BFX9 U48 ( .A(n321), .Z(n2) );
  HS65_LS_BFX9 U49 ( .A(n8), .Z(n145) );
  HS65_LS_BFX9 U50 ( .A(n8), .Z(n9) );
  HS65_LS_BFX9 U51 ( .A(n147), .Z(n149) );
  HS65_LS_BFX9 U52 ( .A(n147), .Z(n148) );
  HS65_LS_BFX9 U53 ( .A(n321), .Z(n4) );
  HS65_LS_BFX9 U54 ( .A(n322), .Z(n7) );
  HS65_LS_BFX9 U55 ( .A(n8), .Z(n146) );
  HS65_LS_BFX9 U56 ( .A(n147), .Z(n150) );
  HS65_LS_IVX9 U57 ( .A(n326), .Z(n160) );
  HS65_LS_IVX9 U58 ( .A(n325), .Z(n155) );
  HS65_LS_IVX9 U59 ( .A(wr_addr[1]), .Z(n190) );
  HS65_LS_NAND3X5 U60 ( .A(wr_addr[0]), .B(wr_ena), .C(wr_addr[1]), .Z(n325)
         );
  HS65_LS_NAND3X5 U61 ( .A(wr_ena), .B(n191), .C(wr_addr[1]), .Z(n326) );
  HS65_LS_BFX9 U62 ( .A(n324), .Z(n147) );
  HS65_LS_NOR2X6 U63 ( .A(rd_addr[0]), .B(rd_addr[1]), .Z(n324) );
  HS65_LS_BFX9 U64 ( .A(n323), .Z(n8) );
  HS65_LS_NOR2X6 U65 ( .A(n192), .B(rd_addr[1]), .Z(n323) );
  HS65_LS_IVX9 U66 ( .A(rd_addr[0]), .Z(n192) );
  HS65_LS_MX41X7 U67 ( .D0(n150), .S0(\mem[0][0] ), .D1(n146), .S1(\mem[1][0] ), .D2(n7), .S2(\mem[2][0] ), .D3(n4), .S3(\mem[3][0] ), .Z(N48) );
  HS65_LS_MX41X7 U68 ( .D0(n150), .S0(\mem[0][1] ), .D1(n146), .S1(\mem[1][1] ), .D2(n7), .S2(\mem[2][1] ), .D3(n4), .S3(\mem[3][1] ), .Z(N47) );
  HS65_LS_MX41X7 U69 ( .D0(n150), .S0(\mem[0][2] ), .D1(n146), .S1(\mem[1][2] ), .D2(n7), .S2(\mem[2][2] ), .D3(n4), .S3(\mem[3][2] ), .Z(N46) );
  HS65_LS_MX41X7 U70 ( .D0(n150), .S0(\mem[0][3] ), .D1(n146), .S1(\mem[1][3] ), .D2(n7), .S2(\mem[2][3] ), .D3(n4), .S3(\mem[3][3] ), .Z(N45) );
  HS65_LS_MX41X7 U71 ( .D0(n150), .S0(\mem[0][4] ), .D1(n146), .S1(\mem[1][4] ), .D2(n7), .S2(\mem[2][4] ), .D3(n4), .S3(\mem[3][4] ), .Z(N44) );
  HS65_LS_MX41X7 U72 ( .D0(n150), .S0(\mem[0][5] ), .D1(n146), .S1(\mem[1][5] ), .D2(n7), .S2(\mem[2][5] ), .D3(n4), .S3(\mem[3][5] ), .Z(N43) );
  HS65_LS_MX41X7 U73 ( .D0(n150), .S0(\mem[0][6] ), .D1(n146), .S1(\mem[1][6] ), .D2(n6), .S2(\mem[2][6] ), .D3(n4), .S3(\mem[3][6] ), .Z(N42) );
  HS65_LS_MX41X7 U74 ( .D0(n150), .S0(\mem[0][7] ), .D1(n146), .S1(\mem[1][7] ), .D2(n6), .S2(\mem[2][7] ), .D3(n4), .S3(\mem[3][7] ), .Z(N41) );
  HS65_LS_MX41X7 U75 ( .D0(n149), .S0(\mem[0][8] ), .D1(n145), .S1(\mem[1][8] ), .D2(n6), .S2(\mem[2][8] ), .D3(n3), .S3(\mem[3][8] ), .Z(N40) );
  HS65_LS_MX41X7 U76 ( .D0(n149), .S0(\mem[0][9] ), .D1(n145), .S1(\mem[1][9] ), .D2(n6), .S2(\mem[2][9] ), .D3(n3), .S3(\mem[3][9] ), .Z(N39) );
  HS65_LS_MX41X7 U77 ( .D0(n149), .S0(\mem[0][10] ), .D1(n145), .S1(
        \mem[1][10] ), .D2(n6), .S2(\mem[2][10] ), .D3(n3), .S3(\mem[3][10] ), 
        .Z(N38) );
  HS65_LS_MX41X7 U78 ( .D0(n149), .S0(\mem[0][11] ), .D1(n145), .S1(
        \mem[1][11] ), .D2(n6), .S2(\mem[2][11] ), .D3(n3), .S3(\mem[3][11] ), 
        .Z(N37) );
  HS65_LS_MX41X7 U79 ( .D0(n149), .S0(\mem[0][12] ), .D1(n145), .S1(
        \mem[1][12] ), .D2(n6), .S2(\mem[2][12] ), .D3(n3), .S3(\mem[3][12] ), 
        .Z(N36) );
  HS65_LS_MX41X7 U80 ( .D0(n149), .S0(\mem[0][13] ), .D1(n145), .S1(
        \mem[1][13] ), .D2(n6), .S2(\mem[2][13] ), .D3(n3), .S3(\mem[3][13] ), 
        .Z(N35) );
  HS65_LS_MX41X7 U81 ( .D0(n149), .S0(\mem[0][14] ), .D1(n145), .S1(
        \mem[1][14] ), .D2(n6), .S2(\mem[2][14] ), .D3(n3), .S3(\mem[3][14] ), 
        .Z(N34) );
  HS65_LS_MX41X7 U82 ( .D0(n149), .S0(\mem[0][15] ), .D1(n145), .S1(
        \mem[1][15] ), .D2(n6), .S2(\mem[2][15] ), .D3(n3), .S3(\mem[3][15] ), 
        .Z(N33) );
  HS65_LS_MX41X7 U83 ( .D0(n149), .S0(\mem[0][16] ), .D1(n145), .S1(
        \mem[1][16] ), .D2(n6), .S2(\mem[2][16] ), .D3(n3), .S3(\mem[3][16] ), 
        .Z(N32) );
  HS65_LS_MX41X7 U84 ( .D0(n149), .S0(\mem[0][17] ), .D1(n145), .S1(
        \mem[1][17] ), .D2(n6), .S2(\mem[2][17] ), .D3(n3), .S3(\mem[3][17] ), 
        .Z(N31) );
  HS65_LS_MX41X7 U85 ( .D0(n149), .S0(\mem[0][18] ), .D1(n145), .S1(
        \mem[1][18] ), .D2(n6), .S2(\mem[2][18] ), .D3(n3), .S3(\mem[3][18] ), 
        .Z(N30) );
  HS65_LS_MX41X7 U86 ( .D0(n149), .S0(\mem[0][19] ), .D1(n145), .S1(
        \mem[1][19] ), .D2(n5), .S2(\mem[2][19] ), .D3(n3), .S3(\mem[3][19] ), 
        .Z(N29) );
  HS65_LS_MX41X7 U87 ( .D0(n148), .S0(\mem[0][20] ), .D1(n9), .S1(\mem[1][20] ), .D2(n5), .S2(\mem[2][20] ), .D3(n2), .S3(\mem[3][20] ), .Z(N28) );
  HS65_LS_MX41X7 U88 ( .D0(n148), .S0(\mem[0][21] ), .D1(n9), .S1(\mem[1][21] ), .D2(n5), .S2(\mem[2][21] ), .D3(n2), .S3(\mem[3][21] ), .Z(N27) );
  HS65_LS_MX41X7 U89 ( .D0(n148), .S0(\mem[0][22] ), .D1(n9), .S1(\mem[1][22] ), .D2(n5), .S2(\mem[2][22] ), .D3(n2), .S3(\mem[3][22] ), .Z(N26) );
  HS65_LS_MX41X7 U90 ( .D0(n148), .S0(\mem[0][23] ), .D1(n9), .S1(\mem[1][23] ), .D2(n5), .S2(\mem[2][23] ), .D3(n2), .S3(\mem[3][23] ), .Z(N25) );
  HS65_LS_MX41X7 U91 ( .D0(n148), .S0(\mem[0][24] ), .D1(n9), .S1(\mem[1][24] ), .D2(n5), .S2(\mem[2][24] ), .D3(n2), .S3(\mem[3][24] ), .Z(N24) );
  HS65_LS_MX41X7 U92 ( .D0(n148), .S0(\mem[0][25] ), .D1(n9), .S1(\mem[1][25] ), .D2(n5), .S2(\mem[2][25] ), .D3(n2), .S3(\mem[3][25] ), .Z(N23) );
  HS65_LS_MX41X7 U93 ( .D0(n148), .S0(\mem[0][26] ), .D1(n9), .S1(\mem[1][26] ), .D2(n5), .S2(\mem[2][26] ), .D3(n2), .S3(\mem[3][26] ), .Z(N22) );
  HS65_LS_MX41X7 U94 ( .D0(n148), .S0(\mem[0][27] ), .D1(n9), .S1(\mem[1][27] ), .D2(n5), .S2(\mem[2][27] ), .D3(n2), .S3(\mem[3][27] ), .Z(N21) );
  HS65_LS_MX41X7 U95 ( .D0(n148), .S0(\mem[0][28] ), .D1(n9), .S1(\mem[1][28] ), .D2(n5), .S2(\mem[2][28] ), .D3(n2), .S3(\mem[3][28] ), .Z(N20) );
  HS65_LS_MX41X7 U96 ( .D0(n148), .S0(\mem[0][29] ), .D1(n9), .S1(\mem[1][29] ), .D2(n5), .S2(\mem[2][29] ), .D3(n2), .S3(\mem[3][29] ), .Z(N19) );
  HS65_LS_MX41X7 U97 ( .D0(n148), .S0(\mem[0][30] ), .D1(n9), .S1(\mem[1][30] ), .D2(n5), .S2(\mem[2][30] ), .D3(n2), .S3(\mem[3][30] ), .Z(N18) );
  HS65_LS_MX41X7 U98 ( .D0(n148), .S0(\mem[0][31] ), .D1(n9), .S1(\mem[1][31] ), .D2(n5), .S2(\mem[2][31] ), .D3(n2), .S3(\mem[3][31] ), .Z(N17) );
  HS65_LS_AO22X9 U99 ( .A(wr_data[0]), .B(n154), .C(n151), .D(\mem[3][0] ), 
        .Z(n224) );
  HS65_LS_AO22X9 U100 ( .A(wr_data[1]), .B(n154), .C(n151), .D(\mem[3][1] ), 
        .Z(n223) );
  HS65_LS_AO22X9 U101 ( .A(wr_data[2]), .B(n154), .C(n151), .D(\mem[3][2] ), 
        .Z(n222) );
  HS65_LS_AO22X9 U102 ( .A(wr_data[3]), .B(n154), .C(n151), .D(\mem[3][3] ), 
        .Z(n221) );
  HS65_LS_AO22X9 U103 ( .A(wr_data[4]), .B(n154), .C(n151), .D(\mem[3][4] ), 
        .Z(n220) );
  HS65_LS_AO22X9 U104 ( .A(wr_data[5]), .B(n154), .C(n151), .D(\mem[3][5] ), 
        .Z(n219) );
  HS65_LS_AO22X9 U105 ( .A(wr_data[6]), .B(n154), .C(n151), .D(\mem[3][6] ), 
        .Z(n218) );
  HS65_LS_AO22X9 U106 ( .A(wr_data[7]), .B(n154), .C(n151), .D(\mem[3][7] ), 
        .Z(n217) );
  HS65_LS_AO22X9 U107 ( .A(wr_data[8]), .B(n154), .C(n151), .D(\mem[3][8] ), 
        .Z(n216) );
  HS65_LS_AO22X9 U108 ( .A(wr_data[9]), .B(n154), .C(n151), .D(\mem[3][9] ), 
        .Z(n215) );
  HS65_LS_AO22X9 U109 ( .A(wr_data[10]), .B(n154), .C(n151), .D(\mem[3][10] ), 
        .Z(n214) );
  HS65_LS_AO22X9 U110 ( .A(wr_data[11]), .B(n153), .C(n151), .D(\mem[3][11] ), 
        .Z(n213) );
  HS65_LS_AO22X9 U111 ( .A(wr_data[12]), .B(n153), .C(n151), .D(\mem[3][12] ), 
        .Z(n212) );
  HS65_LS_AO22X9 U112 ( .A(wr_data[13]), .B(n153), .C(n151), .D(\mem[3][13] ), 
        .Z(n211) );
  HS65_LS_AO22X9 U113 ( .A(wr_data[14]), .B(n153), .C(n151), .D(\mem[3][14] ), 
        .Z(n210) );
  HS65_LS_AO22X9 U114 ( .A(wr_data[15]), .B(n153), .C(n151), .D(\mem[3][15] ), 
        .Z(n209) );
  HS65_LS_AO22X9 U115 ( .A(wr_data[16]), .B(n153), .C(n151), .D(\mem[3][16] ), 
        .Z(n208) );
  HS65_LS_AO22X9 U116 ( .A(wr_data[17]), .B(n153), .C(n151), .D(\mem[3][17] ), 
        .Z(n207) );
  HS65_LS_AO22X9 U117 ( .A(wr_data[18]), .B(n153), .C(n151), .D(\mem[3][18] ), 
        .Z(n206) );
  HS65_LS_AO22X9 U118 ( .A(wr_data[19]), .B(n153), .C(n151), .D(\mem[3][19] ), 
        .Z(n205) );
  HS65_LS_AO22X9 U119 ( .A(wr_data[20]), .B(n153), .C(n325), .D(\mem[3][20] ), 
        .Z(n204) );
  HS65_LS_AO22X9 U120 ( .A(wr_data[21]), .B(n153), .C(n325), .D(\mem[3][21] ), 
        .Z(n203) );
  HS65_LS_AO22X9 U121 ( .A(wr_data[22]), .B(n153), .C(n325), .D(\mem[3][22] ), 
        .Z(n202) );
  HS65_LS_AO22X9 U122 ( .A(wr_data[23]), .B(n153), .C(n325), .D(\mem[3][23] ), 
        .Z(n201) );
  HS65_LS_AO22X9 U123 ( .A(wr_data[24]), .B(n153), .C(n325), .D(\mem[3][24] ), 
        .Z(n200) );
  HS65_LS_AO22X9 U124 ( .A(wr_data[25]), .B(n153), .C(n325), .D(\mem[3][25] ), 
        .Z(n199) );
  HS65_LS_AO22X9 U125 ( .A(wr_data[26]), .B(n153), .C(n325), .D(\mem[3][26] ), 
        .Z(n198) );
  HS65_LS_AO22X9 U126 ( .A(wr_data[27]), .B(n153), .C(n325), .D(\mem[3][27] ), 
        .Z(n197) );
  HS65_LS_AO22X9 U127 ( .A(wr_data[28]), .B(n153), .C(n325), .D(\mem[3][28] ), 
        .Z(n196) );
  HS65_LS_AO22X9 U128 ( .A(wr_data[29]), .B(n153), .C(n325), .D(\mem[3][29] ), 
        .Z(n195) );
  HS65_LS_AO22X9 U129 ( .A(wr_data[30]), .B(n153), .C(n325), .D(\mem[3][30] ), 
        .Z(n194) );
  HS65_LS_AO22X9 U130 ( .A(wr_data[31]), .B(n152), .C(n325), .D(\mem[3][31] ), 
        .Z(n193) );
  HS65_LS_AO22X9 U131 ( .A(wr_data[0]), .B(n164), .C(n161), .D(\mem[1][0] ), 
        .Z(n288) );
  HS65_LS_AO22X9 U132 ( .A(wr_data[1]), .B(n164), .C(n161), .D(\mem[1][1] ), 
        .Z(n287) );
  HS65_LS_AO22X9 U133 ( .A(wr_data[2]), .B(n164), .C(n161), .D(\mem[1][2] ), 
        .Z(n286) );
  HS65_LS_AO22X9 U134 ( .A(wr_data[3]), .B(n164), .C(n161), .D(\mem[1][3] ), 
        .Z(n285) );
  HS65_LS_AO22X9 U135 ( .A(wr_data[4]), .B(n164), .C(n161), .D(\mem[1][4] ), 
        .Z(n284) );
  HS65_LS_AO22X9 U136 ( .A(wr_data[5]), .B(n164), .C(n161), .D(\mem[1][5] ), 
        .Z(n283) );
  HS65_LS_AO22X9 U137 ( .A(wr_data[6]), .B(n164), .C(n161), .D(\mem[1][6] ), 
        .Z(n282) );
  HS65_LS_AO22X9 U138 ( .A(wr_data[7]), .B(n164), .C(n161), .D(\mem[1][7] ), 
        .Z(n281) );
  HS65_LS_AO22X9 U139 ( .A(wr_data[8]), .B(n164), .C(n161), .D(\mem[1][8] ), 
        .Z(n280) );
  HS65_LS_AO22X9 U140 ( .A(wr_data[9]), .B(n164), .C(n161), .D(\mem[1][9] ), 
        .Z(n279) );
  HS65_LS_AO22X9 U141 ( .A(wr_data[10]), .B(n164), .C(n161), .D(\mem[1][10] ), 
        .Z(n278) );
  HS65_LS_AO22X9 U142 ( .A(wr_data[11]), .B(n163), .C(n161), .D(\mem[1][11] ), 
        .Z(n277) );
  HS65_LS_AO22X9 U143 ( .A(wr_data[12]), .B(n163), .C(n161), .D(\mem[1][12] ), 
        .Z(n276) );
  HS65_LS_AO22X9 U144 ( .A(wr_data[13]), .B(n163), .C(n161), .D(\mem[1][13] ), 
        .Z(n275) );
  HS65_LS_AO22X9 U145 ( .A(wr_data[14]), .B(n163), .C(n161), .D(\mem[1][14] ), 
        .Z(n274) );
  HS65_LS_AO22X9 U146 ( .A(wr_data[15]), .B(n163), .C(n161), .D(\mem[1][15] ), 
        .Z(n273) );
  HS65_LS_AO22X9 U147 ( .A(wr_data[16]), .B(n163), .C(n161), .D(\mem[1][16] ), 
        .Z(n272) );
  HS65_LS_AO22X9 U148 ( .A(wr_data[17]), .B(n163), .C(n161), .D(\mem[1][17] ), 
        .Z(n271) );
  HS65_LS_AO22X9 U149 ( .A(wr_data[18]), .B(n163), .C(n161), .D(\mem[1][18] ), 
        .Z(n270) );
  HS65_LS_AO22X9 U150 ( .A(wr_data[19]), .B(n163), .C(n161), .D(\mem[1][19] ), 
        .Z(n269) );
  HS65_LS_AO22X9 U151 ( .A(wr_data[20]), .B(n163), .C(n327), .D(\mem[1][20] ), 
        .Z(n268) );
  HS65_LS_AO22X9 U152 ( .A(wr_data[21]), .B(n163), .C(n327), .D(\mem[1][21] ), 
        .Z(n267) );
  HS65_LS_AO22X9 U153 ( .A(wr_data[22]), .B(n163), .C(n327), .D(\mem[1][22] ), 
        .Z(n266) );
  HS65_LS_AO22X9 U154 ( .A(wr_data[23]), .B(n163), .C(n327), .D(\mem[1][23] ), 
        .Z(n265) );
  HS65_LS_AO22X9 U155 ( .A(wr_data[24]), .B(n163), .C(n327), .D(\mem[1][24] ), 
        .Z(n264) );
  HS65_LS_AO22X9 U156 ( .A(wr_data[25]), .B(n163), .C(n327), .D(\mem[1][25] ), 
        .Z(n263) );
  HS65_LS_AO22X9 U157 ( .A(wr_data[26]), .B(n163), .C(n327), .D(\mem[1][26] ), 
        .Z(n262) );
  HS65_LS_AO22X9 U158 ( .A(wr_data[27]), .B(n163), .C(n327), .D(\mem[1][27] ), 
        .Z(n261) );
  HS65_LS_AO22X9 U159 ( .A(wr_data[28]), .B(n163), .C(n327), .D(\mem[1][28] ), 
        .Z(n260) );
  HS65_LS_AO22X9 U160 ( .A(wr_data[29]), .B(n163), .C(n327), .D(\mem[1][29] ), 
        .Z(n259) );
  HS65_LS_AO22X9 U161 ( .A(wr_data[30]), .B(n163), .C(n327), .D(\mem[1][30] ), 
        .Z(n258) );
  HS65_LS_AO22X9 U162 ( .A(wr_data[31]), .B(n162), .C(n327), .D(\mem[1][31] ), 
        .Z(n257) );
  HS65_LS_AO22X9 U163 ( .A(n170), .B(wr_data[0]), .C(n167), .D(\mem[0][0] ), 
        .Z(n320) );
  HS65_LS_AO22X9 U164 ( .A(n170), .B(wr_data[1]), .C(n166), .D(\mem[0][1] ), 
        .Z(n319) );
  HS65_LS_AO22X9 U165 ( .A(n170), .B(wr_data[2]), .C(n167), .D(\mem[0][2] ), 
        .Z(n318) );
  HS65_LS_AO22X9 U166 ( .A(n170), .B(wr_data[3]), .C(n166), .D(\mem[0][3] ), 
        .Z(n317) );
  HS65_LS_AO22X9 U167 ( .A(n170), .B(wr_data[4]), .C(n167), .D(\mem[0][4] ), 
        .Z(n316) );
  HS65_LS_AO22X9 U168 ( .A(n170), .B(wr_data[5]), .C(n166), .D(\mem[0][5] ), 
        .Z(n315) );
  HS65_LS_AO22X9 U169 ( .A(n170), .B(wr_data[6]), .C(n167), .D(\mem[0][6] ), 
        .Z(n314) );
  HS65_LS_AO22X9 U170 ( .A(n170), .B(wr_data[7]), .C(n167), .D(\mem[0][7] ), 
        .Z(n313) );
  HS65_LS_AO22X9 U171 ( .A(n170), .B(wr_data[8]), .C(n167), .D(\mem[0][8] ), 
        .Z(n312) );
  HS65_LS_AO22X9 U172 ( .A(n170), .B(wr_data[9]), .C(n167), .D(\mem[0][9] ), 
        .Z(n311) );
  HS65_LS_AO22X9 U173 ( .A(n170), .B(wr_data[10]), .C(n167), .D(\mem[0][10] ), 
        .Z(n310) );
  HS65_LS_AO22X9 U174 ( .A(n169), .B(wr_data[11]), .C(n167), .D(\mem[0][11] ), 
        .Z(n309) );
  HS65_LS_AO22X9 U175 ( .A(n169), .B(wr_data[12]), .C(n167), .D(\mem[0][12] ), 
        .Z(n308) );
  HS65_LS_AO22X9 U176 ( .A(n169), .B(wr_data[13]), .C(n167), .D(\mem[0][13] ), 
        .Z(n307) );
  HS65_LS_AO22X9 U177 ( .A(n169), .B(wr_data[14]), .C(n167), .D(\mem[0][14] ), 
        .Z(n306) );
  HS65_LS_AO22X9 U178 ( .A(n169), .B(wr_data[15]), .C(n167), .D(\mem[0][15] ), 
        .Z(n305) );
  HS65_LS_AO22X9 U179 ( .A(n169), .B(wr_data[16]), .C(n167), .D(\mem[0][16] ), 
        .Z(n304) );
  HS65_LS_AO22X9 U180 ( .A(n169), .B(wr_data[17]), .C(n167), .D(\mem[0][17] ), 
        .Z(n303) );
  HS65_LS_AO22X9 U181 ( .A(n169), .B(wr_data[18]), .C(n167), .D(\mem[0][18] ), 
        .Z(n302) );
  HS65_LS_AO22X9 U182 ( .A(n169), .B(wr_data[19]), .C(n166), .D(\mem[0][19] ), 
        .Z(n301) );
  HS65_LS_AO22X9 U183 ( .A(n169), .B(wr_data[20]), .C(n166), .D(\mem[0][20] ), 
        .Z(n300) );
  HS65_LS_AO22X9 U184 ( .A(n169), .B(wr_data[21]), .C(n166), .D(\mem[0][21] ), 
        .Z(n299) );
  HS65_LS_AO22X9 U185 ( .A(n169), .B(wr_data[22]), .C(n166), .D(\mem[0][22] ), 
        .Z(n298) );
  HS65_LS_AO22X9 U186 ( .A(n169), .B(wr_data[23]), .C(n166), .D(\mem[0][23] ), 
        .Z(n297) );
  HS65_LS_AO22X9 U187 ( .A(n169), .B(wr_data[24]), .C(n166), .D(\mem[0][24] ), 
        .Z(n296) );
  HS65_LS_AO22X9 U188 ( .A(n169), .B(wr_data[25]), .C(n166), .D(\mem[0][25] ), 
        .Z(n295) );
  HS65_LS_AO22X9 U189 ( .A(n169), .B(wr_data[26]), .C(n166), .D(\mem[0][26] ), 
        .Z(n294) );
  HS65_LS_AO22X9 U190 ( .A(n169), .B(wr_data[27]), .C(n166), .D(\mem[0][27] ), 
        .Z(n293) );
  HS65_LS_AO22X9 U191 ( .A(n169), .B(wr_data[28]), .C(n166), .D(\mem[0][28] ), 
        .Z(n292) );
  HS65_LS_AO22X9 U192 ( .A(n169), .B(wr_data[29]), .C(n166), .D(\mem[0][29] ), 
        .Z(n291) );
  HS65_LS_AO22X9 U193 ( .A(n169), .B(wr_data[30]), .C(n166), .D(\mem[0][30] ), 
        .Z(n290) );
  HS65_LS_AO22X9 U194 ( .A(n168), .B(wr_data[31]), .C(n166), .D(\mem[0][31] ), 
        .Z(n289) );
  HS65_LS_AO22X9 U195 ( .A(wr_data[0]), .B(n159), .C(n156), .D(\mem[2][0] ), 
        .Z(n256) );
  HS65_LS_AO22X9 U196 ( .A(wr_data[1]), .B(n159), .C(n156), .D(\mem[2][1] ), 
        .Z(n255) );
  HS65_LS_AO22X9 U197 ( .A(wr_data[2]), .B(n159), .C(n156), .D(\mem[2][2] ), 
        .Z(n254) );
  HS65_LS_AO22X9 U198 ( .A(wr_data[3]), .B(n159), .C(n156), .D(\mem[2][3] ), 
        .Z(n253) );
  HS65_LS_AO22X9 U199 ( .A(wr_data[4]), .B(n159), .C(n156), .D(\mem[2][4] ), 
        .Z(n252) );
  HS65_LS_AO22X9 U200 ( .A(wr_data[5]), .B(n159), .C(n156), .D(\mem[2][5] ), 
        .Z(n251) );
  HS65_LS_AO22X9 U201 ( .A(wr_data[6]), .B(n159), .C(n156), .D(\mem[2][6] ), 
        .Z(n250) );
  HS65_LS_AO22X9 U202 ( .A(wr_data[7]), .B(n159), .C(n156), .D(\mem[2][7] ), 
        .Z(n249) );
  HS65_LS_AO22X9 U203 ( .A(wr_data[8]), .B(n159), .C(n156), .D(\mem[2][8] ), 
        .Z(n248) );
  HS65_LS_AO22X9 U204 ( .A(wr_data[9]), .B(n159), .C(n156), .D(\mem[2][9] ), 
        .Z(n247) );
  HS65_LS_AO22X9 U205 ( .A(wr_data[10]), .B(n159), .C(n156), .D(\mem[2][10] ), 
        .Z(n246) );
  HS65_LS_AO22X9 U206 ( .A(wr_data[11]), .B(n158), .C(n156), .D(\mem[2][11] ), 
        .Z(n245) );
  HS65_LS_AO22X9 U207 ( .A(wr_data[12]), .B(n158), .C(n156), .D(\mem[2][12] ), 
        .Z(n244) );
  HS65_LS_AO22X9 U208 ( .A(wr_data[13]), .B(n158), .C(n156), .D(\mem[2][13] ), 
        .Z(n243) );
  HS65_LS_AO22X9 U209 ( .A(wr_data[14]), .B(n158), .C(n156), .D(\mem[2][14] ), 
        .Z(n242) );
  HS65_LS_AO22X9 U210 ( .A(wr_data[15]), .B(n158), .C(n156), .D(\mem[2][15] ), 
        .Z(n241) );
  HS65_LS_AO22X9 U211 ( .A(wr_data[16]), .B(n158), .C(n156), .D(\mem[2][16] ), 
        .Z(n240) );
  HS65_LS_AO22X9 U212 ( .A(wr_data[17]), .B(n158), .C(n156), .D(\mem[2][17] ), 
        .Z(n239) );
  HS65_LS_AO22X9 U213 ( .A(wr_data[18]), .B(n158), .C(n156), .D(\mem[2][18] ), 
        .Z(n238) );
  HS65_LS_AO22X9 U214 ( .A(wr_data[19]), .B(n158), .C(n156), .D(\mem[2][19] ), 
        .Z(n237) );
  HS65_LS_AO22X9 U215 ( .A(wr_data[20]), .B(n158), .C(n326), .D(\mem[2][20] ), 
        .Z(n236) );
  HS65_LS_AO22X9 U216 ( .A(wr_data[21]), .B(n158), .C(n326), .D(\mem[2][21] ), 
        .Z(n235) );
  HS65_LS_AO22X9 U217 ( .A(wr_data[22]), .B(n158), .C(n326), .D(\mem[2][22] ), 
        .Z(n234) );
  HS65_LS_AO22X9 U218 ( .A(wr_data[23]), .B(n158), .C(n326), .D(\mem[2][23] ), 
        .Z(n233) );
  HS65_LS_AO22X9 U219 ( .A(wr_data[24]), .B(n158), .C(n326), .D(\mem[2][24] ), 
        .Z(n232) );
  HS65_LS_AO22X9 U220 ( .A(wr_data[25]), .B(n158), .C(n326), .D(\mem[2][25] ), 
        .Z(n231) );
  HS65_LS_AO22X9 U221 ( .A(wr_data[26]), .B(n158), .C(n326), .D(\mem[2][26] ), 
        .Z(n230) );
  HS65_LS_AO22X9 U222 ( .A(wr_data[27]), .B(n158), .C(n326), .D(\mem[2][27] ), 
        .Z(n229) );
  HS65_LS_AO22X9 U223 ( .A(wr_data[28]), .B(n158), .C(n326), .D(\mem[2][28] ), 
        .Z(n228) );
  HS65_LS_AO22X9 U224 ( .A(wr_data[29]), .B(n158), .C(n326), .D(\mem[2][29] ), 
        .Z(n227) );
  HS65_LS_AO22X9 U225 ( .A(wr_data[30]), .B(n158), .C(n326), .D(\mem[2][30] ), 
        .Z(n226) );
  HS65_LS_AO22X9 U226 ( .A(wr_data[31]), .B(n157), .C(n326), .D(\mem[2][31] ), 
        .Z(n225) );
endmodule


module bram_DATA16_ADDR2_3 ( clk, reset, rd_addr, wr_addr, wr_data, wr_ena, 
        rd_data );
  input [1:0] rd_addr;
  input [1:0] wr_addr;
  input [15:0] wr_data;
  output [15:0] rd_data;
  input clk, reset, wr_ena;
  wire   \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] ,
         \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][15] , \mem[1][14] , \mem[1][13] ,
         \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] , \mem[1][8] ,
         \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] ,
         \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][15] , \mem[0][14] ,
         \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] ,
         \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] ,
         \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, n1,
         n2, n3, n4, n5, n6, n7, n8, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162;

  HS65_LS_DFPRQX9 \mem_reg[3][15]  ( .D(n91), .CP(clk), .RN(n1), .Q(
        \mem[3][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][14]  ( .D(n92), .CP(clk), .RN(n1), .Q(
        \mem[3][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][13]  ( .D(n93), .CP(clk), .RN(n1), .Q(
        \mem[3][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][12]  ( .D(n94), .CP(clk), .RN(n1), .Q(
        \mem[3][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][11]  ( .D(n95), .CP(clk), .RN(n1), .Q(
        \mem[3][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][10]  ( .D(n96), .CP(clk), .RN(n1), .Q(
        \mem[3][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][9]  ( .D(n97), .CP(clk), .RN(n1), .Q(\mem[3][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][8]  ( .D(n98), .CP(clk), .RN(n1), .Q(\mem[3][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][7]  ( .D(n99), .CP(clk), .RN(n1), .Q(\mem[3][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][6]  ( .D(n100), .CP(clk), .RN(n1), .Q(
        \mem[3][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][5]  ( .D(n101), .CP(clk), .RN(n1), .Q(
        \mem[3][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][4]  ( .D(n102), .CP(clk), .RN(n1), .Q(
        \mem[3][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][3]  ( .D(n103), .CP(clk), .RN(n1), .Q(
        \mem[3][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][2]  ( .D(n104), .CP(clk), .RN(n2), .Q(
        \mem[3][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][1]  ( .D(n105), .CP(clk), .RN(n2), .Q(
        \mem[3][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][0]  ( .D(n106), .CP(clk), .RN(n2), .Q(
        \mem[3][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][15]  ( .D(n107), .CP(clk), .RN(n2), .Q(
        \mem[2][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][14]  ( .D(n108), .CP(clk), .RN(n2), .Q(
        \mem[2][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][13]  ( .D(n109), .CP(clk), .RN(n2), .Q(
        \mem[2][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][12]  ( .D(n110), .CP(clk), .RN(n2), .Q(
        \mem[2][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][11]  ( .D(n111), .CP(clk), .RN(n2), .Q(
        \mem[2][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][10]  ( .D(n112), .CP(clk), .RN(n2), .Q(
        \mem[2][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][9]  ( .D(n113), .CP(clk), .RN(n2), .Q(
        \mem[2][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][8]  ( .D(n114), .CP(clk), .RN(n2), .Q(
        \mem[2][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][7]  ( .D(n115), .CP(clk), .RN(n2), .Q(
        \mem[2][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][6]  ( .D(n116), .CP(clk), .RN(n2), .Q(
        \mem[2][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][5]  ( .D(n117), .CP(clk), .RN(n3), .Q(
        \mem[2][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][4]  ( .D(n118), .CP(clk), .RN(n3), .Q(
        \mem[2][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][3]  ( .D(n119), .CP(clk), .RN(n3), .Q(
        \mem[2][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][2]  ( .D(n120), .CP(clk), .RN(n3), .Q(
        \mem[2][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][1]  ( .D(n121), .CP(clk), .RN(n3), .Q(
        \mem[2][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][0]  ( .D(n122), .CP(clk), .RN(n3), .Q(
        \mem[2][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][15]  ( .D(n123), .CP(clk), .RN(n3), .Q(
        \mem[1][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][14]  ( .D(n124), .CP(clk), .RN(n3), .Q(
        \mem[1][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][13]  ( .D(n125), .CP(clk), .RN(n3), .Q(
        \mem[1][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][12]  ( .D(n126), .CP(clk), .RN(n3), .Q(
        \mem[1][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][11]  ( .D(n127), .CP(clk), .RN(n3), .Q(
        \mem[1][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][10]  ( .D(n128), .CP(clk), .RN(n3), .Q(
        \mem[1][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][9]  ( .D(n129), .CP(clk), .RN(n3), .Q(
        \mem[1][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][8]  ( .D(n130), .CP(clk), .RN(n4), .Q(
        \mem[1][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][7]  ( .D(n131), .CP(clk), .RN(n4), .Q(
        \mem[1][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][6]  ( .D(n132), .CP(clk), .RN(n4), .Q(
        \mem[1][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][5]  ( .D(n133), .CP(clk), .RN(n4), .Q(
        \mem[1][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][4]  ( .D(n134), .CP(clk), .RN(n4), .Q(
        \mem[1][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][3]  ( .D(n135), .CP(clk), .RN(n4), .Q(
        \mem[1][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][2]  ( .D(n136), .CP(clk), .RN(n4), .Q(
        \mem[1][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][1]  ( .D(n137), .CP(clk), .RN(n4), .Q(
        \mem[1][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][0]  ( .D(n138), .CP(clk), .RN(n4), .Q(
        \mem[1][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][15]  ( .D(n139), .CP(clk), .RN(n4), .Q(
        \mem[0][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][14]  ( .D(n140), .CP(clk), .RN(n4), .Q(
        \mem[0][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][13]  ( .D(n141), .CP(clk), .RN(n4), .Q(
        \mem[0][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][12]  ( .D(n142), .CP(clk), .RN(n4), .Q(
        \mem[0][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][11]  ( .D(n143), .CP(clk), .RN(n5), .Q(
        \mem[0][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][10]  ( .D(n144), .CP(clk), .RN(n5), .Q(
        \mem[0][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][9]  ( .D(n145), .CP(clk), .RN(n5), .Q(
        \mem[0][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][8]  ( .D(n146), .CP(clk), .RN(n5), .Q(
        \mem[0][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][7]  ( .D(n147), .CP(clk), .RN(n5), .Q(
        \mem[0][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][6]  ( .D(n148), .CP(clk), .RN(n5), .Q(
        \mem[0][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][5]  ( .D(n149), .CP(clk), .RN(n5), .Q(
        \mem[0][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][4]  ( .D(n150), .CP(clk), .RN(n5), .Q(
        \mem[0][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][3]  ( .D(n151), .CP(clk), .RN(n5), .Q(
        \mem[0][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][2]  ( .D(n152), .CP(clk), .RN(n5), .Q(
        \mem[0][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][1]  ( .D(n153), .CP(clk), .RN(n5), .Q(
        \mem[0][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][0]  ( .D(n154), .CP(clk), .RN(n5), .Q(
        \mem[0][0] ) );
  HS65_LS_DFPRQX9 \rd_data_reg[15]  ( .D(N17), .CP(clk), .RN(n5), .Q(
        rd_data[15]) );
  HS65_LS_DFPRQX9 \rd_data_reg[14]  ( .D(N18), .CP(clk), .RN(n6), .Q(
        rd_data[14]) );
  HS65_LS_DFPRQX9 \rd_data_reg[13]  ( .D(N19), .CP(clk), .RN(n6), .Q(
        rd_data[13]) );
  HS65_LS_DFPRQX9 \rd_data_reg[12]  ( .D(N20), .CP(clk), .RN(n6), .Q(
        rd_data[12]) );
  HS65_LS_DFPRQX9 \rd_data_reg[11]  ( .D(N21), .CP(clk), .RN(n6), .Q(
        rd_data[11]) );
  HS65_LS_DFPRQX9 \rd_data_reg[10]  ( .D(N22), .CP(clk), .RN(n6), .Q(
        rd_data[10]) );
  HS65_LS_DFPRQX9 \rd_data_reg[9]  ( .D(N23), .CP(clk), .RN(n6), .Q(rd_data[9]) );
  HS65_LS_DFPRQX9 \rd_data_reg[8]  ( .D(N24), .CP(clk), .RN(n6), .Q(rd_data[8]) );
  HS65_LS_DFPRQX9 \rd_data_reg[7]  ( .D(N25), .CP(clk), .RN(n6), .Q(rd_data[7]) );
  HS65_LS_DFPRQX9 \rd_data_reg[6]  ( .D(N26), .CP(clk), .RN(n6), .Q(rd_data[6]) );
  HS65_LS_DFPRQX9 \rd_data_reg[5]  ( .D(N27), .CP(clk), .RN(n6), .Q(rd_data[5]) );
  HS65_LS_DFPRQX9 \rd_data_reg[4]  ( .D(N28), .CP(clk), .RN(n6), .Q(rd_data[4]) );
  HS65_LS_DFPRQX9 \rd_data_reg[3]  ( .D(N29), .CP(clk), .RN(n6), .Q(rd_data[3]) );
  HS65_LS_DFPRQX9 \rd_data_reg[2]  ( .D(N30), .CP(clk), .RN(n6), .Q(rd_data[2]) );
  HS65_LS_DFPRQX9 \rd_data_reg[1]  ( .D(N31), .CP(clk), .RN(n7), .Q(rd_data[1]) );
  HS65_LS_DFPRQX9 \rd_data_reg[0]  ( .D(N32), .CP(clk), .RN(n7), .Q(rd_data[0]) );
  HS65_LS_BFX9 U3 ( .A(n81), .Z(n4) );
  HS65_LS_BFX9 U4 ( .A(n81), .Z(n3) );
  HS65_LS_BFX9 U5 ( .A(n81), .Z(n2) );
  HS65_LS_BFX9 U6 ( .A(n83), .Z(n81) );
  HS65_LS_BFX9 U7 ( .A(n8), .Z(n6) );
  HS65_LS_BFX9 U8 ( .A(n8), .Z(n5) );
  HS65_LS_BFX9 U9 ( .A(n82), .Z(n1) );
  HS65_LS_BFX9 U10 ( .A(n83), .Z(n82) );
  HS65_LS_BFX9 U11 ( .A(n8), .Z(n7) );
  HS65_LS_BFX9 U12 ( .A(n83), .Z(n8) );
  HS65_LS_IVX9 U13 ( .A(reset), .Z(n83) );
  HS65_LS_IVX9 U14 ( .A(n161), .Z(n85) );
  HS65_LS_IVX9 U15 ( .A(n162), .Z(n84) );
  HS65_LS_NAND3X5 U16 ( .A(wr_ena), .B(n86), .C(wr_addr[0]), .Z(n161) );
  HS65_LS_IVX9 U17 ( .A(wr_addr[0]), .Z(n89) );
  HS65_LS_NAND3X5 U18 ( .A(n89), .B(n86), .C(wr_ena), .Z(n162) );
  HS65_LS_IVX9 U19 ( .A(n160), .Z(n88) );
  HS65_LS_IVX9 U20 ( .A(n159), .Z(n87) );
  HS65_LS_NAND3X5 U21 ( .A(wr_ena), .B(n89), .C(wr_addr[1]), .Z(n160) );
  HS65_LS_NOR2X6 U22 ( .A(n90), .B(rd_addr[1]), .Z(n157) );
  HS65_LS_NOR2X6 U23 ( .A(rd_addr[0]), .B(rd_addr[1]), .Z(n158) );
  HS65_LS_IVX9 U24 ( .A(wr_addr[1]), .Z(n86) );
  HS65_LS_NAND3X5 U25 ( .A(wr_addr[0]), .B(wr_ena), .C(wr_addr[1]), .Z(n159)
         );
  HS65_LS_AND2X4 U26 ( .A(rd_addr[1]), .B(n90), .Z(n156) );
  HS65_LS_IVX9 U27 ( .A(rd_addr[0]), .Z(n90) );
  HS65_LS_AND2X4 U28 ( .A(rd_addr[1]), .B(rd_addr[0]), .Z(n155) );
  HS65_LS_MX41X7 U29 ( .D0(n158), .S0(\mem[0][0] ), .D1(n157), .S1(\mem[1][0] ), .D2(n156), .S2(\mem[2][0] ), .D3(n155), .S3(\mem[3][0] ), .Z(N32) );
  HS65_LS_MX41X7 U30 ( .D0(n158), .S0(\mem[0][1] ), .D1(n157), .S1(\mem[1][1] ), .D2(n156), .S2(\mem[2][1] ), .D3(n155), .S3(\mem[3][1] ), .Z(N31) );
  HS65_LS_MX41X7 U31 ( .D0(n158), .S0(\mem[0][2] ), .D1(n157), .S1(\mem[1][2] ), .D2(n156), .S2(\mem[2][2] ), .D3(n155), .S3(\mem[3][2] ), .Z(N30) );
  HS65_LS_MX41X7 U32 ( .D0(n158), .S0(\mem[0][3] ), .D1(n157), .S1(\mem[1][3] ), .D2(n156), .S2(\mem[2][3] ), .D3(n155), .S3(\mem[3][3] ), .Z(N29) );
  HS65_LS_MX41X7 U33 ( .D0(n158), .S0(\mem[0][4] ), .D1(n157), .S1(\mem[1][4] ), .D2(n156), .S2(\mem[2][4] ), .D3(n155), .S3(\mem[3][4] ), .Z(N28) );
  HS65_LS_MX41X7 U34 ( .D0(n158), .S0(\mem[0][5] ), .D1(n157), .S1(\mem[1][5] ), .D2(n156), .S2(\mem[2][5] ), .D3(n155), .S3(\mem[3][5] ), .Z(N27) );
  HS65_LS_MX41X7 U35 ( .D0(n158), .S0(\mem[0][6] ), .D1(n157), .S1(\mem[1][6] ), .D2(n156), .S2(\mem[2][6] ), .D3(n155), .S3(\mem[3][6] ), .Z(N26) );
  HS65_LS_MX41X7 U36 ( .D0(n158), .S0(\mem[0][7] ), .D1(n157), .S1(\mem[1][7] ), .D2(n156), .S2(\mem[2][7] ), .D3(n155), .S3(\mem[3][7] ), .Z(N25) );
  HS65_LS_MX41X7 U37 ( .D0(n158), .S0(\mem[0][8] ), .D1(n157), .S1(\mem[1][8] ), .D2(n156), .S2(\mem[2][8] ), .D3(n155), .S3(\mem[3][8] ), .Z(N24) );
  HS65_LS_MX41X7 U38 ( .D0(n158), .S0(\mem[0][9] ), .D1(n157), .S1(\mem[1][9] ), .D2(n156), .S2(\mem[2][9] ), .D3(n155), .S3(\mem[3][9] ), .Z(N23) );
  HS65_LS_MX41X7 U39 ( .D0(n158), .S0(\mem[0][10] ), .D1(n157), .S1(
        \mem[1][10] ), .D2(n156), .S2(\mem[2][10] ), .D3(n155), .S3(
        \mem[3][10] ), .Z(N22) );
  HS65_LS_MX41X7 U40 ( .D0(n158), .S0(\mem[0][11] ), .D1(n157), .S1(
        \mem[1][11] ), .D2(n156), .S2(\mem[2][11] ), .D3(n155), .S3(
        \mem[3][11] ), .Z(N21) );
  HS65_LS_MX41X7 U41 ( .D0(n158), .S0(\mem[0][12] ), .D1(n157), .S1(
        \mem[1][12] ), .D2(n156), .S2(\mem[2][12] ), .D3(n155), .S3(
        \mem[3][12] ), .Z(N20) );
  HS65_LS_MX41X7 U42 ( .D0(n158), .S0(\mem[0][13] ), .D1(n157), .S1(
        \mem[1][13] ), .D2(n156), .S2(\mem[2][13] ), .D3(n155), .S3(
        \mem[3][13] ), .Z(N19) );
  HS65_LS_MX41X7 U43 ( .D0(n158), .S0(\mem[0][14] ), .D1(n157), .S1(
        \mem[1][14] ), .D2(n156), .S2(\mem[2][14] ), .D3(n155), .S3(
        \mem[3][14] ), .Z(N18) );
  HS65_LS_MX41X7 U44 ( .D0(n158), .S0(\mem[0][15] ), .D1(n157), .S1(
        \mem[1][15] ), .D2(n156), .S2(\mem[2][15] ), .D3(n155), .S3(
        \mem[3][15] ), .Z(N17) );
  HS65_LS_AO22X9 U45 ( .A(wr_data[0]), .B(n85), .C(n161), .D(\mem[1][0] ), .Z(
        n138) );
  HS65_LS_AO22X9 U46 ( .A(wr_data[1]), .B(n85), .C(n161), .D(\mem[1][1] ), .Z(
        n137) );
  HS65_LS_AO22X9 U47 ( .A(wr_data[2]), .B(n85), .C(n161), .D(\mem[1][2] ), .Z(
        n136) );
  HS65_LS_AO22X9 U48 ( .A(wr_data[3]), .B(n85), .C(n161), .D(\mem[1][3] ), .Z(
        n135) );
  HS65_LS_AO22X9 U49 ( .A(wr_data[4]), .B(n85), .C(n161), .D(\mem[1][4] ), .Z(
        n134) );
  HS65_LS_AO22X9 U50 ( .A(wr_data[5]), .B(n85), .C(n161), .D(\mem[1][5] ), .Z(
        n133) );
  HS65_LS_AO22X9 U51 ( .A(wr_data[6]), .B(n85), .C(n161), .D(\mem[1][6] ), .Z(
        n132) );
  HS65_LS_AO22X9 U52 ( .A(wr_data[7]), .B(n85), .C(n161), .D(\mem[1][7] ), .Z(
        n131) );
  HS65_LS_AO22X9 U53 ( .A(wr_data[8]), .B(n85), .C(n161), .D(\mem[1][8] ), .Z(
        n130) );
  HS65_LS_AO22X9 U54 ( .A(wr_data[9]), .B(n85), .C(n161), .D(\mem[1][9] ), .Z(
        n129) );
  HS65_LS_AO22X9 U55 ( .A(wr_data[10]), .B(n85), .C(n161), .D(\mem[1][10] ), 
        .Z(n128) );
  HS65_LS_AO22X9 U56 ( .A(wr_data[11]), .B(n85), .C(n161), .D(\mem[1][11] ), 
        .Z(n127) );
  HS65_LS_AO22X9 U57 ( .A(wr_data[12]), .B(n85), .C(n161), .D(\mem[1][12] ), 
        .Z(n126) );
  HS65_LS_AO22X9 U58 ( .A(wr_data[13]), .B(n85), .C(n161), .D(\mem[1][13] ), 
        .Z(n125) );
  HS65_LS_AO22X9 U59 ( .A(wr_data[14]), .B(n85), .C(n161), .D(\mem[1][14] ), 
        .Z(n124) );
  HS65_LS_AO22X9 U60 ( .A(wr_data[15]), .B(n85), .C(n161), .D(\mem[1][15] ), 
        .Z(n123) );
  HS65_LS_AO22X9 U61 ( .A(wr_data[0]), .B(n88), .C(n160), .D(\mem[2][0] ), .Z(
        n122) );
  HS65_LS_AO22X9 U62 ( .A(wr_data[1]), .B(n88), .C(n160), .D(\mem[2][1] ), .Z(
        n121) );
  HS65_LS_AO22X9 U63 ( .A(wr_data[2]), .B(n88), .C(n160), .D(\mem[2][2] ), .Z(
        n120) );
  HS65_LS_AO22X9 U64 ( .A(wr_data[3]), .B(n88), .C(n160), .D(\mem[2][3] ), .Z(
        n119) );
  HS65_LS_AO22X9 U65 ( .A(wr_data[4]), .B(n88), .C(n160), .D(\mem[2][4] ), .Z(
        n118) );
  HS65_LS_AO22X9 U66 ( .A(wr_data[5]), .B(n88), .C(n160), .D(\mem[2][5] ), .Z(
        n117) );
  HS65_LS_AO22X9 U67 ( .A(wr_data[6]), .B(n88), .C(n160), .D(\mem[2][6] ), .Z(
        n116) );
  HS65_LS_AO22X9 U68 ( .A(wr_data[7]), .B(n88), .C(n160), .D(\mem[2][7] ), .Z(
        n115) );
  HS65_LS_AO22X9 U69 ( .A(wr_data[8]), .B(n88), .C(n160), .D(\mem[2][8] ), .Z(
        n114) );
  HS65_LS_AO22X9 U70 ( .A(wr_data[9]), .B(n88), .C(n160), .D(\mem[2][9] ), .Z(
        n113) );
  HS65_LS_AO22X9 U71 ( .A(wr_data[10]), .B(n88), .C(n160), .D(\mem[2][10] ), 
        .Z(n112) );
  HS65_LS_AO22X9 U72 ( .A(wr_data[11]), .B(n88), .C(n160), .D(\mem[2][11] ), 
        .Z(n111) );
  HS65_LS_AO22X9 U73 ( .A(wr_data[12]), .B(n88), .C(n160), .D(\mem[2][12] ), 
        .Z(n110) );
  HS65_LS_AO22X9 U74 ( .A(wr_data[13]), .B(n88), .C(n160), .D(\mem[2][13] ), 
        .Z(n109) );
  HS65_LS_AO22X9 U75 ( .A(wr_data[14]), .B(n88), .C(n160), .D(\mem[2][14] ), 
        .Z(n108) );
  HS65_LS_AO22X9 U76 ( .A(wr_data[15]), .B(n88), .C(n160), .D(\mem[2][15] ), 
        .Z(n107) );
  HS65_LS_AO22X9 U77 ( .A(n84), .B(wr_data[0]), .C(n162), .D(\mem[0][0] ), .Z(
        n154) );
  HS65_LS_AO22X9 U78 ( .A(n84), .B(wr_data[1]), .C(n162), .D(\mem[0][1] ), .Z(
        n153) );
  HS65_LS_AO22X9 U79 ( .A(n84), .B(wr_data[2]), .C(n162), .D(\mem[0][2] ), .Z(
        n152) );
  HS65_LS_AO22X9 U80 ( .A(n84), .B(wr_data[3]), .C(n162), .D(\mem[0][3] ), .Z(
        n151) );
  HS65_LS_AO22X9 U81 ( .A(n84), .B(wr_data[4]), .C(n162), .D(\mem[0][4] ), .Z(
        n150) );
  HS65_LS_AO22X9 U82 ( .A(n84), .B(wr_data[5]), .C(n162), .D(\mem[0][5] ), .Z(
        n149) );
  HS65_LS_AO22X9 U83 ( .A(n84), .B(wr_data[6]), .C(n162), .D(\mem[0][6] ), .Z(
        n148) );
  HS65_LS_AO22X9 U84 ( .A(n84), .B(wr_data[7]), .C(n162), .D(\mem[0][7] ), .Z(
        n147) );
  HS65_LS_AO22X9 U85 ( .A(n84), .B(wr_data[8]), .C(n162), .D(\mem[0][8] ), .Z(
        n146) );
  HS65_LS_AO22X9 U86 ( .A(n84), .B(wr_data[9]), .C(n162), .D(\mem[0][9] ), .Z(
        n145) );
  HS65_LS_AO22X9 U87 ( .A(n84), .B(wr_data[10]), .C(n162), .D(\mem[0][10] ), 
        .Z(n144) );
  HS65_LS_AO22X9 U88 ( .A(n84), .B(wr_data[11]), .C(n162), .D(\mem[0][11] ), 
        .Z(n143) );
  HS65_LS_AO22X9 U89 ( .A(n84), .B(wr_data[12]), .C(n162), .D(\mem[0][12] ), 
        .Z(n142) );
  HS65_LS_AO22X9 U90 ( .A(n84), .B(wr_data[13]), .C(n162), .D(\mem[0][13] ), 
        .Z(n141) );
  HS65_LS_AO22X9 U91 ( .A(n84), .B(wr_data[14]), .C(n162), .D(\mem[0][14] ), 
        .Z(n140) );
  HS65_LS_AO22X9 U92 ( .A(n84), .B(wr_data[15]), .C(n162), .D(\mem[0][15] ), 
        .Z(n139) );
  HS65_LS_AO22X9 U93 ( .A(wr_data[0]), .B(n87), .C(n159), .D(\mem[3][0] ), .Z(
        n106) );
  HS65_LS_AO22X9 U94 ( .A(wr_data[1]), .B(n87), .C(n159), .D(\mem[3][1] ), .Z(
        n105) );
  HS65_LS_AO22X9 U95 ( .A(wr_data[2]), .B(n87), .C(n159), .D(\mem[3][2] ), .Z(
        n104) );
  HS65_LS_AO22X9 U96 ( .A(wr_data[3]), .B(n87), .C(n159), .D(\mem[3][3] ), .Z(
        n103) );
  HS65_LS_AO22X9 U97 ( .A(wr_data[4]), .B(n87), .C(n159), .D(\mem[3][4] ), .Z(
        n102) );
  HS65_LS_AO22X9 U98 ( .A(wr_data[5]), .B(n87), .C(n159), .D(\mem[3][5] ), .Z(
        n101) );
  HS65_LS_AO22X9 U99 ( .A(wr_data[6]), .B(n87), .C(n159), .D(\mem[3][6] ), .Z(
        n100) );
  HS65_LS_AO22X9 U100 ( .A(wr_data[7]), .B(n87), .C(n159), .D(\mem[3][7] ), 
        .Z(n99) );
  HS65_LS_AO22X9 U101 ( .A(wr_data[8]), .B(n87), .C(n159), .D(\mem[3][8] ), 
        .Z(n98) );
  HS65_LS_AO22X9 U102 ( .A(wr_data[9]), .B(n87), .C(n159), .D(\mem[3][9] ), 
        .Z(n97) );
  HS65_LS_AO22X9 U103 ( .A(wr_data[10]), .B(n87), .C(n159), .D(\mem[3][10] ), 
        .Z(n96) );
  HS65_LS_AO22X9 U104 ( .A(wr_data[11]), .B(n87), .C(n159), .D(\mem[3][11] ), 
        .Z(n95) );
  HS65_LS_AO22X9 U105 ( .A(wr_data[12]), .B(n87), .C(n159), .D(\mem[3][12] ), 
        .Z(n94) );
  HS65_LS_AO22X9 U106 ( .A(wr_data[13]), .B(n87), .C(n159), .D(\mem[3][13] ), 
        .Z(n93) );
  HS65_LS_AO22X9 U107 ( .A(wr_data[14]), .B(n87), .C(n159), .D(\mem[3][14] ), 
        .Z(n92) );
  HS65_LS_AO22X9 U108 ( .A(wr_data[15]), .B(n87), .C(n159), .D(\mem[3][15] ), 
        .Z(n91) );
endmodule


module dma_sdp_DATA64_ADDR2_2 ( clk, reset, ren, wen, waddr, wdata, raddr, 
        rdata );
  input [2:0] ren;
  input [2:0] wen;
  input [1:0] waddr;
  input [63:0] wdata;
  input [1:0] raddr;
  output [63:0] rdata;
  input clk, reset;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n41, n42, n43, n44, n45, n46, n47, n48;
  wire   [2:0] sel_out;
  wire   [15:0] rdata0;
  wire   [31:0] rdata1;
  wire   [15:0] rdata2;

  HS65_LS_DFPRQX9 \sel_out_reg[2]  ( .D(ren[2]), .CP(clk), .RN(n5), .Q(
        sel_out[2]) );
  HS65_LS_DFPRQX9 \sel_out_reg[1]  ( .D(ren[1]), .CP(clk), .RN(n5), .Q(
        sel_out[1]) );
  HS65_LS_DFPRQX9 \sel_out_reg[0]  ( .D(ren[0]), .CP(clk), .RN(n5), .Q(
        sel_out[0]) );
  bram_DATA16_ADDR2_4 dma0 ( .clk(clk), .reset(reset), .rd_addr(raddr), 
        .wr_addr(waddr), .wr_data(wdata[63:48]), .wr_ena(wen[2]), .rd_data(
        rdata0) );
  bram_DATA32_ADDR2_2 dma1 ( .clk(clk), .reset(reset), .rd_addr(raddr), 
        .wr_addr(waddr), .wr_data(wdata[47:16]), .wr_ena(wen[1]), .rd_data(
        rdata1) );
  bram_DATA16_ADDR2_3 dma2 ( .clk(clk), .reset(reset), .rd_addr(raddr), 
        .wr_addr(waddr), .wr_data(wdata[15:0]), .wr_ena(wen[0]), .rd_data(
        rdata2) );
  HS65_LS_NAND3X5 U3 ( .A(sel_out[2]), .B(sel_out[1]), .C(sel_out[0]), .Z(n46)
         );
  HS65_LS_IVX9 U4 ( .A(reset), .Z(n5) );
  HS65_LS_NOR2X6 U5 ( .A(n2), .B(n13), .Z(rdata[40]) );
  HS65_LS_NOR2X6 U6 ( .A(n2), .B(n12), .Z(rdata[41]) );
  HS65_LS_NOR2X6 U7 ( .A(n2), .B(n11), .Z(rdata[42]) );
  HS65_LS_NOR2X6 U8 ( .A(n2), .B(n10), .Z(rdata[43]) );
  HS65_LS_NOR2X6 U9 ( .A(n2), .B(n9), .Z(rdata[44]) );
  HS65_LS_NOR2X6 U10 ( .A(n2), .B(n8), .Z(rdata[45]) );
  HS65_LS_NOR2X6 U11 ( .A(n2), .B(n14), .Z(rdata[39]) );
  HS65_LS_BFX9 U12 ( .A(n46), .Z(n2) );
  HS65_LS_NOR2X6 U13 ( .A(n2), .B(n15), .Z(rdata[38]) );
  HS65_LS_NOR2X6 U14 ( .A(n3), .B(n19), .Z(rdata[34]) );
  HS65_LS_NOR2X6 U15 ( .A(n2), .B(n18), .Z(rdata[35]) );
  HS65_LS_NOR2X6 U16 ( .A(n3), .B(n17), .Z(rdata[36]) );
  HS65_LS_NOR2X6 U17 ( .A(n2), .B(n16), .Z(rdata[37]) );
  HS65_LS_NOR2X6 U18 ( .A(n3), .B(n20), .Z(rdata[33]) );
  HS65_LS_BFX9 U19 ( .A(n46), .Z(n3) );
  HS65_LS_BFX9 U20 ( .A(n46), .Z(n1) );
  HS65_LS_BFX9 U21 ( .A(n46), .Z(n4) );
  HS65_LS_IVX9 U22 ( .A(n45), .Z(n42) );
  HS65_LS_NOR2X6 U23 ( .A(n2), .B(n7), .Z(rdata[46]) );
  HS65_LS_NOR2X6 U24 ( .A(n2), .B(n6), .Z(rdata[47]) );
  HS65_LS_NAND3X5 U25 ( .A(n44), .B(n43), .C(sel_out[1]), .Z(n45) );
  HS65_LS_IVX9 U26 ( .A(sel_out[0]), .Z(n44) );
  HS65_LS_IVX9 U27 ( .A(sel_out[2]), .Z(n43) );
  HS65_LS_OAI22X6 U28 ( .A(n45), .B(n19), .C(n1), .D(n35), .Z(rdata[18]) );
  HS65_LS_IVX9 U29 ( .A(rdata1[2]), .Z(n35) );
  HS65_LS_OAI22X6 U30 ( .A(n45), .B(n18), .C(n1), .D(n34), .Z(rdata[19]) );
  HS65_LS_IVX9 U31 ( .A(rdata1[3]), .Z(n34) );
  HS65_LS_OAI22X6 U32 ( .A(n45), .B(n17), .C(n1), .D(n33), .Z(rdata[20]) );
  HS65_LS_IVX9 U33 ( .A(rdata1[4]), .Z(n33) );
  HS65_LS_OAI22X6 U34 ( .A(n45), .B(n16), .C(n1), .D(n32), .Z(rdata[21]) );
  HS65_LS_IVX9 U35 ( .A(rdata1[5]), .Z(n32) );
  HS65_LS_OAI22X6 U36 ( .A(n45), .B(n15), .C(n31), .D(n3), .Z(rdata[22]) );
  HS65_LS_IVX9 U37 ( .A(rdata1[6]), .Z(n31) );
  HS65_LS_OAI22X6 U38 ( .A(n45), .B(n14), .C(n30), .D(n3), .Z(rdata[23]) );
  HS65_LS_IVX9 U39 ( .A(rdata1[7]), .Z(n30) );
  HS65_LS_OAI22X6 U40 ( .A(n45), .B(n13), .C(n29), .D(n3), .Z(rdata[24]) );
  HS65_LS_IVX9 U41 ( .A(rdata1[8]), .Z(n29) );
  HS65_LS_OAI22X6 U42 ( .A(n45), .B(n12), .C(n28), .D(n3), .Z(rdata[25]) );
  HS65_LS_IVX9 U43 ( .A(rdata1[9]), .Z(n28) );
  HS65_LS_OAI22X6 U44 ( .A(n45), .B(n11), .C(n1), .D(n27), .Z(rdata[26]) );
  HS65_LS_IVX9 U45 ( .A(rdata1[10]), .Z(n27) );
  HS65_LS_OAI22X6 U46 ( .A(n45), .B(n10), .C(n1), .D(n26), .Z(rdata[27]) );
  HS65_LS_IVX9 U47 ( .A(rdata1[11]), .Z(n26) );
  HS65_LS_OAI22X6 U48 ( .A(n45), .B(n20), .C(n1), .D(n36), .Z(rdata[17]) );
  HS65_LS_IVX9 U49 ( .A(rdata1[1]), .Z(n36) );
  HS65_LS_NOR2X6 U50 ( .A(n3), .B(n21), .Z(rdata[32]) );
  HS65_LS_NOR2AX3 U51 ( .A(rdata0[15]), .B(n3), .Z(rdata[63]) );
  HS65_LS_IVX9 U52 ( .A(rdata1[18]), .Z(n19) );
  HS65_LS_IVX9 U53 ( .A(rdata1[19]), .Z(n18) );
  HS65_LS_IVX9 U54 ( .A(rdata1[17]), .Z(n20) );
  HS65_LS_NOR2AX3 U55 ( .A(rdata0[3]), .B(n3), .Z(rdata[51]) );
  HS65_LS_NOR2AX3 U56 ( .A(rdata0[4]), .B(n4), .Z(rdata[52]) );
  HS65_LS_NOR2AX3 U57 ( .A(rdata0[7]), .B(n4), .Z(rdata[55]) );
  HS65_LS_NOR2AX3 U58 ( .A(rdata0[8]), .B(n4), .Z(rdata[56]) );
  HS65_LS_NOR2AX3 U59 ( .A(rdata0[10]), .B(n4), .Z(rdata[58]) );
  HS65_LS_NOR2AX3 U60 ( .A(rdata0[1]), .B(n3), .Z(rdata[49]) );
  HS65_LS_NOR2AX3 U61 ( .A(rdata0[2]), .B(n3), .Z(rdata[50]) );
  HS65_LS_NOR2AX3 U62 ( .A(rdata0[5]), .B(n4), .Z(rdata[53]) );
  HS65_LS_NOR2AX3 U63 ( .A(rdata0[6]), .B(n4), .Z(rdata[54]) );
  HS65_LS_NOR2AX3 U64 ( .A(rdata0[9]), .B(n4), .Z(rdata[57]) );
  HS65_LS_NOR2AX3 U65 ( .A(rdata0[11]), .B(n4), .Z(rdata[59]) );
  HS65_LS_NOR2AX3 U66 ( .A(rdata0[14]), .B(n4), .Z(rdata[62]) );
  HS65_LS_OAI31X5 U67 ( .A(n44), .B(sel_out[2]), .C(sel_out[1]), .D(n2), .Z(
        n47) );
  HS65_LS_NOR3X4 U68 ( .A(sel_out[0]), .B(sel_out[1]), .C(n43), .Z(n48) );
  HS65_LS_OAI22X6 U69 ( .A(n45), .B(n9), .C(n1), .D(n25), .Z(rdata[28]) );
  HS65_LS_IVX9 U70 ( .A(rdata1[12]), .Z(n25) );
  HS65_LS_OAI22X6 U71 ( .A(n45), .B(n8), .C(n1), .D(n24), .Z(rdata[29]) );
  HS65_LS_IVX9 U72 ( .A(rdata1[13]), .Z(n24) );
  HS65_LS_OAI22X6 U73 ( .A(n45), .B(n7), .C(n1), .D(n23), .Z(rdata[30]) );
  HS65_LS_IVX9 U74 ( .A(rdata1[14]), .Z(n23) );
  HS65_LS_OAI22X6 U75 ( .A(n45), .B(n6), .C(n1), .D(n22), .Z(rdata[31]) );
  HS65_LS_IVX9 U76 ( .A(rdata1[15]), .Z(n22) );
  HS65_LS_OAI22X6 U77 ( .A(n45), .B(n21), .C(n1), .D(n41), .Z(rdata[16]) );
  HS65_LS_IVX9 U78 ( .A(rdata1[0]), .Z(n41) );
  HS65_LS_NOR2AX3 U79 ( .A(rdata0[0]), .B(n3), .Z(rdata[48]) );
  HS65_LS_IVX9 U80 ( .A(rdata1[20]), .Z(n17) );
  HS65_LS_IVX9 U81 ( .A(rdata1[21]), .Z(n16) );
  HS65_LS_IVX9 U82 ( .A(rdata1[22]), .Z(n15) );
  HS65_LS_IVX9 U83 ( .A(rdata1[23]), .Z(n14) );
  HS65_LS_IVX9 U84 ( .A(rdata1[24]), .Z(n13) );
  HS65_LS_IVX9 U85 ( .A(rdata1[25]), .Z(n12) );
  HS65_LS_IVX9 U86 ( .A(rdata1[26]), .Z(n11) );
  HS65_LS_IVX9 U87 ( .A(rdata1[27]), .Z(n10) );
  HS65_LS_IVX9 U88 ( .A(rdata1[28]), .Z(n9) );
  HS65_LS_IVX9 U89 ( .A(rdata1[29]), .Z(n8) );
  HS65_LS_IVX9 U90 ( .A(rdata1[30]), .Z(n7) );
  HS65_LS_IVX9 U91 ( .A(rdata1[31]), .Z(n6) );
  HS65_LS_IVX9 U92 ( .A(rdata1[16]), .Z(n21) );
  HS65_LS_AO222X4 U93 ( .A(rdata0[0]), .B(n48), .C(rdata1[0]), .D(n42), .E(
        rdata2[0]), .F(n47), .Z(rdata[0]) );
  HS65_LS_AO222X4 U94 ( .A(rdata0[1]), .B(n48), .C(rdata1[1]), .D(n42), .E(
        rdata2[1]), .F(n47), .Z(rdata[1]) );
  HS65_LS_AO222X4 U95 ( .A(rdata0[2]), .B(n48), .C(rdata1[2]), .D(n42), .E(
        rdata2[2]), .F(n47), .Z(rdata[2]) );
  HS65_LS_AO222X4 U96 ( .A(rdata0[3]), .B(n48), .C(rdata1[3]), .D(n42), .E(
        rdata2[3]), .F(n47), .Z(rdata[3]) );
  HS65_LS_AO222X4 U97 ( .A(rdata0[4]), .B(n48), .C(rdata1[4]), .D(n42), .E(
        rdata2[4]), .F(n47), .Z(rdata[4]) );
  HS65_LS_AO222X4 U98 ( .A(rdata0[5]), .B(n48), .C(rdata1[5]), .D(n42), .E(
        rdata2[5]), .F(n47), .Z(rdata[5]) );
  HS65_LS_AO222X4 U99 ( .A(rdata0[6]), .B(n48), .C(rdata1[6]), .D(n42), .E(
        rdata2[6]), .F(n47), .Z(rdata[6]) );
  HS65_LS_AO222X4 U100 ( .A(rdata0[7]), .B(n48), .C(rdata1[7]), .D(n42), .E(
        rdata2[7]), .F(n47), .Z(rdata[7]) );
  HS65_LS_AO222X4 U101 ( .A(rdata0[8]), .B(n48), .C(rdata1[8]), .D(n42), .E(
        rdata2[8]), .F(n47), .Z(rdata[8]) );
  HS65_LS_AO222X4 U102 ( .A(rdata0[9]), .B(n48), .C(rdata1[9]), .D(n42), .E(
        rdata2[9]), .F(n47), .Z(rdata[9]) );
  HS65_LS_AO222X4 U103 ( .A(rdata0[10]), .B(n48), .C(rdata1[10]), .D(n42), .E(
        rdata2[10]), .F(n47), .Z(rdata[10]) );
  HS65_LS_AO222X4 U104 ( .A(rdata0[11]), .B(n48), .C(rdata1[11]), .D(n42), .E(
        rdata2[11]), .F(n47), .Z(rdata[11]) );
  HS65_LS_AO222X4 U105 ( .A(rdata0[12]), .B(n48), .C(rdata1[12]), .D(n42), .E(
        rdata2[12]), .F(n47), .Z(rdata[12]) );
  HS65_LS_AO222X4 U106 ( .A(rdata0[13]), .B(n48), .C(rdata1[13]), .D(n42), .E(
        rdata2[13]), .F(n47), .Z(rdata[13]) );
  HS65_LS_AO222X4 U107 ( .A(rdata0[14]), .B(n48), .C(rdata1[14]), .D(n42), .E(
        rdata2[14]), .F(n47), .Z(rdata[14]) );
  HS65_LS_AO222X4 U108 ( .A(rdata0[15]), .B(n48), .C(rdata1[15]), .D(n42), .E(
        rdata2[15]), .F(n47), .Z(rdata[15]) );
  HS65_LS_NOR2AX3 U109 ( .A(rdata0[12]), .B(n4), .Z(rdata[60]) );
  HS65_LS_NOR2AX3 U110 ( .A(rdata0[13]), .B(n4), .Z(rdata[61]) );
endmodule


module bram_DATA5_ADDR3_2 ( clk, reset, rd_addr, wr_addr, wr_data, wr_ena, 
        rd_data );
  input [2:0] rd_addr;
  input [2:0] wr_addr;
  input [4:0] wr_data;
  output [4:0] rd_data;
  input clk, reset, wr_ena;
  wire   \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N34,
         N35, N36, N37, N38, n1, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218;

  HS65_LS_DFPRQX9 \mem_reg[5][4]  ( .D(n131), .CP(clk), .RN(n1), .Q(
        \mem[5][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[5][3]  ( .D(n132), .CP(clk), .RN(n1), .Q(
        \mem[5][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[5][2]  ( .D(n133), .CP(clk), .RN(n1), .Q(
        \mem[5][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[5][1]  ( .D(n134), .CP(clk), .RN(n1), .Q(
        \mem[5][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[5][0]  ( .D(n135), .CP(clk), .RN(n22), .Q(
        \mem[5][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[4][4]  ( .D(n136), .CP(clk), .RN(n22), .Q(
        \mem[4][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[4][3]  ( .D(n137), .CP(clk), .RN(n22), .Q(
        \mem[4][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[4][2]  ( .D(n138), .CP(clk), .RN(n22), .Q(
        \mem[4][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[4][1]  ( .D(n139), .CP(clk), .RN(n22), .Q(
        \mem[4][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[4][0]  ( .D(n140), .CP(clk), .RN(n22), .Q(
        \mem[4][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][4]  ( .D(n151), .CP(clk), .RN(n22), .Q(
        \mem[1][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][3]  ( .D(n152), .CP(clk), .RN(n22), .Q(
        \mem[1][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][2]  ( .D(n153), .CP(clk), .RN(n22), .Q(
        \mem[1][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][1]  ( .D(n154), .CP(clk), .RN(n22), .Q(
        \mem[1][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][0]  ( .D(n155), .CP(clk), .RN(n22), .Q(
        \mem[1][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][4]  ( .D(n156), .CP(clk), .RN(n22), .Q(
        \mem[0][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][3]  ( .D(n157), .CP(clk), .RN(n1), .Q(
        \mem[0][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][2]  ( .D(n158), .CP(clk), .RN(n1), .Q(
        \mem[0][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][1]  ( .D(n159), .CP(clk), .RN(n1), .Q(
        \mem[0][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][0]  ( .D(n160), .CP(clk), .RN(n1), .Q(
        \mem[0][0] ) );
  HS65_LS_DFPRQX9 \rd_data_reg[4]  ( .D(N34), .CP(clk), .RN(n1), .Q(rd_data[4]) );
  HS65_LS_DFPRQX9 \rd_data_reg[3]  ( .D(N35), .CP(clk), .RN(n1), .Q(rd_data[3]) );
  HS65_LS_DFPRQX9 \rd_data_reg[2]  ( .D(N36), .CP(clk), .RN(n1), .Q(rd_data[2]) );
  HS65_LS_DFPRQX9 \rd_data_reg[1]  ( .D(N37), .CP(clk), .RN(n1), .Q(rd_data[1]) );
  HS65_LS_DFPRQX9 \rd_data_reg[0]  ( .D(N38), .CP(clk), .RN(n1), .Q(rd_data[0]) );
  HS65_LS_DFPRQNX9 \mem_reg[7][4]  ( .D(n121), .CP(clk), .RN(n23), .QN(n218)
         );
  HS65_LS_DFPRQNX9 \mem_reg[7][3]  ( .D(n122), .CP(clk), .RN(n22), .QN(n217)
         );
  HS65_LS_DFPRQNX9 \mem_reg[7][2]  ( .D(n123), .CP(clk), .RN(n24), .QN(n216)
         );
  HS65_LS_DFPRQNX9 \mem_reg[7][1]  ( .D(n124), .CP(clk), .RN(n24), .QN(n215)
         );
  HS65_LS_DFPRQNX9 \mem_reg[7][0]  ( .D(n125), .CP(clk), .RN(n24), .QN(n214)
         );
  HS65_LS_DFPRQNX9 \mem_reg[3][4]  ( .D(n141), .CP(clk), .RN(n23), .QN(n208)
         );
  HS65_LS_DFPRQNX9 \mem_reg[3][3]  ( .D(n142), .CP(clk), .RN(n23), .QN(n207)
         );
  HS65_LS_DFPRQNX9 \mem_reg[3][2]  ( .D(n143), .CP(clk), .RN(n23), .QN(n206)
         );
  HS65_LS_DFPRQNX9 \mem_reg[3][1]  ( .D(n144), .CP(clk), .RN(n23), .QN(n205)
         );
  HS65_LS_DFPRQNX9 \mem_reg[3][0]  ( .D(n145), .CP(clk), .RN(n23), .QN(n204)
         );
  HS65_LS_DFPRQNX9 \mem_reg[6][4]  ( .D(n126), .CP(clk), .RN(n24), .QN(n213)
         );
  HS65_LS_DFPRQNX9 \mem_reg[6][3]  ( .D(n127), .CP(clk), .RN(n24), .QN(n212)
         );
  HS65_LS_DFPRQNX9 \mem_reg[6][2]  ( .D(n128), .CP(clk), .RN(n23), .QN(n211)
         );
  HS65_LS_DFPRQNX9 \mem_reg[6][1]  ( .D(n129), .CP(clk), .RN(n23), .QN(n210)
         );
  HS65_LS_DFPRQNX9 \mem_reg[6][0]  ( .D(n130), .CP(clk), .RN(n23), .QN(n209)
         );
  HS65_LS_DFPRQNX9 \mem_reg[2][4]  ( .D(n146), .CP(clk), .RN(n23), .QN(n203)
         );
  HS65_LS_DFPRQNX9 \mem_reg[2][3]  ( .D(n147), .CP(clk), .RN(n23), .QN(n202)
         );
  HS65_LS_DFPRQNX9 \mem_reg[2][2]  ( .D(n148), .CP(clk), .RN(n23), .QN(n201)
         );
  HS65_LS_DFPRQNX9 \mem_reg[2][1]  ( .D(n149), .CP(clk), .RN(n23), .QN(n200)
         );
  HS65_LS_DFPRQNX9 \mem_reg[2][0]  ( .D(n150), .CP(clk), .RN(n23), .QN(n199)
         );
  HS65_LS_BFX9 U3 ( .A(n25), .Z(n1) );
  HS65_LS_BFX9 U4 ( .A(n25), .Z(n22) );
  HS65_LS_BFX9 U5 ( .A(n25), .Z(n23) );
  HS65_LS_BFX9 U6 ( .A(n25), .Z(n24) );
  HS65_LS_IVX9 U7 ( .A(reset), .Z(n25) );
  HS65_LS_IVX9 U8 ( .A(n198), .Z(n35) );
  HS65_LS_IVX9 U9 ( .A(n193), .Z(n31) );
  HS65_LS_IVX9 U10 ( .A(n194), .Z(n32) );
  HS65_LS_IVX9 U11 ( .A(n190), .Z(n29) );
  HS65_LS_IVX9 U12 ( .A(n189), .Z(n28) );
  HS65_LS_IVX9 U13 ( .A(n195), .Z(n33) );
  HS65_LS_NAND3X5 U14 ( .A(n37), .B(n36), .C(n197), .Z(n198) );
  HS65_LS_NAND3X5 U15 ( .A(n37), .B(n36), .C(n192), .Z(n193) );
  HS65_LS_IVX9 U16 ( .A(n191), .Z(n30) );
  HS65_LS_IVX9 U17 ( .A(n196), .Z(n34) );
  HS65_LS_NOR3X4 U18 ( .A(n26), .B(rd_addr[1]), .C(n27), .Z(n186) );
  HS65_LS_NOR3X4 U19 ( .A(rd_addr[1]), .B(rd_addr[2]), .C(n26), .Z(n181) );
  HS65_LS_NOR3X4 U20 ( .A(rd_addr[1]), .B(rd_addr[2]), .C(rd_addr[0]), .Z(n180) );
  HS65_LS_NOR3X4 U21 ( .A(rd_addr[0]), .B(rd_addr[1]), .C(n27), .Z(n185) );
  HS65_LS_NAND3X5 U22 ( .A(n26), .B(n27), .C(rd_addr[1]), .Z(n178) );
  HS65_LS_NAND3X5 U23 ( .A(rd_addr[0]), .B(n27), .C(rd_addr[1]), .Z(n177) );
  HS65_LS_NAND3X5 U24 ( .A(rd_addr[1]), .B(n26), .C(rd_addr[2]), .Z(n183) );
  HS65_LS_NAND3X5 U25 ( .A(rd_addr[1]), .B(rd_addr[0]), .C(rd_addr[2]), .Z(
        n182) );
  HS65_LS_OAI22X6 U26 ( .A(n199), .B(n178), .C(n204), .D(n177), .Z(n179) );
  HS65_LS_OAI22X6 U27 ( .A(n200), .B(n178), .C(n205), .D(n177), .Z(n173) );
  HS65_LS_OAI22X6 U28 ( .A(n201), .B(n178), .C(n206), .D(n177), .Z(n169) );
  HS65_LS_OAI22X6 U29 ( .A(n202), .B(n178), .C(n207), .D(n177), .Z(n165) );
  HS65_LS_OAI22X6 U30 ( .A(n203), .B(n178), .C(n208), .D(n177), .Z(n161) );
  HS65_LS_IVX9 U31 ( .A(rd_addr[0]), .Z(n26) );
  HS65_LS_IVX9 U32 ( .A(rd_addr[2]), .Z(n27) );
  HS65_LS_OAI22X6 U33 ( .A(n120), .B(n194), .C(n32), .D(n204), .Z(n145) );
  HS65_LS_OAI22X6 U34 ( .A(n119), .B(n194), .C(n32), .D(n205), .Z(n144) );
  HS65_LS_OAI22X6 U35 ( .A(n118), .B(n194), .C(n32), .D(n206), .Z(n143) );
  HS65_LS_OAI22X6 U36 ( .A(n117), .B(n194), .C(n32), .D(n207), .Z(n142) );
  HS65_LS_OAI22X6 U37 ( .A(n38), .B(n194), .C(n32), .D(n208), .Z(n141) );
  HS65_LS_OAI22X6 U38 ( .A(n120), .B(n190), .C(n29), .D(n209), .Z(n130) );
  HS65_LS_OAI22X6 U39 ( .A(n119), .B(n190), .C(n29), .D(n210), .Z(n129) );
  HS65_LS_OAI22X6 U40 ( .A(n118), .B(n190), .C(n29), .D(n211), .Z(n128) );
  HS65_LS_OAI22X6 U41 ( .A(n117), .B(n190), .C(n29), .D(n212), .Z(n127) );
  HS65_LS_OAI22X6 U42 ( .A(n38), .B(n190), .C(n29), .D(n213), .Z(n126) );
  HS65_LS_OAI22X6 U43 ( .A(n120), .B(n189), .C(n28), .D(n214), .Z(n125) );
  HS65_LS_OAI22X6 U44 ( .A(n119), .B(n189), .C(n28), .D(n215), .Z(n124) );
  HS65_LS_OAI22X6 U45 ( .A(n118), .B(n189), .C(n28), .D(n216), .Z(n123) );
  HS65_LS_OAI22X6 U46 ( .A(n117), .B(n189), .C(n28), .D(n217), .Z(n122) );
  HS65_LS_OAI22X6 U47 ( .A(n38), .B(n189), .C(n28), .D(n218), .Z(n121) );
  HS65_LS_OAI22X6 U48 ( .A(n120), .B(n195), .C(n33), .D(n199), .Z(n150) );
  HS65_LS_OAI22X6 U49 ( .A(n119), .B(n195), .C(n33), .D(n200), .Z(n149) );
  HS65_LS_OAI22X6 U50 ( .A(n118), .B(n195), .C(n33), .D(n201), .Z(n148) );
  HS65_LS_OAI22X6 U51 ( .A(n117), .B(n195), .C(n33), .D(n202), .Z(n147) );
  HS65_LS_OAI22X6 U52 ( .A(n38), .B(n195), .C(n33), .D(n203), .Z(n146) );
  HS65_LS_NAND2X7 U53 ( .A(n188), .B(n187), .Z(N38) );
  HS65_LS_AOI212X4 U54 ( .A(n186), .B(\mem[5][0] ), .C(n185), .D(\mem[4][0] ), 
        .E(n184), .Z(n187) );
  HS65_LS_AOI212X4 U55 ( .A(n181), .B(\mem[1][0] ), .C(n180), .D(\mem[0][0] ), 
        .E(n179), .Z(n188) );
  HS65_LS_OAI22X6 U56 ( .A(n209), .B(n183), .C(n214), .D(n182), .Z(n184) );
  HS65_LS_NAND2X7 U57 ( .A(n176), .B(n175), .Z(N37) );
  HS65_LS_AOI212X4 U58 ( .A(n186), .B(\mem[5][1] ), .C(n185), .D(\mem[4][1] ), 
        .E(n174), .Z(n175) );
  HS65_LS_AOI212X4 U59 ( .A(n181), .B(\mem[1][1] ), .C(n180), .D(\mem[0][1] ), 
        .E(n173), .Z(n176) );
  HS65_LS_OAI22X6 U60 ( .A(n210), .B(n183), .C(n215), .D(n182), .Z(n174) );
  HS65_LS_NAND2X7 U61 ( .A(n172), .B(n171), .Z(N36) );
  HS65_LS_AOI212X4 U62 ( .A(n186), .B(\mem[5][2] ), .C(n185), .D(\mem[4][2] ), 
        .E(n170), .Z(n171) );
  HS65_LS_AOI212X4 U63 ( .A(n181), .B(\mem[1][2] ), .C(n180), .D(\mem[0][2] ), 
        .E(n169), .Z(n172) );
  HS65_LS_OAI22X6 U64 ( .A(n211), .B(n183), .C(n216), .D(n182), .Z(n170) );
  HS65_LS_NAND2X7 U65 ( .A(n168), .B(n167), .Z(N35) );
  HS65_LS_AOI212X4 U66 ( .A(n186), .B(\mem[5][3] ), .C(n185), .D(\mem[4][3] ), 
        .E(n166), .Z(n167) );
  HS65_LS_AOI212X4 U67 ( .A(n181), .B(\mem[1][3] ), .C(n180), .D(\mem[0][3] ), 
        .E(n165), .Z(n168) );
  HS65_LS_OAI22X6 U68 ( .A(n212), .B(n183), .C(n217), .D(n182), .Z(n166) );
  HS65_LS_NAND2X7 U69 ( .A(n164), .B(n163), .Z(N34) );
  HS65_LS_AOI212X4 U70 ( .A(n186), .B(\mem[5][4] ), .C(n185), .D(\mem[4][4] ), 
        .E(n162), .Z(n163) );
  HS65_LS_AOI212X4 U71 ( .A(n181), .B(\mem[1][4] ), .C(n180), .D(\mem[0][4] ), 
        .E(n161), .Z(n164) );
  HS65_LS_OAI22X6 U72 ( .A(n213), .B(n183), .C(n218), .D(n182), .Z(n162) );
  HS65_LS_AO22X9 U73 ( .A(n35), .B(wr_data[0]), .C(n198), .D(\mem[0][0] ), .Z(
        n160) );
  HS65_LS_AO22X9 U74 ( .A(n35), .B(wr_data[1]), .C(n198), .D(\mem[0][1] ), .Z(
        n159) );
  HS65_LS_AO22X9 U75 ( .A(n35), .B(wr_data[2]), .C(n198), .D(\mem[0][2] ), .Z(
        n158) );
  HS65_LS_AO22X9 U76 ( .A(n35), .B(wr_data[3]), .C(n198), .D(\mem[0][3] ), .Z(
        n157) );
  HS65_LS_AO22X9 U77 ( .A(n35), .B(wr_data[4]), .C(n198), .D(\mem[0][4] ), .Z(
        n156) );
  HS65_LS_AO22X9 U78 ( .A(wr_data[0]), .B(n31), .C(n193), .D(\mem[4][0] ), .Z(
        n140) );
  HS65_LS_AO22X9 U79 ( .A(wr_data[1]), .B(n31), .C(n193), .D(\mem[4][1] ), .Z(
        n139) );
  HS65_LS_AO22X9 U80 ( .A(wr_data[2]), .B(n31), .C(n193), .D(\mem[4][2] ), .Z(
        n138) );
  HS65_LS_AO22X9 U81 ( .A(wr_data[3]), .B(n31), .C(n193), .D(\mem[4][3] ), .Z(
        n137) );
  HS65_LS_AO22X9 U82 ( .A(wr_data[4]), .B(n31), .C(n193), .D(\mem[4][4] ), .Z(
        n136) );
  HS65_LS_AO22X9 U83 ( .A(wr_data[0]), .B(n30), .C(n191), .D(\mem[5][0] ), .Z(
        n135) );
  HS65_LS_AO22X9 U84 ( .A(wr_data[1]), .B(n30), .C(n191), .D(\mem[5][1] ), .Z(
        n134) );
  HS65_LS_AO22X9 U85 ( .A(wr_data[2]), .B(n30), .C(n191), .D(\mem[5][2] ), .Z(
        n133) );
  HS65_LS_AO22X9 U86 ( .A(wr_data[3]), .B(n30), .C(n191), .D(\mem[5][3] ), .Z(
        n132) );
  HS65_LS_AO22X9 U87 ( .A(wr_data[4]), .B(n30), .C(n191), .D(\mem[5][4] ), .Z(
        n131) );
  HS65_LS_AO22X9 U88 ( .A(wr_data[0]), .B(n34), .C(n196), .D(\mem[1][0] ), .Z(
        n155) );
  HS65_LS_AO22X9 U89 ( .A(wr_data[1]), .B(n34), .C(n196), .D(\mem[1][1] ), .Z(
        n154) );
  HS65_LS_AO22X9 U90 ( .A(wr_data[2]), .B(n34), .C(n196), .D(\mem[1][2] ), .Z(
        n153) );
  HS65_LS_AO22X9 U91 ( .A(wr_data[3]), .B(n34), .C(n196), .D(\mem[1][3] ), .Z(
        n152) );
  HS65_LS_AO22X9 U92 ( .A(wr_data[4]), .B(n34), .C(n196), .D(\mem[1][4] ), .Z(
        n151) );
  HS65_LS_NAND3X5 U93 ( .A(wr_addr[0]), .B(n197), .C(wr_addr[1]), .Z(n194) );
  HS65_LS_NAND3X5 U94 ( .A(wr_addr[1]), .B(n37), .C(n192), .Z(n190) );
  HS65_LS_NAND3X5 U95 ( .A(wr_addr[1]), .B(wr_addr[0]), .C(n192), .Z(n189) );
  HS65_LS_NAND3X5 U96 ( .A(n197), .B(n37), .C(wr_addr[1]), .Z(n195) );
  HS65_LS_NOR2AX3 U97 ( .A(wr_ena), .B(wr_addr[2]), .Z(n197) );
  HS65_LS_NAND3X5 U98 ( .A(wr_addr[0]), .B(n36), .C(n192), .Z(n191) );
  HS65_LS_NAND3X5 U99 ( .A(n197), .B(n36), .C(wr_addr[0]), .Z(n196) );
  HS65_LS_IVX9 U100 ( .A(wr_addr[0]), .Z(n37) );
  HS65_LS_IVX9 U101 ( .A(wr_data[0]), .Z(n120) );
  HS65_LS_IVX9 U102 ( .A(wr_data[1]), .Z(n119) );
  HS65_LS_IVX9 U103 ( .A(wr_data[2]), .Z(n118) );
  HS65_LS_IVX9 U104 ( .A(wr_data[3]), .Z(n117) );
  HS65_LS_IVX9 U105 ( .A(wr_data[4]), .Z(n38) );
  HS65_LS_IVX9 U106 ( .A(wr_addr[1]), .Z(n36) );
  HS65_LS_AND2X4 U107 ( .A(wr_addr[2]), .B(wr_ena), .Z(n192) );
endmodule


module nAdapter_2 ( na_clk, na_reset, .proc_in({\proc_in[MCMD][1] , 
        \proc_in[MCMD][0] , \proc_in[MADDR][31] , \proc_in[MADDR][30] , 
        \proc_in[MADDR][29] , \proc_in[MADDR][28] , \proc_in[MADDR][27] , 
        \proc_in[MADDR][26] , \proc_in[MADDR][25] , \proc_in[MADDR][24] , 
        \proc_in[MADDR][23] , \proc_in[MADDR][22] , \proc_in[MADDR][21] , 
        \proc_in[MADDR][20] , \proc_in[MADDR][19] , \proc_in[MADDR][18] , 
        \proc_in[MADDR][17] , \proc_in[MADDR][16] , \proc_in[MADDR][15] , 
        \proc_in[MADDR][14] , \proc_in[MADDR][13] , \proc_in[MADDR][12] , 
        \proc_in[MADDR][11] , \proc_in[MADDR][10] , \proc_in[MADDR][9] , 
        \proc_in[MADDR][8] , \proc_in[MADDR][7] , \proc_in[MADDR][6] , 
        \proc_in[MADDR][5] , \proc_in[MADDR][4] , \proc_in[MADDR][3] , 
        \proc_in[MADDR][2] , \proc_in[MADDR][1] , \proc_in[MADDR][0] , 
        \proc_in[MDATA][31] , \proc_in[MDATA][30] , \proc_in[MDATA][29] , 
        \proc_in[MDATA][28] , \proc_in[MDATA][27] , \proc_in[MDATA][26] , 
        \proc_in[MDATA][25] , \proc_in[MDATA][24] , \proc_in[MDATA][23] , 
        \proc_in[MDATA][22] , \proc_in[MDATA][21] , \proc_in[MDATA][20] , 
        \proc_in[MDATA][19] , \proc_in[MDATA][18] , \proc_in[MDATA][17] , 
        \proc_in[MDATA][16] , \proc_in[MDATA][15] , \proc_in[MDATA][14] , 
        \proc_in[MDATA][13] , \proc_in[MDATA][12] , \proc_in[MDATA][11] , 
        \proc_in[MDATA][10] , \proc_in[MDATA][9] , \proc_in[MDATA][8] , 
        \proc_in[MDATA][7] , \proc_in[MDATA][6] , \proc_in[MDATA][5] , 
        \proc_in[MDATA][4] , \proc_in[MDATA][3] , \proc_in[MDATA][2] , 
        \proc_in[MDATA][1] , \proc_in[MDATA][0] }), .proc_out({
        \proc_out[SCMDACCEPT] , \proc_out[SRESP] , \proc_out[SDATA][31] , 
        \proc_out[SDATA][30] , \proc_out[SDATA][29] , \proc_out[SDATA][28] , 
        \proc_out[SDATA][27] , \proc_out[SDATA][26] , \proc_out[SDATA][25] , 
        \proc_out[SDATA][24] , \proc_out[SDATA][23] , \proc_out[SDATA][22] , 
        \proc_out[SDATA][21] , \proc_out[SDATA][20] , \proc_out[SDATA][19] , 
        \proc_out[SDATA][18] , \proc_out[SDATA][17] , \proc_out[SDATA][16] , 
        \proc_out[SDATA][15] , \proc_out[SDATA][14] , \proc_out[SDATA][13] , 
        \proc_out[SDATA][12] , \proc_out[SDATA][11] , \proc_out[SDATA][10] , 
        \proc_out[SDATA][9] , \proc_out[SDATA][8] , \proc_out[SDATA][7] , 
        \proc_out[SDATA][6] , \proc_out[SDATA][5] , \proc_out[SDATA][4] , 
        \proc_out[SDATA][3] , \proc_out[SDATA][2] , \proc_out[SDATA][1] , 
        \proc_out[SDATA][0] }), .spm_in({\spm_in[SCMDACCEPT] , \spm_in[SRESP] , 
        \spm_in[SDATA][63] , \spm_in[SDATA][62] , \spm_in[SDATA][61] , 
        \spm_in[SDATA][60] , \spm_in[SDATA][59] , \spm_in[SDATA][58] , 
        \spm_in[SDATA][57] , \spm_in[SDATA][56] , \spm_in[SDATA][55] , 
        \spm_in[SDATA][54] , \spm_in[SDATA][53] , \spm_in[SDATA][52] , 
        \spm_in[SDATA][51] , \spm_in[SDATA][50] , \spm_in[SDATA][49] , 
        \spm_in[SDATA][48] , \spm_in[SDATA][47] , \spm_in[SDATA][46] , 
        \spm_in[SDATA][45] , \spm_in[SDATA][44] , \spm_in[SDATA][43] , 
        \spm_in[SDATA][42] , \spm_in[SDATA][41] , \spm_in[SDATA][40] , 
        \spm_in[SDATA][39] , \spm_in[SDATA][38] , \spm_in[SDATA][37] , 
        \spm_in[SDATA][36] , \spm_in[SDATA][35] , \spm_in[SDATA][34] , 
        \spm_in[SDATA][33] , \spm_in[SDATA][32] , \spm_in[SDATA][31] , 
        \spm_in[SDATA][30] , \spm_in[SDATA][29] , \spm_in[SDATA][28] , 
        \spm_in[SDATA][27] , \spm_in[SDATA][26] , \spm_in[SDATA][25] , 
        \spm_in[SDATA][24] , \spm_in[SDATA][23] , \spm_in[SDATA][22] , 
        \spm_in[SDATA][21] , \spm_in[SDATA][20] , \spm_in[SDATA][19] , 
        \spm_in[SDATA][18] , \spm_in[SDATA][17] , \spm_in[SDATA][16] , 
        \spm_in[SDATA][15] , \spm_in[SDATA][14] , \spm_in[SDATA][13] , 
        \spm_in[SDATA][12] , \spm_in[SDATA][11] , \spm_in[SDATA][10] , 
        \spm_in[SDATA][9] , \spm_in[SDATA][8] , \spm_in[SDATA][7] , 
        \spm_in[SDATA][6] , \spm_in[SDATA][5] , \spm_in[SDATA][4] , 
        \spm_in[SDATA][3] , \spm_in[SDATA][2] , \spm_in[SDATA][1] , 
        \spm_in[SDATA][0] }), .spm_out({\spm_out[MCMD][1] , \spm_out[MCMD][0] , 
        \spm_out[MADDR][31] , \spm_out[MADDR][30] , \spm_out[MADDR][29] , 
        \spm_out[MADDR][28] , \spm_out[MADDR][27] , \spm_out[MADDR][26] , 
        \spm_out[MADDR][25] , \spm_out[MADDR][24] , \spm_out[MADDR][23] , 
        \spm_out[MADDR][22] , \spm_out[MADDR][21] , \spm_out[MADDR][20] , 
        \spm_out[MADDR][19] , \spm_out[MADDR][18] , \spm_out[MADDR][17] , 
        \spm_out[MADDR][16] , \spm_out[MADDR][15] , \spm_out[MADDR][14] , 
        \spm_out[MADDR][13] , \spm_out[MADDR][12] , \spm_out[MADDR][11] , 
        \spm_out[MADDR][10] , \spm_out[MADDR][9] , \spm_out[MADDR][8] , 
        \spm_out[MADDR][7] , \spm_out[MADDR][6] , \spm_out[MADDR][5] , 
        \spm_out[MADDR][4] , \spm_out[MADDR][3] , \spm_out[MADDR][2] , 
        \spm_out[MADDR][1] , \spm_out[MADDR][0] , \spm_out[MDATA][63] , 
        \spm_out[MDATA][62] , \spm_out[MDATA][61] , \spm_out[MDATA][60] , 
        \spm_out[MDATA][59] , \spm_out[MDATA][58] , \spm_out[MDATA][57] , 
        \spm_out[MDATA][56] , \spm_out[MDATA][55] , \spm_out[MDATA][54] , 
        \spm_out[MDATA][53] , \spm_out[MDATA][52] , \spm_out[MDATA][51] , 
        \spm_out[MDATA][50] , \spm_out[MDATA][49] , \spm_out[MDATA][48] , 
        \spm_out[MDATA][47] , \spm_out[MDATA][46] , \spm_out[MDATA][45] , 
        \spm_out[MDATA][44] , \spm_out[MDATA][43] , \spm_out[MDATA][42] , 
        \spm_out[MDATA][41] , \spm_out[MDATA][40] , \spm_out[MDATA][39] , 
        \spm_out[MDATA][38] , \spm_out[MDATA][37] , \spm_out[MDATA][36] , 
        \spm_out[MDATA][35] , \spm_out[MDATA][34] , \spm_out[MDATA][33] , 
        \spm_out[MDATA][32] , \spm_out[MDATA][31] , \spm_out[MDATA][30] , 
        \spm_out[MDATA][29] , \spm_out[MDATA][28] , \spm_out[MDATA][27] , 
        \spm_out[MDATA][26] , \spm_out[MDATA][25] , \spm_out[MDATA][24] , 
        \spm_out[MDATA][23] , \spm_out[MDATA][22] , \spm_out[MDATA][21] , 
        \spm_out[MDATA][20] , \spm_out[MDATA][19] , \spm_out[MDATA][18] , 
        \spm_out[MDATA][17] , \spm_out[MDATA][16] , \spm_out[MDATA][15] , 
        \spm_out[MDATA][14] , \spm_out[MDATA][13] , \spm_out[MDATA][12] , 
        \spm_out[MDATA][11] , \spm_out[MDATA][10] , \spm_out[MDATA][9] , 
        \spm_out[MDATA][8] , \spm_out[MDATA][7] , \spm_out[MDATA][6] , 
        \spm_out[MDATA][5] , \spm_out[MDATA][4] , \spm_out[MDATA][3] , 
        \spm_out[MDATA][2] , \spm_out[MDATA][1] , \spm_out[MDATA][0] }), 
        pkt_in, pkt_out );
  input [34:0] pkt_in;
  output [34:0] pkt_out;
  input na_clk, na_reset, \proc_in[MCMD][1] , \proc_in[MCMD][0] ,
         \proc_in[MADDR][31] , \proc_in[MADDR][30] , \proc_in[MADDR][29] ,
         \proc_in[MADDR][28] , \proc_in[MADDR][27] , \proc_in[MADDR][26] ,
         \proc_in[MADDR][25] , \proc_in[MADDR][24] , \proc_in[MADDR][23] ,
         \proc_in[MADDR][22] , \proc_in[MADDR][21] , \proc_in[MADDR][20] ,
         \proc_in[MADDR][19] , \proc_in[MADDR][18] , \proc_in[MADDR][17] ,
         \proc_in[MADDR][16] , \proc_in[MADDR][15] , \proc_in[MADDR][14] ,
         \proc_in[MADDR][13] , \proc_in[MADDR][12] , \proc_in[MADDR][11] ,
         \proc_in[MADDR][10] , \proc_in[MADDR][9] , \proc_in[MADDR][8] ,
         \proc_in[MADDR][7] , \proc_in[MADDR][6] , \proc_in[MADDR][5] ,
         \proc_in[MADDR][4] , \proc_in[MADDR][3] , \proc_in[MADDR][2] ,
         \proc_in[MADDR][1] , \proc_in[MADDR][0] , \proc_in[MDATA][31] ,
         \proc_in[MDATA][30] , \proc_in[MDATA][29] , \proc_in[MDATA][28] ,
         \proc_in[MDATA][27] , \proc_in[MDATA][26] , \proc_in[MDATA][25] ,
         \proc_in[MDATA][24] , \proc_in[MDATA][23] , \proc_in[MDATA][22] ,
         \proc_in[MDATA][21] , \proc_in[MDATA][20] , \proc_in[MDATA][19] ,
         \proc_in[MDATA][18] , \proc_in[MDATA][17] , \proc_in[MDATA][16] ,
         \proc_in[MDATA][15] , \proc_in[MDATA][14] , \proc_in[MDATA][13] ,
         \proc_in[MDATA][12] , \proc_in[MDATA][11] , \proc_in[MDATA][10] ,
         \proc_in[MDATA][9] , \proc_in[MDATA][8] , \proc_in[MDATA][7] ,
         \proc_in[MDATA][6] , \proc_in[MDATA][5] , \proc_in[MDATA][4] ,
         \proc_in[MDATA][3] , \proc_in[MDATA][2] , \proc_in[MDATA][1] ,
         \proc_in[MDATA][0] , \spm_in[SCMDACCEPT] , \spm_in[SRESP] ,
         \spm_in[SDATA][63] , \spm_in[SDATA][62] , \spm_in[SDATA][61] ,
         \spm_in[SDATA][60] , \spm_in[SDATA][59] , \spm_in[SDATA][58] ,
         \spm_in[SDATA][57] , \spm_in[SDATA][56] , \spm_in[SDATA][55] ,
         \spm_in[SDATA][54] , \spm_in[SDATA][53] , \spm_in[SDATA][52] ,
         \spm_in[SDATA][51] , \spm_in[SDATA][50] , \spm_in[SDATA][49] ,
         \spm_in[SDATA][48] , \spm_in[SDATA][47] , \spm_in[SDATA][46] ,
         \spm_in[SDATA][45] , \spm_in[SDATA][44] , \spm_in[SDATA][43] ,
         \spm_in[SDATA][42] , \spm_in[SDATA][41] , \spm_in[SDATA][40] ,
         \spm_in[SDATA][39] , \spm_in[SDATA][38] , \spm_in[SDATA][37] ,
         \spm_in[SDATA][36] , \spm_in[SDATA][35] , \spm_in[SDATA][34] ,
         \spm_in[SDATA][33] , \spm_in[SDATA][32] , \spm_in[SDATA][31] ,
         \spm_in[SDATA][30] , \spm_in[SDATA][29] , \spm_in[SDATA][28] ,
         \spm_in[SDATA][27] , \spm_in[SDATA][26] , \spm_in[SDATA][25] ,
         \spm_in[SDATA][24] , \spm_in[SDATA][23] , \spm_in[SDATA][22] ,
         \spm_in[SDATA][21] , \spm_in[SDATA][20] , \spm_in[SDATA][19] ,
         \spm_in[SDATA][18] , \spm_in[SDATA][17] , \spm_in[SDATA][16] ,
         \spm_in[SDATA][15] , \spm_in[SDATA][14] , \spm_in[SDATA][13] ,
         \spm_in[SDATA][12] , \spm_in[SDATA][11] , \spm_in[SDATA][10] ,
         \spm_in[SDATA][9] , \spm_in[SDATA][8] , \spm_in[SDATA][7] ,
         \spm_in[SDATA][6] , \spm_in[SDATA][5] , \spm_in[SDATA][4] ,
         \spm_in[SDATA][3] , \spm_in[SDATA][2] , \spm_in[SDATA][1] ,
         \spm_in[SDATA][0] ;
  output \proc_out[SCMDACCEPT] , \proc_out[SRESP] , \proc_out[SDATA][31] ,
         \proc_out[SDATA][30] , \proc_out[SDATA][29] , \proc_out[SDATA][28] ,
         \proc_out[SDATA][27] , \proc_out[SDATA][26] , \proc_out[SDATA][25] ,
         \proc_out[SDATA][24] , \proc_out[SDATA][23] , \proc_out[SDATA][22] ,
         \proc_out[SDATA][21] , \proc_out[SDATA][20] , \proc_out[SDATA][19] ,
         \proc_out[SDATA][18] , \proc_out[SDATA][17] , \proc_out[SDATA][16] ,
         \proc_out[SDATA][15] , \proc_out[SDATA][14] , \proc_out[SDATA][13] ,
         \proc_out[SDATA][12] , \proc_out[SDATA][11] , \proc_out[SDATA][10] ,
         \proc_out[SDATA][9] , \proc_out[SDATA][8] , \proc_out[SDATA][7] ,
         \proc_out[SDATA][6] , \proc_out[SDATA][5] , \proc_out[SDATA][4] ,
         \proc_out[SDATA][3] , \proc_out[SDATA][2] , \proc_out[SDATA][1] ,
         \proc_out[SDATA][0] , \spm_out[MCMD][1] , \spm_out[MCMD][0] ,
         \spm_out[MADDR][31] , \spm_out[MADDR][30] , \spm_out[MADDR][29] ,
         \spm_out[MADDR][28] , \spm_out[MADDR][27] , \spm_out[MADDR][26] ,
         \spm_out[MADDR][25] , \spm_out[MADDR][24] , \spm_out[MADDR][23] ,
         \spm_out[MADDR][22] , \spm_out[MADDR][21] , \spm_out[MADDR][20] ,
         \spm_out[MADDR][19] , \spm_out[MADDR][18] , \spm_out[MADDR][17] ,
         \spm_out[MADDR][16] , \spm_out[MADDR][15] , \spm_out[MADDR][14] ,
         \spm_out[MADDR][13] , \spm_out[MADDR][12] , \spm_out[MADDR][11] ,
         \spm_out[MADDR][10] , \spm_out[MADDR][9] , \spm_out[MADDR][8] ,
         \spm_out[MADDR][7] , \spm_out[MADDR][6] , \spm_out[MADDR][5] ,
         \spm_out[MADDR][4] , \spm_out[MADDR][3] , \spm_out[MADDR][2] ,
         \spm_out[MADDR][1] , \spm_out[MADDR][0] , \spm_out[MDATA][63] ,
         \spm_out[MDATA][62] , \spm_out[MDATA][61] , \spm_out[MDATA][60] ,
         \spm_out[MDATA][59] , \spm_out[MDATA][58] , \spm_out[MDATA][57] ,
         \spm_out[MDATA][56] , \spm_out[MDATA][55] , \spm_out[MDATA][54] ,
         \spm_out[MDATA][53] , \spm_out[MDATA][52] , \spm_out[MDATA][51] ,
         \spm_out[MDATA][50] , \spm_out[MDATA][49] , \spm_out[MDATA][48] ,
         \spm_out[MDATA][47] , \spm_out[MDATA][46] , \spm_out[MDATA][45] ,
         \spm_out[MDATA][44] , \spm_out[MDATA][43] , \spm_out[MDATA][42] ,
         \spm_out[MDATA][41] , \spm_out[MDATA][40] , \spm_out[MDATA][39] ,
         \spm_out[MDATA][38] , \spm_out[MDATA][37] , \spm_out[MDATA][36] ,
         \spm_out[MDATA][35] , \spm_out[MDATA][34] , \spm_out[MDATA][33] ,
         \spm_out[MDATA][32] , \spm_out[MDATA][31] , \spm_out[MDATA][30] ,
         \spm_out[MDATA][29] , \spm_out[MDATA][28] , \spm_out[MDATA][27] ,
         \spm_out[MDATA][26] , \spm_out[MDATA][25] , \spm_out[MDATA][24] ,
         \spm_out[MDATA][23] , \spm_out[MDATA][22] , \spm_out[MDATA][21] ,
         \spm_out[MDATA][20] , \spm_out[MDATA][19] , \spm_out[MDATA][18] ,
         \spm_out[MDATA][17] , \spm_out[MDATA][16] , \spm_out[MDATA][15] ,
         \spm_out[MDATA][14] , \spm_out[MDATA][13] , \spm_out[MDATA][12] ,
         \spm_out[MDATA][11] , \spm_out[MDATA][10] , \spm_out[MDATA][9] ,
         \spm_out[MDATA][8] , \spm_out[MDATA][7] , \spm_out[MDATA][6] ,
         \spm_out[MDATA][5] , \spm_out[MDATA][4] , \spm_out[MDATA][3] ,
         \spm_out[MDATA][2] , \spm_out[MDATA][1] , \spm_out[MDATA][0] ;
  wire   \spm_out[MCMD][0] , \phase_prev[0] , \phase_next[1] , vld_pkt,
         \add_545/A[8] , \add_545/A[9] , \add_545/A[10] , \add_545/A[11] ,
         \add_545/A[12] , \add_545/A[13] , \add_545/A[14] , \add_545/A[15] ,
         \sub_544/A[1] , \sub_544/A[2] , \sub_544/A[3] , \sub_544/A[4] ,
         \sub_544/A[5] , \sub_544/A[6] , \sub_544/A[7] , \sub_544/A[8] ,
         \sub_544/A[9] , \sub_544/A[10] , \sub_544/A[11] , \sub_544/A[12] , n1,
         n2, n3, n4, n5, n6, n15, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n34, n35, n37, n39, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n62, n64, n72, n73, n74, n75, n77, n78, n79, n80, n84, n87,
         n88, n89, n90, n91, n93, n94, n95, n101, n102, n103, n104, n105, n106,
         n108, n109, n111, n112, n113, n114, n116, n117, n118, n120, n122,
         n124, n125, n127, n128, n129, n130, n132, n133, n134, n136, n137,
         n138, n139, n140, n142, n144, n149, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n310, n311,
         n312, n313, n314, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883;
  wire   [2:0] slt_index;
  wire   [2:0] dma_ren;
  wire   [2:0] dma_wen;
  wire   [1:0] dma_waddr;
  wire   [63:0] dma_wdata;
  wire   [1:0] dma_raddr;
  wire   [63:0] dma_rdata;
  wire   [4:0] slt_entry;
  wire   [1:0] state_cnt;
  wire   [4:0] config_reg;
  wire   [70:64] flit_buf;
  wire   [34:0] phitIn;
  wire   [31:0] mux_out;
  wire   [31:0] dOut_l;
  wire   [34:32] phit_togo;
  wire   [34:0] phitOut0;
  wire   [34:0] phitOut1;
  wire   [34:0] phitOut2;
  wire   [13:0] dma_cnt_new;
  wire   [15:0] dma_rp_new;
  wire   [15:0] dma_wp_new;
  wire   [6:0] address;
  wire   [31:0] dIn_h;
  assign \spm_out[MADDR][15]  = 1'b0;
  assign \spm_out[MADDR][16]  = 1'b0;
  assign \spm_out[MADDR][17]  = 1'b0;
  assign \spm_out[MADDR][18]  = 1'b0;
  assign \spm_out[MADDR][19]  = 1'b0;
  assign \spm_out[MADDR][20]  = 1'b0;
  assign \spm_out[MADDR][21]  = 1'b0;
  assign \spm_out[MADDR][22]  = 1'b0;
  assign \spm_out[MADDR][23]  = 1'b0;
  assign \spm_out[MADDR][24]  = 1'b0;
  assign \spm_out[MADDR][25]  = 1'b0;
  assign \spm_out[MADDR][26]  = 1'b0;
  assign \spm_out[MADDR][27]  = 1'b0;
  assign \spm_out[MADDR][28]  = 1'b0;
  assign \spm_out[MADDR][29]  = 1'b0;
  assign \spm_out[MADDR][30]  = 1'b0;
  assign \spm_out[MADDR][31]  = 1'b0;
  assign \spm_out[MCMD][1]  = \spm_out[MCMD][0] ;

  HS65_LS_DFPRQX9 \phase_next_reg[1]  ( .D(n681), .CP(na_clk), .RN(n348), .Q(
        \phase_next[1] ) );
  HS65_LS_DFPRQX9 \dOut_l_reg[31]  ( .D(n691), .CP(na_clk), .RN(n352), .Q(
        dOut_l[31]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[30]  ( .D(n692), .CP(na_clk), .RN(n350), .Q(
        dOut_l[30]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[29]  ( .D(n693), .CP(na_clk), .RN(n348), .Q(
        dOut_l[29]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[28]  ( .D(n694), .CP(na_clk), .RN(n346), .Q(
        dOut_l[28]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[27]  ( .D(n695), .CP(na_clk), .RN(n351), .Q(
        dOut_l[27]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[26]  ( .D(n696), .CP(na_clk), .RN(n341), .Q(
        dOut_l[26]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[25]  ( .D(n697), .CP(na_clk), .RN(n354), .Q(
        dOut_l[25]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[24]  ( .D(n698), .CP(na_clk), .RN(n353), .Q(
        dOut_l[24]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[23]  ( .D(n699), .CP(na_clk), .RN(n349), .Q(
        dOut_l[23]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[22]  ( .D(n700), .CP(na_clk), .RN(n347), .Q(
        dOut_l[22]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[21]  ( .D(n701), .CP(na_clk), .RN(n346), .Q(
        dOut_l[21]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[20]  ( .D(n702), .CP(na_clk), .RN(n344), .Q(
        dOut_l[20]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[19]  ( .D(n703), .CP(na_clk), .RN(n343), .Q(
        dOut_l[19]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[18]  ( .D(n704), .CP(na_clk), .RN(n342), .Q(
        dOut_l[18]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[17]  ( .D(n705), .CP(na_clk), .RN(n344), .Q(
        dOut_l[17]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[16]  ( .D(n706), .CP(na_clk), .RN(n343), .Q(
        dOut_l[16]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[15]  ( .D(n707), .CP(na_clk), .RN(n342), .Q(
        dOut_l[15]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[14]  ( .D(n708), .CP(na_clk), .RN(n345), .Q(
        dOut_l[14]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[13]  ( .D(n709), .CP(na_clk), .RN(n355), .Q(
        dOut_l[13]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[12]  ( .D(n710), .CP(na_clk), .RN(n351), .Q(
        dOut_l[12]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[11]  ( .D(n711), .CP(na_clk), .RN(n341), .Q(
        dOut_l[11]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[10]  ( .D(n712), .CP(na_clk), .RN(n354), .Q(
        dOut_l[10]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[9]  ( .D(n713), .CP(na_clk), .RN(n353), .Q(
        dOut_l[9]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[8]  ( .D(n714), .CP(na_clk), .RN(n349), .Q(
        dOut_l[8]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[7]  ( .D(n715), .CP(na_clk), .RN(n347), .Q(
        dOut_l[7]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[6]  ( .D(n716), .CP(na_clk), .RN(n346), .Q(
        dOut_l[6]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[5]  ( .D(n717), .CP(na_clk), .RN(n344), .Q(
        dOut_l[5]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[4]  ( .D(n718), .CP(na_clk), .RN(n343), .Q(
        dOut_l[4]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[3]  ( .D(n719), .CP(na_clk), .RN(n342), .Q(
        dOut_l[3]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[2]  ( .D(n720), .CP(na_clk), .RN(n345), .Q(
        dOut_l[2]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[1]  ( .D(n721), .CP(na_clk), .RN(n355), .Q(
        dOut_l[1]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[0]  ( .D(n722), .CP(na_clk), .RN(n348), .Q(
        dOut_l[0]) );
  HS65_LS_DFPRQX9 \phitIn_reg[34]  ( .D(pkt_in[34]), .CP(na_clk), .RN(n342), 
        .Q(phitIn[34]) );
  HS65_LS_DFPRQX9 \phitIn_reg[33]  ( .D(pkt_in[33]), .CP(na_clk), .RN(n343), 
        .Q(phitIn[33]) );
  HS65_LS_DFPRQX9 vld_pkt_reg ( .D(n684), .CP(na_clk), .RN(n344), .Q(vld_pkt)
         );
  HS65_LS_DFPRQX9 \phitIn_reg[32]  ( .D(pkt_in[32]), .CP(na_clk), .RN(n346), 
        .Q(phitIn[32]) );
  HS65_LS_DFPRQX9 \phitIn_reg[31]  ( .D(pkt_in[31]), .CP(na_clk), .RN(n347), 
        .Q(phitIn[31]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[31]  ( .D(n723), .CP(na_clk), .RN(n349), .Q(
        dIn_h[31]) );
  HS65_LS_DFPRQX9 \phitIn_reg[30]  ( .D(pkt_in[30]), .CP(na_clk), .RN(n353), 
        .Q(phitIn[30]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[30]  ( .D(n724), .CP(na_clk), .RN(n354), .Q(
        dIn_h[30]) );
  HS65_LS_DFPRQX9 \phitIn_reg[29]  ( .D(pkt_in[29]), .CP(na_clk), .RN(n341), 
        .Q(phitIn[29]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[29]  ( .D(n725), .CP(na_clk), .RN(n351), .Q(
        dIn_h[29]) );
  HS65_LS_DFPRQX9 \phitIn_reg[28]  ( .D(pkt_in[28]), .CP(na_clk), .RN(n350), 
        .Q(phitIn[28]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[28]  ( .D(n726), .CP(na_clk), .RN(n352), .Q(
        dIn_h[28]) );
  HS65_LS_DFPRQX9 \phitIn_reg[27]  ( .D(pkt_in[27]), .CP(na_clk), .RN(n350), 
        .Q(phitIn[27]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[27]  ( .D(n727), .CP(na_clk), .RN(n350), .Q(
        dIn_h[27]) );
  HS65_LS_DFPRQX9 \phitIn_reg[26]  ( .D(pkt_in[26]), .CP(na_clk), .RN(n350), 
        .Q(phitIn[26]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[26]  ( .D(n728), .CP(na_clk), .RN(n350), .Q(
        dIn_h[26]) );
  HS65_LS_DFPRQX9 \phitIn_reg[25]  ( .D(pkt_in[25]), .CP(na_clk), .RN(n350), 
        .Q(phitIn[25]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[25]  ( .D(n729), .CP(na_clk), .RN(n350), .Q(
        dIn_h[25]) );
  HS65_LS_DFPRQX9 \phitIn_reg[24]  ( .D(pkt_in[24]), .CP(na_clk), .RN(n350), 
        .Q(phitIn[24]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[24]  ( .D(n730), .CP(na_clk), .RN(n350), .Q(
        dIn_h[24]) );
  HS65_LS_DFPRQX9 \phitIn_reg[23]  ( .D(pkt_in[23]), .CP(na_clk), .RN(n350), 
        .Q(phitIn[23]) );
  HS65_LS_DFPRQX9 \address_reg[6]  ( .D(n731), .CP(na_clk), .RN(n350), .Q(
        address[6]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[23]  ( .D(n732), .CP(na_clk), .RN(n350), .Q(
        dIn_h[23]) );
  HS65_LS_DFPRQX9 \phitIn_reg[22]  ( .D(pkt_in[22]), .CP(na_clk), .RN(n350), 
        .Q(phitIn[22]) );
  HS65_LS_DFPRQX9 \address_reg[5]  ( .D(n733), .CP(na_clk), .RN(n350), .Q(
        address[5]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[22]  ( .D(n734), .CP(na_clk), .RN(n350), .Q(
        dIn_h[22]) );
  HS65_LS_DFPRQX9 \phitIn_reg[21]  ( .D(pkt_in[21]), .CP(na_clk), .RN(n350), 
        .Q(phitIn[21]) );
  HS65_LS_DFPRQX9 \address_reg[4]  ( .D(n735), .CP(na_clk), .RN(n351), .Q(
        address[4]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[21]  ( .D(n736), .CP(na_clk), .RN(n351), .Q(
        dIn_h[21]) );
  HS65_LS_DFPRQX9 \phitIn_reg[20]  ( .D(pkt_in[20]), .CP(na_clk), .RN(n351), 
        .Q(phitIn[20]) );
  HS65_LS_DFPRQX9 \address_reg[3]  ( .D(n737), .CP(na_clk), .RN(n351), .Q(
        address[3]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[20]  ( .D(n738), .CP(na_clk), .RN(n351), .Q(
        dIn_h[20]) );
  HS65_LS_DFPRQX9 \phitIn_reg[19]  ( .D(pkt_in[19]), .CP(na_clk), .RN(n351), 
        .Q(phitIn[19]) );
  HS65_LS_DFPRQX9 \address_reg[2]  ( .D(n739), .CP(na_clk), .RN(n351), .Q(
        address[2]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[19]  ( .D(n740), .CP(na_clk), .RN(n351), .Q(
        dIn_h[19]) );
  HS65_LS_DFPRQX9 \phitIn_reg[18]  ( .D(pkt_in[18]), .CP(na_clk), .RN(n351), 
        .Q(phitIn[18]) );
  HS65_LS_DFPRQX9 \address_reg[1]  ( .D(n741), .CP(na_clk), .RN(n351), .Q(
        address[1]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[18]  ( .D(n742), .CP(na_clk), .RN(n351), .Q(
        dIn_h[18]) );
  HS65_LS_DFPRQX9 \phitIn_reg[17]  ( .D(pkt_in[17]), .CP(na_clk), .RN(n351), 
        .Q(phitIn[17]) );
  HS65_LS_DFPRQX9 \address_reg[0]  ( .D(n743), .CP(na_clk), .RN(n351), .Q(
        address[0]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[17]  ( .D(n744), .CP(na_clk), .RN(n351), .Q(
        dIn_h[17]) );
  HS65_LS_DFPRQX9 \phitIn_reg[16]  ( .D(pkt_in[16]), .CP(na_clk), .RN(n352), 
        .Q(phitIn[16]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[16]  ( .D(n745), .CP(na_clk), .RN(n352), .Q(
        dIn_h[16]) );
  HS65_LS_DFPRQX9 \phitIn_reg[15]  ( .D(pkt_in[15]), .CP(na_clk), .RN(n352), 
        .Q(phitIn[15]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[15]  ( .D(n746), .CP(na_clk), .RN(n352), .Q(
        dIn_h[15]) );
  HS65_LS_DFPRQX9 \phitIn_reg[14]  ( .D(pkt_in[14]), .CP(na_clk), .RN(n352), 
        .Q(phitIn[14]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[14]  ( .D(n747), .CP(na_clk), .RN(n352), .Q(
        dIn_h[14]) );
  HS65_LS_DFPRQX9 \phitIn_reg[13]  ( .D(pkt_in[13]), .CP(na_clk), .RN(n352), 
        .Q(phitIn[13]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[13]  ( .D(n748), .CP(na_clk), .RN(n352), .Q(
        dIn_h[13]) );
  HS65_LS_DFPRQX9 \phitIn_reg[12]  ( .D(pkt_in[12]), .CP(na_clk), .RN(n352), 
        .Q(phitIn[12]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[12]  ( .D(n749), .CP(na_clk), .RN(n352), .Q(
        dIn_h[12]) );
  HS65_LS_DFPRQX9 \phitIn_reg[11]  ( .D(pkt_in[11]), .CP(na_clk), .RN(n352), 
        .Q(phitIn[11]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[11]  ( .D(n750), .CP(na_clk), .RN(n352), .Q(
        dIn_h[11]) );
  HS65_LS_DFPRQX9 \phitIn_reg[10]  ( .D(pkt_in[10]), .CP(na_clk), .RN(n352), 
        .Q(phitIn[10]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[10]  ( .D(n751), .CP(na_clk), .RN(n352), .Q(
        dIn_h[10]) );
  HS65_LS_DFPRQX9 \phitIn_reg[9]  ( .D(pkt_in[9]), .CP(na_clk), .RN(n352), .Q(
        phitIn[9]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[9]  ( .D(n752), .CP(na_clk), .RN(n353), .Q(
        dIn_h[9]) );
  HS65_LS_DFPRQX9 \phitIn_reg[8]  ( .D(pkt_in[8]), .CP(na_clk), .RN(n353), .Q(
        phitIn[8]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[8]  ( .D(n753), .CP(na_clk), .RN(n353), .Q(
        dIn_h[8]) );
  HS65_LS_DFPRQX9 \phitIn_reg[7]  ( .D(pkt_in[7]), .CP(na_clk), .RN(n353), .Q(
        phitIn[7]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[7]  ( .D(n754), .CP(na_clk), .RN(n353), .Q(
        dIn_h[7]) );
  HS65_LS_DFPRQX9 \phitIn_reg[6]  ( .D(pkt_in[6]), .CP(na_clk), .RN(n353), .Q(
        phitIn[6]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[6]  ( .D(n755), .CP(na_clk), .RN(n353), .Q(
        dIn_h[6]) );
  HS65_LS_DFPRQX9 \phitIn_reg[5]  ( .D(pkt_in[5]), .CP(na_clk), .RN(n353), .Q(
        phitIn[5]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[5]  ( .D(n756), .CP(na_clk), .RN(n353), .Q(
        dIn_h[5]) );
  HS65_LS_DFPRQX9 \phitIn_reg[4]  ( .D(pkt_in[4]), .CP(na_clk), .RN(n353), .Q(
        phitIn[4]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[4]  ( .D(n757), .CP(na_clk), .RN(n353), .Q(
        dIn_h[4]) );
  HS65_LS_DFPRQX9 \phitIn_reg[3]  ( .D(pkt_in[3]), .CP(na_clk), .RN(n353), .Q(
        phitIn[3]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[3]  ( .D(n758), .CP(na_clk), .RN(n353), .Q(
        dIn_h[3]) );
  HS65_LS_DFPRQX9 \phitIn_reg[2]  ( .D(pkt_in[2]), .CP(na_clk), .RN(n353), .Q(
        phitIn[2]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[2]  ( .D(n759), .CP(na_clk), .RN(n353), .Q(
        dIn_h[2]) );
  HS65_LS_DFPRQX9 \phitIn_reg[1]  ( .D(pkt_in[1]), .CP(na_clk), .RN(n354), .Q(
        phitIn[1]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[1]  ( .D(n760), .CP(na_clk), .RN(n354), .Q(
        dIn_h[1]) );
  HS65_LS_DFPRQX9 \phitIn_reg[0]  ( .D(pkt_in[0]), .CP(na_clk), .RN(n354), .Q(
        phitIn[0]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[0]  ( .D(n761), .CP(na_clk), .RN(n354), .Q(
        dIn_h[0]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[34]  ( .D(phit_togo[34]), .CP(na_clk), .RN(
        n354), .Q(phitOut0[34]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[33]  ( .D(n333), .CP(na_clk), .RN(n354), .Q(
        phitOut0[33]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[32]  ( .D(phit_togo[32]), .CP(na_clk), .RN(
        n354), .Q(phitOut0[32]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[31]  ( .D(mux_out[31]), .CP(na_clk), .RN(n354), 
        .Q(phitOut0[31]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[30]  ( .D(mux_out[30]), .CP(na_clk), .RN(n354), 
        .Q(phitOut0[30]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[29]  ( .D(mux_out[29]), .CP(na_clk), .RN(n354), 
        .Q(phitOut0[29]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[28]  ( .D(mux_out[28]), .CP(na_clk), .RN(n354), 
        .Q(phitOut0[28]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[27]  ( .D(mux_out[27]), .CP(na_clk), .RN(n354), 
        .Q(phitOut0[27]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[26]  ( .D(mux_out[26]), .CP(na_clk), .RN(n354), 
        .Q(phitOut0[26]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[25]  ( .D(mux_out[25]), .CP(na_clk), .RN(n354), 
        .Q(phitOut0[25]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[24]  ( .D(mux_out[24]), .CP(na_clk), .RN(n354), 
        .Q(phitOut0[24]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[23]  ( .D(mux_out[23]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[23]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[22]  ( .D(mux_out[22]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[22]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[21]  ( .D(mux_out[21]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[21]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[20]  ( .D(mux_out[20]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[20]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[19]  ( .D(mux_out[19]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[19]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[18]  ( .D(mux_out[18]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[18]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[17]  ( .D(mux_out[17]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[17]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[16]  ( .D(mux_out[16]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[16]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[15]  ( .D(mux_out[15]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[15]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[14]  ( .D(mux_out[14]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[14]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[13]  ( .D(mux_out[13]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[13]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[12]  ( .D(mux_out[12]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[12]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[11]  ( .D(mux_out[11]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[11]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[10]  ( .D(mux_out[10]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[10]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[9]  ( .D(mux_out[9]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[9]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[8]  ( .D(mux_out[8]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[8]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[7]  ( .D(mux_out[7]), .CP(na_clk), .RN(n348), 
        .Q(phitOut0[7]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[6]  ( .D(mux_out[6]), .CP(na_clk), .RN(n345), 
        .Q(phitOut0[6]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[5]  ( .D(mux_out[5]), .CP(na_clk), .RN(n342), 
        .Q(phitOut0[5]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[4]  ( .D(mux_out[4]), .CP(na_clk), .RN(n343), 
        .Q(phitOut0[4]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[3]  ( .D(mux_out[3]), .CP(na_clk), .RN(n344), 
        .Q(phitOut0[3]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[2]  ( .D(mux_out[2]), .CP(na_clk), .RN(n346), 
        .Q(phitOut0[2]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[1]  ( .D(mux_out[1]), .CP(na_clk), .RN(n347), 
        .Q(phitOut0[1]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[0]  ( .D(mux_out[0]), .CP(na_clk), .RN(n341), 
        .Q(phitOut0[0]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[34]  ( .D(phitOut0[34]), .CP(na_clk), .RN(n345), .Q(phitOut1[34]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[33]  ( .D(phitOut0[33]), .CP(na_clk), .RN(n341), .Q(phitOut1[33]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[32]  ( .D(phitOut0[32]), .CP(na_clk), .RN(n341), .Q(phitOut1[32]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[31]  ( .D(phitOut0[31]), .CP(na_clk), .RN(n341), .Q(phitOut1[31]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[30]  ( .D(phitOut0[30]), .CP(na_clk), .RN(n341), .Q(phitOut1[30]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[29]  ( .D(phitOut0[29]), .CP(na_clk), .RN(n341), .Q(phitOut1[29]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[28]  ( .D(phitOut0[28]), .CP(na_clk), .RN(n341), .Q(phitOut1[28]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[27]  ( .D(phitOut0[27]), .CP(na_clk), .RN(n341), .Q(phitOut1[27]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[26]  ( .D(phitOut0[26]), .CP(na_clk), .RN(n341), .Q(phitOut1[26]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[25]  ( .D(phitOut0[25]), .CP(na_clk), .RN(n341), .Q(phitOut1[25]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[24]  ( .D(phitOut0[24]), .CP(na_clk), .RN(n341), .Q(phitOut1[24]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[23]  ( .D(phitOut0[23]), .CP(na_clk), .RN(n341), .Q(phitOut1[23]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[22]  ( .D(phitOut0[22]), .CP(na_clk), .RN(n341), .Q(phitOut1[22]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[21]  ( .D(phitOut0[21]), .CP(na_clk), .RN(n355), .Q(phitOut1[21]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[20]  ( .D(phitOut0[20]), .CP(na_clk), .RN(n350), .Q(phitOut1[20]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[19]  ( .D(phitOut0[19]), .CP(na_clk), .RN(n352), .Q(phitOut1[19]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[18]  ( .D(phitOut0[18]), .CP(na_clk), .RN(n348), .Q(phitOut1[18]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[17]  ( .D(phitOut0[17]), .CP(na_clk), .RN(n353), .Q(phitOut1[17]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[16]  ( .D(phitOut0[16]), .CP(na_clk), .RN(n354), .Q(phitOut1[16]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[15]  ( .D(phitOut0[15]), .CP(na_clk), .RN(n349), .Q(phitOut1[15]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[14]  ( .D(phitOut0[14]), .CP(na_clk), .RN(n341), .Q(phitOut1[14]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[13]  ( .D(phitOut0[13]), .CP(na_clk), .RN(n345), .Q(phitOut1[13]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[12]  ( .D(phitOut0[12]), .CP(na_clk), .RN(n355), .Q(phitOut1[12]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[11]  ( .D(phitOut0[11]), .CP(na_clk), .RN(n351), .Q(phitOut1[11]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[10]  ( .D(phitOut0[10]), .CP(na_clk), .RN(n347), .Q(phitOut1[10]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[9]  ( .D(phitOut0[9]), .CP(na_clk), .RN(n345), 
        .Q(phitOut1[9]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[8]  ( .D(phitOut0[8]), .CP(na_clk), .RN(n350), 
        .Q(phitOut1[8]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[7]  ( .D(phitOut0[7]), .CP(na_clk), .RN(n352), 
        .Q(phitOut1[7]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[6]  ( .D(phitOut0[6]), .CP(na_clk), .RN(n342), 
        .Q(phitOut1[6]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[5]  ( .D(phitOut0[5]), .CP(na_clk), .RN(n342), 
        .Q(phitOut1[5]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[4]  ( .D(phitOut0[4]), .CP(na_clk), .RN(n342), 
        .Q(phitOut1[4]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[3]  ( .D(phitOut0[3]), .CP(na_clk), .RN(n342), 
        .Q(phitOut1[3]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[2]  ( .D(phitOut0[2]), .CP(na_clk), .RN(n342), 
        .Q(phitOut1[2]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[1]  ( .D(phitOut0[1]), .CP(na_clk), .RN(n342), 
        .Q(phitOut1[1]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[0]  ( .D(phitOut0[0]), .CP(na_clk), .RN(n342), 
        .Q(phitOut1[0]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[34]  ( .D(phitOut1[34]), .CP(na_clk), .RN(n342), .Q(phitOut2[34]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[33]  ( .D(phitOut1[33]), .CP(na_clk), .RN(n342), .Q(phitOut2[33]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[32]  ( .D(phitOut1[32]), .CP(na_clk), .RN(n342), .Q(phitOut2[32]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[31]  ( .D(phitOut1[31]), .CP(na_clk), .RN(n342), .Q(phitOut2[31]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[30]  ( .D(phitOut1[30]), .CP(na_clk), .RN(n342), .Q(phitOut2[30]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[29]  ( .D(phitOut1[29]), .CP(na_clk), .RN(n342), .Q(phitOut2[29]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[28]  ( .D(phitOut1[28]), .CP(na_clk), .RN(n342), .Q(phitOut2[28]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[27]  ( .D(phitOut1[27]), .CP(na_clk), .RN(n342), .Q(phitOut2[27]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[26]  ( .D(phitOut1[26]), .CP(na_clk), .RN(n343), .Q(phitOut2[26]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[25]  ( .D(phitOut1[25]), .CP(na_clk), .RN(n343), .Q(phitOut2[25]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[24]  ( .D(phitOut1[24]), .CP(na_clk), .RN(n343), .Q(phitOut2[24]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[23]  ( .D(phitOut1[23]), .CP(na_clk), .RN(n343), .Q(phitOut2[23]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[22]  ( .D(phitOut1[22]), .CP(na_clk), .RN(n343), .Q(phitOut2[22]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[21]  ( .D(phitOut1[21]), .CP(na_clk), .RN(n343), .Q(phitOut2[21]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[20]  ( .D(phitOut1[20]), .CP(na_clk), .RN(n343), .Q(phitOut2[20]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[19]  ( .D(phitOut1[19]), .CP(na_clk), .RN(n343), .Q(phitOut2[19]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[18]  ( .D(phitOut1[18]), .CP(na_clk), .RN(n343), .Q(phitOut2[18]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[17]  ( .D(phitOut1[17]), .CP(na_clk), .RN(n343), .Q(phitOut2[17]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[16]  ( .D(phitOut1[16]), .CP(na_clk), .RN(n343), .Q(phitOut2[16]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[15]  ( .D(phitOut1[15]), .CP(na_clk), .RN(n343), .Q(phitOut2[15]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[14]  ( .D(phitOut1[14]), .CP(na_clk), .RN(n343), .Q(phitOut2[14]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[13]  ( .D(phitOut1[13]), .CP(na_clk), .RN(n343), .Q(phitOut2[13]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[12]  ( .D(phitOut1[12]), .CP(na_clk), .RN(n343), .Q(phitOut2[12]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[11]  ( .D(phitOut1[11]), .CP(na_clk), .RN(n344), .Q(phitOut2[11]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[10]  ( .D(phitOut1[10]), .CP(na_clk), .RN(n344), .Q(phitOut2[10]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[9]  ( .D(phitOut1[9]), .CP(na_clk), .RN(n344), 
        .Q(phitOut2[9]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[8]  ( .D(phitOut1[8]), .CP(na_clk), .RN(n344), 
        .Q(phitOut2[8]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[7]  ( .D(phitOut1[7]), .CP(na_clk), .RN(n344), 
        .Q(phitOut2[7]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[6]  ( .D(phitOut1[6]), .CP(na_clk), .RN(n344), 
        .Q(phitOut2[6]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[5]  ( .D(phitOut1[5]), .CP(na_clk), .RN(n344), 
        .Q(phitOut2[5]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[4]  ( .D(phitOut1[4]), .CP(na_clk), .RN(n344), 
        .Q(phitOut2[4]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[3]  ( .D(phitOut1[3]), .CP(na_clk), .RN(n344), 
        .Q(phitOut2[3]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[2]  ( .D(phitOut1[2]), .CP(na_clk), .RN(n344), 
        .Q(phitOut2[2]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[1]  ( .D(phitOut1[1]), .CP(na_clk), .RN(n344), 
        .Q(phitOut2[1]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[0]  ( .D(phitOut1[0]), .CP(na_clk), .RN(n344), 
        .Q(phitOut2[0]) );
  HS65_LS_DFPRQX9 \config_reg_reg[4]  ( .D(\proc_in[MCMD][1] ), .CP(na_clk), 
        .RN(n344), .Q(config_reg[4]) );
  HS65_LS_DFPRQX9 \config_reg_reg[3]  ( .D(n680), .CP(na_clk), .RN(n344), .Q(
        config_reg[3]) );
  HS65_LS_DFPRQX9 \config_reg_reg[2]  ( .D(n657), .CP(na_clk), .RN(n344), .Q(
        config_reg[2]) );
  HS65_LS_DFPRQX9 \config_reg_reg[1]  ( .D(n658), .CP(na_clk), .RN(n345), .Q(
        config_reg[1]) );
  HS65_LS_DFPRQX9 \config_reg_reg[0]  ( .D(n656), .CP(na_clk), .RN(n345), .Q(
        config_reg[0]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[70]  ( .D(n762), .CP(na_clk), .RN(n345), .Q(
        flit_buf[70]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[69]  ( .D(n763), .CP(na_clk), .RN(n345), .Q(
        flit_buf[69]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[68]  ( .D(n764), .CP(na_clk), .RN(n345), .Q(
        flit_buf[68]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[67]  ( .D(n765), .CP(na_clk), .RN(n345), .Q(
        flit_buf[67]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[66]  ( .D(n766), .CP(na_clk), .RN(n345), .Q(
        flit_buf[66]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[65]  ( .D(n767), .CP(na_clk), .RN(n345), .Q(
        flit_buf[65]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[64]  ( .D(n768), .CP(na_clk), .RN(n345), .Q(
        flit_buf[64]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[63]  ( .D(n769), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][63] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[62]  ( .D(n770), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][62] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[61]  ( .D(n771), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][61] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[60]  ( .D(n772), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][60] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[59]  ( .D(n773), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][59] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[58]  ( .D(n774), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][58] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[57]  ( .D(n775), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][57] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[56]  ( .D(n776), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][56] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[55]  ( .D(n777), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][55] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[54]  ( .D(n778), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][54] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[53]  ( .D(n779), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][53] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[52]  ( .D(n780), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][52] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[51]  ( .D(n781), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][51] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[50]  ( .D(n782), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][50] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[49]  ( .D(n783), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][49] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[48]  ( .D(n784), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][48] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[47]  ( .D(n785), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][47] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[46]  ( .D(n786), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][46] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[45]  ( .D(n787), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][45] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[44]  ( .D(n788), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][44] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[43]  ( .D(n789), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][43] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[42]  ( .D(n790), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][42] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[41]  ( .D(n791), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][41] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[40]  ( .D(n792), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][40] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[39]  ( .D(n793), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][39] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[38]  ( .D(n794), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][38] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[37]  ( .D(n795), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][37] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[36]  ( .D(n796), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][36] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[35]  ( .D(n797), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][35] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[34]  ( .D(n798), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][34] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[33]  ( .D(n799), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][33] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[32]  ( .D(n800), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][32] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[31]  ( .D(n801), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][31] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[30]  ( .D(n802), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][30] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[29]  ( .D(n803), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][29] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[28]  ( .D(n804), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][28] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[27]  ( .D(n805), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][27] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[26]  ( .D(n806), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][26] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[25]  ( .D(n807), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][25] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[24]  ( .D(n808), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][24] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[23]  ( .D(n809), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][23] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[22]  ( .D(n810), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][22] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[21]  ( .D(n811), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][21] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[20]  ( .D(n812), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][20] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[19]  ( .D(n813), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][19] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[18]  ( .D(n814), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][18] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[17]  ( .D(n815), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][17] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[16]  ( .D(n816), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][16] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[15]  ( .D(n817), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][15] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[14]  ( .D(n818), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][14] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[13]  ( .D(n819), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][13] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[12]  ( .D(n820), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][12] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[11]  ( .D(n821), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][11] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[10]  ( .D(n822), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][10] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[9]  ( .D(n823), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][9] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[8]  ( .D(n824), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][8] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[7]  ( .D(n825), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][7] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[6]  ( .D(n826), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][6] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[5]  ( .D(n827), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][5] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[4]  ( .D(n828), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][4] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[3]  ( .D(n829), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][3] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[2]  ( .D(n830), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][2] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[1]  ( .D(n831), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][1] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[0]  ( .D(n832), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][0] ) );
  HS65_LS_DFPRQX9 \phase_prev_reg[0]  ( .D(n687), .CP(na_clk), .RN(n349), .Q(
        \phase_prev[0] ) );
  counter_WIDTH3_2 slt_cnt ( .clk(na_clk), .reset(n356), .enable(n652), .cnt(
        slt_index) );
  dma_sdp_DATA64_ADDR2_2 dma_table ( .clk(na_clk), .reset(n357), .ren(dma_ren), 
        .wen(dma_wen), .waddr(dma_waddr), .wdata(dma_wdata), .raddr(dma_raddr), 
        .rdata(dma_rdata) );
  bram_DATA5_ADDR3_2 slt_table ( .clk(na_clk), .reset(n356), .rd_addr(
        slt_index), .wr_addr({\proc_in[MADDR][2] , \proc_in[MADDR][1] , 
        \proc_in[MADDR][0] }), .wr_data({\proc_in[MDATA][4] , 
        \proc_in[MDATA][3] , \proc_in[MDATA][2] , \proc_in[MDATA][1] , 
        \proc_in[MDATA][0] }), .wr_ena(n655), .rd_data(slt_entry) );
  HS65_LS_DFPRQNX9 vld_buf_reg ( .D(n685), .CP(na_clk), .RN(n349), .QN(n688)
         );
  HS65_LS_DFPRQNX9 dma_ctrl_reg_reg ( .D(n683), .CP(na_clk), .RN(n353), .QN(
        n689) );
  HS65_LS_DFPRQX9 \state_cnt_reg[0]  ( .D(n34), .CP(na_clk), .RN(n341), .Q(
        state_cnt[0]) );
  HS65_LS_DFPRQX9 \state_cnt_reg[1]  ( .D(n602), .CP(na_clk), .RN(n351), .Q(
        state_cnt[1]) );
  HS65_LS_DFPRQNX9 \phase_next_reg[0]  ( .D(n682), .CP(na_clk), .RN(n354), 
        .QN(n690) );
  HS65_LS_DFPRQX9 \phase_prev_reg[1]  ( .D(n686), .CP(na_clk), .RN(n341), .Q(
        n23) );
  HS65_LS_IVX31 U3 ( .A(n46), .Z(n30) );
  HS65_LS_BFX31 U4 ( .A(n575), .Z(n47) );
  HS65_LS_BFX13 U5 ( .A(n32), .Z(n21) );
  HS65_LS_NAND2X14 U6 ( .A(n577), .B(n472), .Z(n31) );
  HS65_LS_OAI12X6 U7 ( .A(n6), .B(n580), .C(n579), .Z(pkt_out[34]) );
  HS65_LS_NAND2X29 U8 ( .A(n481), .B(n41), .Z(n468) );
  HS65_LS_NAND2X14 U9 ( .A(n43), .B(n479), .Z(n35) );
  HS65_LS_NAND2X11 U10 ( .A(n46), .B(phitOut0[2]), .Z(n43) );
  HS65_LS_IVX31 U11 ( .A(n472), .Z(n26) );
  HS65_LS_BFX40 U12 ( .A(n575), .Z(n48) );
  HS65_LS_NAND2X14 U13 ( .A(n577), .B(n26), .Z(n575) );
  HS65_LS_NAND2X14 U14 ( .A(n577), .B(n472), .Z(n32) );
  HS65_LS_NAND2X5 U15 ( .A(n20), .B(n467), .Z(n450) );
  HS65_LS_IVX4 U16 ( .A(n467), .Z(n456) );
  HS65_LS_NAND3X13 U17 ( .A(n139), .B(n456), .C(n455), .Z(n457) );
  HS65_LH_OAI222X2 U18 ( .A(n662), .B(n855), .C(n650), .D(n451), .E(n661), .F(
        n857), .Z(dma_waddr[1]) );
  HS65_LH_OAI222X2 U19 ( .A(n663), .B(n855), .C(n651), .D(n451), .E(n662), .F(
        n857), .Z(dma_waddr[0]) );
  HS65_LS_IVX27 U20 ( .A(n468), .Z(n577) );
  HS65_LS_AND2X4 U21 ( .A(\proc_in[MCMD][0] ), .B(n597), .Z(n1) );
  HS65_LS_IVX22 U22 ( .A(n575), .Z(n46) );
  HS65_LS_AND2X4 U23 ( .A(n616), .B(n73), .Z(n2) );
  HS65_LS_AND2X4 U24 ( .A(\add_545/A[14] ), .B(n89), .Z(n3) );
  HS65_LH_BFX4 U25 ( .A(n139), .Z(n140) );
  HS65_LS_AND2X4 U26 ( .A(n142), .B(n415), .Z(n4) );
  HS65_LS_IVX2 U27 ( .A(n44), .Z(n20) );
  HS65_LH_IVX2 U28 ( .A(n454), .Z(n5) );
  HS65_LS_NAND2X7 U29 ( .A(phitOut2[2]), .B(n101), .Z(n479) );
  HS65_LS_NAND2X5 U30 ( .A(phitOut2[1]), .B(n101), .Z(n476) );
  HS65_LS_NAND2X5 U31 ( .A(phitOut2[0]), .B(n101), .Z(n473) );
  HS65_LS_NAND2X4 U32 ( .A(phitOut2[11]), .B(n517), .Z(n506) );
  HS65_LS_NAND2X5 U33 ( .A(phitOut2[23]), .B(n25), .Z(n542) );
  HS65_LS_NAND2X5 U34 ( .A(phitOut2[27]), .B(n25), .Z(n554) );
  HS65_LS_NAND2X5 U35 ( .A(phitOut2[4]), .B(n25), .Z(n485) );
  HS65_LS_NAND2X5 U36 ( .A(phitOut2[12]), .B(n25), .Z(n508) );
  HS65_LS_IVX18 U37 ( .A(n28), .Z(n6) );
  HS65_LS_IVX22 U38 ( .A(n28), .Z(n15) );
  HS65_LS_IVX27 U39 ( .A(n28), .Z(n29) );
  HS65_LS_IVX31 U40 ( .A(n17), .Z(n25) );
  HS65_LS_NAND2X29 U41 ( .A(n471), .B(n129), .Z(n472) );
  HS65_LS_NAND2X21 U42 ( .A(n468), .B(n26), .Z(n17) );
  HS65_LS_NAND2X14 U43 ( .A(n46), .B(phitOut0[11]), .Z(n51) );
  HS65_LS_NAND2X7 U44 ( .A(phitOut2[15]), .B(n572), .Z(n518) );
  HS65_LS_OR2X9 U45 ( .A(n21), .B(n480), .Z(n42) );
  HS65_LS_CBI4I1X11 U46 ( .A(n459), .B(n49), .C(n690), .D(n462), .Z(n469) );
  HS65_LS_IVX4 U47 ( .A(state_cnt[1]), .Z(n19) );
  HS65_LS_NAND2X5 U48 ( .A(state_cnt[1]), .B(n448), .Z(n451) );
  HS65_LS_NAND2X5 U49 ( .A(state_cnt[0]), .B(state_cnt[1]), .Z(n462) );
  HS65_LS_NAND2X5 U50 ( .A(phitOut2[21]), .B(n25), .Z(n536) );
  HS65_LS_NAND2X5 U51 ( .A(phitOut2[7]), .B(n25), .Z(n494) );
  HS65_LS_NAND2X5 U52 ( .A(phitOut2[19]), .B(n25), .Z(n530) );
  HS65_LS_NAND2X5 U53 ( .A(phitOut2[5]), .B(n25), .Z(n488) );
  HS65_LS_NAND2X5 U54 ( .A(phitOut2[8]), .B(n25), .Z(n497) );
  HS65_LS_NAND2X5 U55 ( .A(phitOut2[25]), .B(n25), .Z(n548) );
  HS65_LS_NAND2X5 U56 ( .A(phitOut2[22]), .B(n25), .Z(n539) );
  HS65_LS_NAND2X5 U57 ( .A(phitOut2[33]), .B(n25), .Z(n573) );
  HS65_LS_NAND2X5 U58 ( .A(phitOut2[29]), .B(n25), .Z(n560) );
  HS65_LS_NAND2X7 U59 ( .A(phitOut2[14]), .B(n517), .Z(n514) );
  HS65_LH_IVX2 U60 ( .A(n466), .Z(n18) );
  HS65_LS_IVX18 U61 ( .A(n460), .Z(n481) );
  HS65_LS_IVX7 U62 ( .A(state_cnt[1]), .Z(n452) );
  HS65_LS_CBI4I1X11 U63 ( .A(n459), .B(n49), .C(n458), .D(n457), .Z(n460) );
  HS65_LS_BFX53 U64 ( .A(n32), .Z(n22) );
  HS65_LS_IVX18 U65 ( .A(n23), .Z(n24) );
  HS65_LS_IVX18 U66 ( .A(n454), .Z(n44) );
  HS65_LS_NAND2X21 U67 ( .A(n454), .B(n466), .Z(n461) );
  HS65_LS_IVX18 U68 ( .A(n24), .Z(n466) );
  HS65_LS_IVX18 U69 ( .A(n470), .Z(n129) );
  HS65_LS_NAND3X13 U70 ( .A(n506), .B(n51), .C(n50), .Z(pkt_out[11]) );
  HS65_LS_IVX9 U71 ( .A(n472), .Z(n578) );
  HS65_LS_IVX9 U72 ( .A(n448), .Z(n27) );
  HS65_LH_MUX21I1X3 U73 ( .D0(n18), .D1(\phase_next[1] ), .S0(n652), .Z(n686)
         );
  HS65_LS_NAND2X11 U74 ( .A(n44), .B(n24), .Z(n45) );
  HS65_LS_IVX27 U75 ( .A(n31), .Z(n28) );
  HS65_LS_NAND2X7 U76 ( .A(n461), .B(n45), .Z(n453) );
  HS65_LH_BFX4 U77 ( .A(n139), .Z(n34) );
  HS65_LS_BFX18 U78 ( .A(n120), .Z(n139) );
  HS65_LS_NAND2X14 U79 ( .A(n37), .B(n42), .Z(pkt_out[2]) );
  HS65_LS_IVX18 U80 ( .A(n35), .Z(n37) );
  HS65_LS_AND2X9 U81 ( .A(n26), .B(n468), .Z(n101) );
  HS65_LS_IVX9 U82 ( .A(n125), .Z(n39) );
  HS65_LS_IVX18 U83 ( .A(n39), .Z(n41) );
  HS65_LS_IVX27 U84 ( .A(n17), .Z(n572) );
  HS65_LS_NAND2X14 U85 ( .A(n461), .B(n45), .Z(n467) );
  HS65_LS_AND2X18 U86 ( .A(n19), .B(n453), .Z(n49) );
  HS65_LS_IVX18 U87 ( .A(\phase_prev[0] ), .Z(n454) );
  HS65_LS_BFX9 U88 ( .A(n335), .Z(n331) );
  HS65_LS_BFX9 U89 ( .A(n335), .Z(n330) );
  HS65_LS_BFX9 U90 ( .A(n324), .Z(n310) );
  HS65_LS_BFX9 U91 ( .A(n324), .Z(n311) );
  HS65_LS_AND2X18 U92 ( .A(n448), .B(n452), .Z(n120) );
  HS65_LS_BFX9 U93 ( .A(n298), .Z(n301) );
  HS65_LS_BFX9 U94 ( .A(n340), .Z(n358) );
  HS65_LS_BFX9 U95 ( .A(n339), .Z(n357) );
  HS65_LS_BFX9 U96 ( .A(n339), .Z(n356) );
  HS65_LH_NAND2X2 U97 ( .A(n27), .B(n19), .Z(n365) );
  HS65_LS_OR2X18 U98 ( .A(n21), .B(n507), .Z(n50) );
  HS65_LS_IVX9 U99 ( .A(n331), .Z(n325) );
  HS65_LS_IVX9 U100 ( .A(n331), .Z(n326) );
  HS65_LS_IVX9 U101 ( .A(n330), .Z(n327) );
  HS65_LS_IVX9 U102 ( .A(n330), .Z(n328) );
  HS65_LS_IVX9 U103 ( .A(n330), .Z(n329) );
  HS65_LS_AND2X4 U104 ( .A(n619), .B(n618), .Z(n52) );
  HS65_LS_AND2X4 U105 ( .A(n605), .B(n90), .Z(n53) );
  HS65_LS_AND2X4 U106 ( .A(n606), .B(n53), .Z(n54) );
  HS65_LS_AND2X4 U107 ( .A(n607), .B(n54), .Z(n55) );
  HS65_LS_AND2X4 U108 ( .A(n608), .B(n55), .Z(n56) );
  HS65_LS_AND2X4 U109 ( .A(n609), .B(n56), .Z(n57) );
  HS65_LS_AND2X4 U110 ( .A(n610), .B(n57), .Z(n58) );
  HS65_LS_AND2X4 U111 ( .A(n611), .B(n58), .Z(n59) );
  HS65_LS_AND2X4 U112 ( .A(n612), .B(n59), .Z(n62) );
  HS65_LS_AND2X4 U113 ( .A(n613), .B(n62), .Z(n64) );
  HS65_LS_AND2X4 U114 ( .A(n614), .B(n64), .Z(n72) );
  HS65_LS_AND2X4 U115 ( .A(n615), .B(n72), .Z(n73) );
  HS65_LS_AND2X4 U116 ( .A(n624), .B(n91), .Z(n74) );
  HS65_LS_AND2X4 U117 ( .A(n620), .B(n52), .Z(n75) );
  HS65_LS_AND2X4 U118 ( .A(n621), .B(n75), .Z(n77) );
  HS65_LS_AND2X4 U119 ( .A(n622), .B(n77), .Z(n78) );
  HS65_LS_AND2X4 U120 ( .A(\add_545/A[8] ), .B(n74), .Z(n79) );
  HS65_LS_AND2X4 U121 ( .A(\add_545/A[9] ), .B(n79), .Z(n80) );
  HS65_LS_AND2X4 U122 ( .A(\add_545/A[10] ), .B(n80), .Z(n84) );
  HS65_LS_AND2X4 U123 ( .A(\add_545/A[11] ), .B(n84), .Z(n87) );
  HS65_LS_AND2X4 U124 ( .A(\add_545/A[12] ), .B(n87), .Z(n88) );
  HS65_LS_AND2X4 U125 ( .A(\add_545/A[13] ), .B(n88), .Z(n89) );
  HS65_LS_AND2X4 U126 ( .A(n604), .B(n603), .Z(n90) );
  HS65_LS_AND2X4 U127 ( .A(n623), .B(n78), .Z(n91) );
  HS65_LS_BFX9 U128 ( .A(n334), .Z(n332) );
  HS65_LS_BFX9 U129 ( .A(n334), .Z(n333) );
  HS65_LS_IVX9 U130 ( .A(n310), .Z(n306) );
  HS65_LS_IVX9 U131 ( .A(n311), .Z(n305) );
  HS65_LS_IVX9 U132 ( .A(n311), .Z(n304) );
  HS65_LS_OAI21X3 U133 ( .A(n871), .B(n859), .C(n325), .Z(dma_wen[2]) );
  HS65_LS_NOR2AX3 U134 ( .A(n857), .B(n601), .Z(n871) );
  HS65_LS_IVX9 U135 ( .A(n855), .Z(n601) );
  HS65_LSS_XNOR2X6 U136 ( .A(n111), .B(\sub_544/A[10] ), .Z(dma_cnt_new[10])
         );
  HS65_LSS_XNOR2X6 U137 ( .A(n104), .B(\sub_544/A[5] ), .Z(dma_cnt_new[5]) );
  HS65_LSS_XNOR2X6 U138 ( .A(n109), .B(\sub_544/A[9] ), .Z(dma_cnt_new[9]) );
  HS65_LSS_XNOR2X6 U139 ( .A(n103), .B(\sub_544/A[4] ), .Z(dma_cnt_new[4]) );
  HS65_LSS_XNOR2X6 U140 ( .A(n108), .B(\sub_544/A[8] ), .Z(dma_cnt_new[8]) );
  HS65_LS_NOR4ABX2 U141 ( .A(n114), .B(n116), .C(n867), .D(dma_cnt_new[13]), 
        .Z(n849) );
  HS65_LSS_XOR2X6 U142 ( .A(n106), .B(\sub_544/A[7] ), .Z(n93) );
  HS65_LSS_XOR2X6 U143 ( .A(n102), .B(\sub_544/A[3] ), .Z(n94) );
  HS65_LSS_XOR2X6 U144 ( .A(n105), .B(\sub_544/A[6] ), .Z(n95) );
  HS65_LS_IVX9 U145 ( .A(n881), .Z(\add_545/A[8] ) );
  HS65_LS_IVX9 U146 ( .A(n882), .Z(\add_545/A[9] ) );
  HS65_LS_IVX9 U147 ( .A(n883), .Z(\add_545/A[10] ) );
  HS65_LS_IVX9 U148 ( .A(n876), .Z(\add_545/A[11] ) );
  HS65_LS_IVX9 U149 ( .A(n877), .Z(\add_545/A[12] ) );
  HS65_LS_IVX9 U150 ( .A(n878), .Z(\add_545/A[13] ) );
  HS65_LS_BFX9 U151 ( .A(n118), .Z(n334) );
  HS65_LS_BFX9 U152 ( .A(n118), .Z(n335) );
  HS65_LS_OR2X9 U153 ( .A(\sub_544/A[2] ), .B(\sub_544/A[1] ), .Z(n102) );
  HS65_LS_OR2X9 U154 ( .A(\sub_544/A[3] ), .B(n102), .Z(n103) );
  HS65_LS_OR2X9 U155 ( .A(\sub_544/A[4] ), .B(n103), .Z(n104) );
  HS65_LS_OR2X9 U156 ( .A(\sub_544/A[5] ), .B(n104), .Z(n105) );
  HS65_LS_OR2X9 U157 ( .A(\sub_544/A[6] ), .B(n105), .Z(n106) );
  HS65_LS_OR2X9 U158 ( .A(\sub_544/A[7] ), .B(n106), .Z(n108) );
  HS65_LS_OR2X9 U159 ( .A(\sub_544/A[8] ), .B(n108), .Z(n109) );
  HS65_LS_OR2X9 U160 ( .A(\sub_544/A[9] ), .B(n109), .Z(n111) );
  HS65_LS_OR2X9 U161 ( .A(\sub_544/A[10] ), .B(n111), .Z(n112) );
  HS65_LS_OR2X9 U162 ( .A(\sub_544/A[11] ), .B(n112), .Z(n113) );
  HS65_LSS_XOR2X6 U163 ( .A(n112), .B(\sub_544/A[11] ), .Z(n114) );
  HS65_LSS_XOR2X6 U164 ( .A(n113), .B(\sub_544/A[12] ), .Z(n116) );
  HS65_LS_BFX9 U165 ( .A(n625), .Z(n144) );
  HS65_LS_BFX9 U166 ( .A(n625), .Z(n149) );
  HS65_LS_BFX9 U167 ( .A(n625), .Z(n293) );
  HS65_LS_BFX9 U168 ( .A(n4), .Z(n130) );
  HS65_LS_BFX9 U169 ( .A(n4), .Z(n132) );
  HS65_LS_BFX9 U170 ( .A(n4), .Z(n133) );
  HS65_LS_IVX9 U171 ( .A(n879), .Z(\add_545/A[14] ) );
  HS65_LS_IVX9 U172 ( .A(n301), .Z(n299) );
  HS65_LS_IVX9 U173 ( .A(n301), .Z(n300) );
  HS65_LSS_XOR2X6 U174 ( .A(\sub_544/A[1] ), .B(\sub_544/A[2] ), .Z(n117) );
  HS65_LS_BFX9 U175 ( .A(n324), .Z(n312) );
  HS65_LS_BFX9 U176 ( .A(n324), .Z(n314) );
  HS65_LS_BFX9 U177 ( .A(n324), .Z(n313) );
  HS65_LS_BFX9 U178 ( .A(n294), .Z(n296) );
  HS65_LS_BFX9 U179 ( .A(n294), .Z(n295) );
  HS65_LS_BFX9 U180 ( .A(n324), .Z(n323) );
  HS65_LS_BFX9 U181 ( .A(n134), .Z(n136) );
  HS65_LS_BFX9 U182 ( .A(n134), .Z(n137) );
  HS65_LS_BFX9 U183 ( .A(n294), .Z(n297) );
  HS65_LS_BFX9 U184 ( .A(n134), .Z(n138) );
  HS65_LS_IVX9 U185 ( .A(n859), .Z(n657) );
  HS65_LS_IVX9 U186 ( .A(\proc_out[SRESP] ), .Z(n336) );
  HS65_LS_IVX9 U187 ( .A(n358), .Z(n349) );
  HS65_LS_IVX9 U188 ( .A(n358), .Z(n348) );
  HS65_LS_IVX9 U189 ( .A(n358), .Z(n352) );
  HS65_LS_IVX9 U190 ( .A(n358), .Z(n350) );
  HS65_LS_IVX9 U191 ( .A(n358), .Z(n351) );
  HS65_LS_IVX9 U192 ( .A(n357), .Z(n347) );
  HS65_LS_IVX9 U193 ( .A(n357), .Z(n346) );
  HS65_LS_IVX9 U194 ( .A(n357), .Z(n344) );
  HS65_LS_IVX9 U195 ( .A(n357), .Z(n343) );
  HS65_LS_IVX9 U196 ( .A(n357), .Z(n342) );
  HS65_LS_IVX9 U197 ( .A(n357), .Z(n345) );
  HS65_LS_IVX9 U198 ( .A(n359), .Z(n355) );
  HS65_LS_IVX9 U199 ( .A(n359), .Z(n354) );
  HS65_LS_IVX9 U200 ( .A(n359), .Z(n353) );
  HS65_LS_IVX9 U201 ( .A(n356), .Z(n341) );
  HS65_LS_NOR2X6 U202 ( .A(n359), .B(n881), .Z(\spm_out[MADDR][7] ) );
  HS65_LS_NOR2X6 U203 ( .A(n359), .B(n882), .Z(\spm_out[MADDR][8] ) );
  HS65_LS_NOR2X6 U204 ( .A(n359), .B(n883), .Z(\spm_out[MADDR][9] ) );
  HS65_LS_NOR2X6 U205 ( .A(n359), .B(n876), .Z(\spm_out[MADDR][10] ) );
  HS65_LS_NOR2X6 U206 ( .A(n359), .B(n877), .Z(\spm_out[MADDR][11] ) );
  HS65_LS_NOR2X6 U207 ( .A(n359), .B(n878), .Z(\spm_out[MADDR][12] ) );
  HS65_LS_NOR2X6 U208 ( .A(n359), .B(n879), .Z(\spm_out[MADDR][13] ) );
  HS65_LS_NOR2X6 U209 ( .A(n359), .B(n880), .Z(\spm_out[MADDR][14] ) );
  HS65_LS_NOR2X6 U210 ( .A(n336), .B(n647), .Z(\proc_out[SDATA][0] ) );
  HS65_LS_NOR2X6 U211 ( .A(n336), .B(n646), .Z(\proc_out[SDATA][1] ) );
  HS65_LS_NOR2X6 U212 ( .A(n336), .B(n645), .Z(\proc_out[SDATA][2] ) );
  HS65_LS_NOR2X6 U213 ( .A(n875), .B(n644), .Z(\proc_out[SDATA][3] ) );
  HS65_LS_NOR2X6 U214 ( .A(n336), .B(n643), .Z(\proc_out[SDATA][4] ) );
  HS65_LS_NOR2X6 U215 ( .A(n875), .B(n642), .Z(\proc_out[SDATA][5] ) );
  HS65_LS_NOR2X6 U216 ( .A(n875), .B(n641), .Z(\proc_out[SDATA][6] ) );
  HS65_LS_NOR2X6 U217 ( .A(n875), .B(n640), .Z(\proc_out[SDATA][7] ) );
  HS65_LS_NOR2X6 U218 ( .A(n336), .B(n639), .Z(\proc_out[SDATA][8] ) );
  HS65_LS_NOR2X6 U219 ( .A(n336), .B(n638), .Z(\proc_out[SDATA][9] ) );
  HS65_LS_NOR2X6 U220 ( .A(n336), .B(n637), .Z(\proc_out[SDATA][10] ) );
  HS65_LS_NOR2X6 U221 ( .A(n336), .B(n636), .Z(\proc_out[SDATA][11] ) );
  HS65_LS_NOR2X6 U222 ( .A(n336), .B(n635), .Z(\proc_out[SDATA][12] ) );
  HS65_LS_NOR2X6 U223 ( .A(n336), .B(n634), .Z(\proc_out[SDATA][13] ) );
  HS65_LS_NOR2X6 U224 ( .A(n336), .B(n633), .Z(\proc_out[SDATA][14] ) );
  HS65_LS_NOR2X6 U225 ( .A(n336), .B(n632), .Z(\proc_out[SDATA][15] ) );
  HS65_LS_OAI222X2 U226 ( .A(n331), .B(n841), .C(n854), .D(n679), .E(n325), 
        .F(n841), .Z(dma_wdata[48]) );
  HS65_LS_NOR2X6 U227 ( .A(n871), .B(n858), .Z(dma_wen[0]) );
  HS65_LS_OAI222X2 U228 ( .A(n331), .B(n842), .C(n854), .D(n676), .E(n325), 
        .F(n94), .Z(dma_wdata[51]) );
  HS65_LS_OAI222X2 U229 ( .A(n331), .B(n843), .C(n854), .D(n675), .E(n325), 
        .F(n631), .Z(dma_wdata[52]) );
  HS65_LS_IVX9 U230 ( .A(dma_cnt_new[4]), .Z(n631) );
  HS65_LS_OAI222X2 U231 ( .A(n331), .B(n844), .C(n672), .D(n854), .E(n325), 
        .F(n93), .Z(dma_wdata[55]) );
  HS65_LS_OAI222X2 U232 ( .A(n331), .B(n845), .C(n671), .D(n854), .E(n325), 
        .F(n629), .Z(dma_wdata[56]) );
  HS65_LS_IVX9 U233 ( .A(dma_cnt_new[8]), .Z(n629) );
  HS65_LS_OAI222X2 U234 ( .A(n331), .B(n846), .C(n854), .D(n669), .E(n326), 
        .F(n627), .Z(dma_wdata[58]) );
  HS65_LS_IVX9 U235 ( .A(dma_cnt_new[10]), .Z(n627) );
  HS65_LS_OAI222X2 U236 ( .A(n330), .B(n847), .C(n854), .D(n667), .E(n326), 
        .F(n116), .Z(dma_wdata[60]) );
  HS65_LS_OAI222X2 U237 ( .A(n331), .B(n848), .C(n854), .D(n666), .E(n325), 
        .F(n626), .Z(dma_wdata[61]) );
  HS65_LS_IVX9 U238 ( .A(dma_cnt_new[13]), .Z(n626) );
  HS65_LS_OAI222X2 U239 ( .A(n331), .B(n867), .C(n854), .D(n678), .E(n325), 
        .F(\sub_544/A[1] ), .Z(dma_wdata[49]) );
  HS65_LS_OAI222X2 U240 ( .A(n331), .B(n866), .C(n854), .D(n677), .E(n325), 
        .F(n117), .Z(dma_wdata[50]) );
  HS65_LS_OAI222X2 U241 ( .A(n331), .B(n865), .C(n854), .D(n674), .E(n325), 
        .F(n630), .Z(dma_wdata[53]) );
  HS65_LS_IVX9 U242 ( .A(dma_cnt_new[5]), .Z(n630) );
  HS65_LS_OAI222X2 U243 ( .A(n331), .B(n864), .C(n673), .D(n854), .E(n325), 
        .F(n95), .Z(dma_wdata[54]) );
  HS65_LS_OAI222X2 U244 ( .A(n331), .B(n863), .C(n670), .D(n854), .E(n325), 
        .F(n628), .Z(dma_wdata[57]) );
  HS65_LS_IVX9 U245 ( .A(dma_cnt_new[9]), .Z(n628) );
  HS65_LS_OAI222X2 U246 ( .A(n331), .B(n862), .C(n854), .D(n668), .E(n325), 
        .F(n114), .Z(dma_wdata[59]) );
  HS65_LS_OAI212X5 U247 ( .A(n854), .B(n665), .C(n856), .D(n649), .E(n853), 
        .Z(dma_wdata[62]) );
  HS65_LS_NAND4ABX3 U248 ( .A(n852), .B(n851), .C(n850), .D(n849), .Z(n853) );
  HS65_LS_NAND4ABX3 U249 ( .A(dma_cnt_new[5]), .B(dma_cnt_new[4]), .C(n117), 
        .D(n94), .Z(n851) );
  HS65_LS_NAND4ABX3 U250 ( .A(dma_cnt_new[9]), .B(dma_cnt_new[8]), .C(n95), 
        .D(n93), .Z(n852) );
  HS65_LS_NAND2X7 U251 ( .A(n656), .B(n1), .Z(n855) );
  HS65_LS_AND3X9 U252 ( .A(dma_rdata[63]), .B(n649), .C(n293), .Z(n118) );
  HS65_LS_OAI21X3 U253 ( .A(n871), .B(n861), .C(n325), .Z(dma_wen[1]) );
  HS65_LS_NAND2X7 U254 ( .A(n365), .B(n128), .Z(n597) );
  HS65_LS_NOR3X4 U255 ( .A(n325), .B(dma_cnt_new[10]), .C(dma_cnt_new[0]), .Z(
        n850) );
  HS65_LS_IVX9 U256 ( .A(n841), .Z(dma_cnt_new[0]) );
  HS65_LS_IVX9 U257 ( .A(n867), .Z(\sub_544/A[1] ) );
  HS65_LS_NAND2X7 U258 ( .A(dma_rdata[40]), .B(n144), .Z(n881) );
  HS65_LS_NAND2X7 U259 ( .A(dma_rdata[41]), .B(n144), .Z(n882) );
  HS65_LS_NAND2X7 U260 ( .A(dma_rdata[42]), .B(n144), .Z(n883) );
  HS65_LS_NAND2X7 U261 ( .A(dma_rdata[43]), .B(n144), .Z(n876) );
  HS65_LS_NAND2X7 U262 ( .A(dma_rdata[44]), .B(n144), .Z(n877) );
  HS65_LS_NAND2X7 U263 ( .A(dma_rdata[45]), .B(n149), .Z(n878) );
  HS65_LS_IVX9 U264 ( .A(n842), .Z(\sub_544/A[3] ) );
  HS65_LS_IVX9 U265 ( .A(n843), .Z(\sub_544/A[4] ) );
  HS65_LS_IVX9 U266 ( .A(n844), .Z(\sub_544/A[7] ) );
  HS65_LS_IVX9 U267 ( .A(n845), .Z(\sub_544/A[8] ) );
  HS65_LS_IVX9 U268 ( .A(n846), .Z(\sub_544/A[10] ) );
  HS65_LS_IVX9 U269 ( .A(n866), .Z(\sub_544/A[2] ) );
  HS65_LS_IVX9 U270 ( .A(n865), .Z(\sub_544/A[5] ) );
  HS65_LS_IVX9 U271 ( .A(n864), .Z(\sub_544/A[6] ) );
  HS65_LS_IVX9 U272 ( .A(n863), .Z(\sub_544/A[9] ) );
  HS65_LS_IVX9 U273 ( .A(n862), .Z(\sub_544/A[11] ) );
  HS65_LSS_XNOR2X6 U274 ( .A(n848), .B(n127), .Z(dma_cnt_new[13]) );
  HS65_LS_NOR2X6 U275 ( .A(\sub_544/A[12] ), .B(n113), .Z(n127) );
  HS65_LS_OAI22X6 U276 ( .A(n856), .B(n648), .C(n854), .D(n664), .Z(
        dma_wdata[63]) );
  HS65_LS_IVX9 U277 ( .A(dma_rdata[63]), .Z(n648) );
  HS65_LS_OAI22X6 U278 ( .A(n856), .B(n647), .C(n855), .D(n679), .Z(
        dma_wdata[0]) );
  HS65_LS_OAI22X6 U279 ( .A(n856), .B(n646), .C(n855), .D(n678), .Z(
        dma_wdata[1]) );
  HS65_LS_OAI22X6 U280 ( .A(n856), .B(n645), .C(n855), .D(n677), .Z(
        dma_wdata[2]) );
  HS65_LS_OAI22X6 U281 ( .A(n856), .B(n644), .C(n855), .D(n676), .Z(
        dma_wdata[3]) );
  HS65_LS_OAI22X6 U282 ( .A(n856), .B(n643), .C(n855), .D(n675), .Z(
        dma_wdata[4]) );
  HS65_LS_OAI22X6 U283 ( .A(n856), .B(n642), .C(n855), .D(n674), .Z(
        dma_wdata[5]) );
  HS65_LS_OAI22X6 U284 ( .A(n856), .B(n641), .C(n855), .D(n673), .Z(
        dma_wdata[6]) );
  HS65_LS_OAI22X6 U285 ( .A(n856), .B(n640), .C(n855), .D(n672), .Z(
        dma_wdata[7]) );
  HS65_LS_OAI22X6 U286 ( .A(n856), .B(n639), .C(n855), .D(n671), .Z(
        dma_wdata[8]) );
  HS65_LS_OAI22X6 U287 ( .A(n856), .B(n638), .C(n855), .D(n670), .Z(
        dma_wdata[9]) );
  HS65_LS_OAI22X6 U288 ( .A(n856), .B(n637), .C(n855), .D(n669), .Z(
        dma_wdata[10]) );
  HS65_LS_OAI22X6 U289 ( .A(n856), .B(n636), .C(n855), .D(n668), .Z(
        dma_wdata[11]) );
  HS65_LS_OAI22X6 U290 ( .A(n856), .B(n635), .C(n855), .D(n667), .Z(
        dma_wdata[12]) );
  HS65_LS_OAI22X6 U291 ( .A(n856), .B(n634), .C(n855), .D(n666), .Z(
        dma_wdata[13]) );
  HS65_LS_OAI22X6 U292 ( .A(n856), .B(n633), .C(n855), .D(n665), .Z(
        dma_wdata[14]) );
  HS65_LS_OAI22X6 U293 ( .A(n856), .B(n632), .C(n855), .D(n664), .Z(
        dma_wdata[15]) );
  HS65_LS_OAI21X3 U294 ( .A(n656), .B(n839), .C(n361), .Z(n598) );
  HS65_LS_NAND2X7 U295 ( .A(n657), .B(n1), .Z(n854) );
  HS65_LS_IVX9 U296 ( .A(n868), .Z(n653) );
  HS65_LS_OAI21X3 U297 ( .A(n858), .B(n598), .C(n365), .Z(dma_ren[0]) );
  HS65_LH_OAI21X2 U298 ( .A(n861), .B(n598), .C(n365), .Z(dma_ren[1]) );
  HS65_LH_OAI21X2 U299 ( .A(n859), .B(n598), .C(n365), .Z(dma_ren[2]) );
  HS65_LS_NAND2X7 U300 ( .A(dma_rdata[46]), .B(n149), .Z(n879) );
  HS65_LS_NAND2X7 U301 ( .A(dma_rdata[47]), .B(n149), .Z(n880) );
  HS65_LS_IVX9 U302 ( .A(dma_rdata[0]), .Z(n647) );
  HS65_LS_IVX9 U303 ( .A(dma_rdata[1]), .Z(n646) );
  HS65_LS_IVX9 U304 ( .A(dma_rdata[2]), .Z(n645) );
  HS65_LS_IVX9 U305 ( .A(dma_rdata[3]), .Z(n644) );
  HS65_LS_IVX9 U306 ( .A(dma_rdata[4]), .Z(n643) );
  HS65_LS_IVX9 U307 ( .A(dma_rdata[5]), .Z(n642) );
  HS65_LS_IVX9 U308 ( .A(dma_rdata[6]), .Z(n641) );
  HS65_LS_IVX9 U309 ( .A(dma_rdata[7]), .Z(n640) );
  HS65_LS_IVX9 U310 ( .A(dma_rdata[8]), .Z(n639) );
  HS65_LS_IVX9 U311 ( .A(dma_rdata[9]), .Z(n638) );
  HS65_LS_IVX9 U312 ( .A(dma_rdata[10]), .Z(n637) );
  HS65_LS_IVX9 U313 ( .A(dma_rdata[11]), .Z(n636) );
  HS65_LS_IVX9 U314 ( .A(dma_rdata[12]), .Z(n635) );
  HS65_LS_IVX9 U315 ( .A(dma_rdata[13]), .Z(n634) );
  HS65_LS_IVX9 U316 ( .A(dma_rdata[14]), .Z(n633) );
  HS65_LS_IVX9 U317 ( .A(dma_rdata[15]), .Z(n632) );
  HS65_LS_IVX9 U318 ( .A(n847), .Z(\sub_544/A[12] ) );
  HS65_LS_BFX9 U319 ( .A(n414), .Z(n134) );
  HS65_LS_BFX9 U320 ( .A(n840), .Z(n294) );
  HS65_LS_NOR2AX3 U321 ( .A(n1), .B(n861), .Z(n840) );
  HS65_LS_BFX9 U322 ( .A(n298), .Z(n302) );
  HS65_LS_IVX9 U323 ( .A(n870), .Z(n324) );
  HS65_LS_BFX9 U324 ( .A(n298), .Z(n303) );
  HS65_LS_NAND3X2 U325 ( .A(n140), .B(n581), .C(n341), .Z(n596) );
  HS65_LS_IVX9 U326 ( .A(n858), .Z(n656) );
  HS65_LS_NAND2X7 U327 ( .A(n859), .B(n861), .Z(n839) );
  HS65_LS_NAND2X7 U328 ( .A(n836), .B(n663), .Z(n859) );
  HS65_LS_BFX9 U329 ( .A(n338), .Z(\proc_out[SRESP] ) );
  HS65_LS_IVX9 U330 ( .A(n875), .Z(n338) );
  HS65_LS_BFX9 U331 ( .A(n340), .Z(n359) );
  HS65_LS_IVX9 U332 ( .A(n872), .Z(n655) );
  HS65_LS_NOR2AX3 U333 ( .A(dma_rdata[16]), .B(n875), .Z(\proc_out[SDATA][16] ) );
  HS65_LS_NOR2AX3 U334 ( .A(dma_rdata[17]), .B(n875), .Z(\proc_out[SDATA][17] ) );
  HS65_LS_NOR2AX3 U335 ( .A(dma_rdata[18]), .B(n875), .Z(\proc_out[SDATA][18] ) );
  HS65_LS_NOR2AX3 U336 ( .A(dma_rdata[19]), .B(n875), .Z(\proc_out[SDATA][19] ) );
  HS65_LS_NOR2AX3 U337 ( .A(dma_rdata[20]), .B(n875), .Z(\proc_out[SDATA][20] ) );
  HS65_LS_NOR2AX3 U338 ( .A(dma_rdata[21]), .B(n875), .Z(\proc_out[SDATA][21] ) );
  HS65_LS_NOR2AX3 U339 ( .A(dma_rdata[22]), .B(n875), .Z(\proc_out[SDATA][22] ) );
  HS65_LS_NOR2AX3 U340 ( .A(dma_rdata[23]), .B(n875), .Z(\proc_out[SDATA][23] ) );
  HS65_LS_NOR2AX3 U341 ( .A(dma_rdata[24]), .B(n875), .Z(\proc_out[SDATA][24] ) );
  HS65_LS_NOR2AX3 U342 ( .A(dma_rdata[25]), .B(n875), .Z(\proc_out[SDATA][25] ) );
  HS65_LS_NOR2AX3 U343 ( .A(dma_rdata[26]), .B(n336), .Z(\proc_out[SDATA][26] ) );
  HS65_LS_NOR2AX3 U344 ( .A(dma_rdata[27]), .B(n875), .Z(\proc_out[SDATA][27] ) );
  HS65_LS_NOR2AX3 U345 ( .A(dma_rdata[28]), .B(n875), .Z(\proc_out[SDATA][28] ) );
  HS65_LS_NOR2AX3 U346 ( .A(dma_rdata[29]), .B(n336), .Z(\proc_out[SDATA][29] ) );
  HS65_LS_NOR2AX3 U347 ( .A(dma_rdata[30]), .B(n875), .Z(\proc_out[SDATA][30] ) );
  HS65_LS_NOR2AX3 U348 ( .A(dma_rdata[31]), .B(n875), .Z(\proc_out[SDATA][31] ) );
  HS65_LS_IVX9 U349 ( .A(n861), .Z(n658) );
  HS65_LS_AOI22X6 U350 ( .A(\proc_in[MADDR][1] ), .B(n656), .C(
        \proc_in[MADDR][2] ), .D(n839), .Z(n838) );
  HS65_LS_IVX9 U351 ( .A(\proc_in[MADDR][2] ), .Z(n661) );
  HS65_LS_NAND2X7 U352 ( .A(slt_entry[4]), .B(n652), .Z(n856) );
  HS65_LS_NAND3X5 U353 ( .A(n128), .B(n581), .C(n306), .Z(n363) );
  HS65_LS_OAI21X3 U354 ( .A(n652), .B(n140), .C(n360), .Z(n362) );
  HS65_LH_MUXI21X2 U355 ( .D0(n690), .D1(n122), .S0(n652), .Z(n682) );
  HS65_LS_NOR2X6 U356 ( .A(slt_entry[0]), .B(n327), .Z(n122) );
  HS65_LS_MUXI21X2 U357 ( .D0(n458), .D1(n124), .S0(n652), .Z(n681) );
  HS65_LS_NOR2X6 U358 ( .A(slt_entry[1]), .B(n327), .Z(n124) );
  HS65_LS_OAI21X3 U359 ( .A(n689), .B(n652), .C(n327), .Z(n683) );
  HS65_LS_MX41X7 U360 ( .D0(n600), .S0(n332), .D1(n600), .S1(n326), .D2(
        \proc_in[MDATA][16] ), .S2(n601), .D3(n295), .S3(\proc_in[MDATA][0] ), 
        .Z(dma_wdata[16]) );
  HS65_LS_MX41X7 U361 ( .D0(n385), .S0(n331), .D1(n603), .S1(n326), .D2(
        \proc_in[MDATA][17] ), .S2(n601), .D3(n295), .S3(\proc_in[MDATA][1] ), 
        .Z(dma_wdata[17]) );
  HS65_LS_MX41X7 U362 ( .D0(dma_wp_new[2]), .S0(n331), .D1(n604), .S1(n326), 
        .D2(\proc_in[MDATA][18] ), .S2(n601), .D3(n295), .S3(
        \proc_in[MDATA][2] ), .Z(dma_wdata[18]) );
  HS65_LSS_XOR2X6 U363 ( .A(n603), .B(n604), .Z(dma_wp_new[2]) );
  HS65_LS_MX41X7 U364 ( .D0(dma_wp_new[3]), .S0(n331), .D1(n605), .S1(n326), 
        .D2(\proc_in[MDATA][19] ), .S2(n601), .D3(n295), .S3(
        \proc_in[MDATA][3] ), .Z(dma_wdata[19]) );
  HS65_LSS_XOR2X6 U365 ( .A(n90), .B(n605), .Z(dma_wp_new[3]) );
  HS65_LS_MX41X7 U366 ( .D0(dma_wp_new[4]), .S0(n331), .D1(n606), .S1(n326), 
        .D2(\proc_in[MDATA][20] ), .S2(n601), .D3(n295), .S3(
        \proc_in[MDATA][4] ), .Z(dma_wdata[20]) );
  HS65_LSS_XOR2X6 U367 ( .A(n53), .B(n606), .Z(dma_wp_new[4]) );
  HS65_LS_MX41X7 U368 ( .D0(dma_wp_new[5]), .S0(n331), .D1(n607), .S1(n326), 
        .D2(\proc_in[MDATA][21] ), .S2(n601), .D3(n295), .S3(
        \proc_in[MDATA][5] ), .Z(dma_wdata[21]) );
  HS65_LSS_XOR2X6 U369 ( .A(n54), .B(n607), .Z(dma_wp_new[5]) );
  HS65_LS_MX41X7 U370 ( .D0(dma_wp_new[6]), .S0(n332), .D1(n608), .S1(n326), 
        .D2(\proc_in[MDATA][22] ), .S2(n601), .D3(n295), .S3(
        \proc_in[MDATA][6] ), .Z(dma_wdata[22]) );
  HS65_LSS_XOR2X6 U371 ( .A(n55), .B(n608), .Z(dma_wp_new[6]) );
  HS65_LS_MX41X7 U372 ( .D0(dma_wp_new[7]), .S0(n332), .D1(n609), .S1(n326), 
        .D2(\proc_in[MDATA][23] ), .S2(n601), .D3(n295), .S3(
        \proc_in[MDATA][7] ), .Z(dma_wdata[23]) );
  HS65_LSS_XOR2X6 U373 ( .A(n56), .B(n609), .Z(dma_wp_new[7]) );
  HS65_LS_MX41X7 U374 ( .D0(dma_wp_new[8]), .S0(n332), .D1(n610), .S1(n326), 
        .D2(\proc_in[MDATA][24] ), .S2(n601), .D3(n295), .S3(
        \proc_in[MDATA][8] ), .Z(dma_wdata[24]) );
  HS65_LSS_XOR2X6 U375 ( .A(n57), .B(n610), .Z(dma_wp_new[8]) );
  HS65_LS_MX41X7 U376 ( .D0(dma_wp_new[9]), .S0(n332), .D1(n611), .S1(n326), 
        .D2(\proc_in[MDATA][25] ), .S2(n601), .D3(n295), .S3(
        \proc_in[MDATA][9] ), .Z(dma_wdata[25]) );
  HS65_LSS_XOR2X6 U377 ( .A(n58), .B(n611), .Z(dma_wp_new[9]) );
  HS65_LS_MX41X7 U378 ( .D0(dma_wp_new[10]), .S0(n332), .D1(n612), .S1(n326), 
        .D2(\proc_in[MDATA][26] ), .S2(n601), .D3(n295), .S3(
        \proc_in[MDATA][10] ), .Z(dma_wdata[26]) );
  HS65_LSS_XOR2X6 U379 ( .A(n59), .B(n612), .Z(dma_wp_new[10]) );
  HS65_LS_MX41X7 U380 ( .D0(dma_wp_new[11]), .S0(n332), .D1(n613), .S1(n326), 
        .D2(\proc_in[MDATA][27] ), .S2(n601), .D3(n295), .S3(
        \proc_in[MDATA][11] ), .Z(dma_wdata[27]) );
  HS65_LSS_XOR2X6 U381 ( .A(n62), .B(n613), .Z(dma_wp_new[11]) );
  HS65_LS_MX41X7 U382 ( .D0(dma_wp_new[12]), .S0(n332), .D1(n614), .S1(n326), 
        .D2(\proc_in[MDATA][28] ), .S2(n601), .D3(n296), .S3(
        \proc_in[MDATA][12] ), .Z(dma_wdata[28]) );
  HS65_LSS_XOR2X6 U383 ( .A(n64), .B(n614), .Z(dma_wp_new[12]) );
  HS65_LS_MX41X7 U384 ( .D0(dma_wp_new[13]), .S0(n332), .D1(n615), .S1(n326), 
        .D2(\proc_in[MDATA][29] ), .S2(n601), .D3(n296), .S3(
        \proc_in[MDATA][13] ), .Z(dma_wdata[29]) );
  HS65_LSS_XOR2X6 U385 ( .A(n72), .B(n615), .Z(dma_wp_new[13]) );
  HS65_LS_MX41X7 U386 ( .D0(dma_wp_new[14]), .S0(n332), .D1(n616), .S1(n326), 
        .D2(\proc_in[MDATA][30] ), .S2(n601), .D3(n296), .S3(
        \proc_in[MDATA][14] ), .Z(dma_wdata[30]) );
  HS65_LSS_XOR2X6 U387 ( .A(n73), .B(n616), .Z(dma_wp_new[14]) );
  HS65_LS_MX41X7 U388 ( .D0(dma_wp_new[15]), .S0(n332), .D1(n617), .S1(n326), 
        .D2(\proc_in[MDATA][31] ), .S2(n601), .D3(n296), .S3(
        \proc_in[MDATA][15] ), .Z(dma_wdata[31]) );
  HS65_LSS_XOR2X6 U389 ( .A(n617), .B(n2), .Z(dma_wp_new[15]) );
  HS65_LS_AO222X4 U390 ( .A(n618), .B(n327), .C(\proc_in[MDATA][17] ), .D(n296), .E(n583), .F(n332), .Z(dma_wdata[33]) );
  HS65_LS_AO222X4 U391 ( .A(n619), .B(n327), .C(\proc_in[MDATA][18] ), .D(n296), .E(dma_rp_new[2]), .F(n332), .Z(dma_wdata[34]) );
  HS65_LSS_XOR2X6 U392 ( .A(n618), .B(n619), .Z(dma_rp_new[2]) );
  HS65_LS_AO222X4 U393 ( .A(n620), .B(n327), .C(\proc_in[MDATA][19] ), .D(n296), .E(dma_rp_new[3]), .F(n332), .Z(dma_wdata[35]) );
  HS65_LSS_XOR2X6 U394 ( .A(n52), .B(n620), .Z(dma_rp_new[3]) );
  HS65_LS_AO222X4 U395 ( .A(n621), .B(n326), .C(\proc_in[MDATA][20] ), .D(n296), .E(dma_rp_new[4]), .F(n332), .Z(dma_wdata[36]) );
  HS65_LSS_XOR2X6 U396 ( .A(n75), .B(n621), .Z(dma_rp_new[4]) );
  HS65_LS_AO222X4 U397 ( .A(n622), .B(n327), .C(\proc_in[MDATA][21] ), .D(n296), .E(dma_rp_new[5]), .F(n332), .Z(dma_wdata[37]) );
  HS65_LSS_XOR2X6 U398 ( .A(n77), .B(n622), .Z(dma_rp_new[5]) );
  HS65_LS_AO222X4 U399 ( .A(n623), .B(n327), .C(\proc_in[MDATA][22] ), .D(n296), .E(dma_rp_new[6]), .F(n332), .Z(dma_wdata[38]) );
  HS65_LSS_XOR2X6 U400 ( .A(n78), .B(n623), .Z(dma_rp_new[6]) );
  HS65_LS_AO222X4 U401 ( .A(n624), .B(n327), .C(\proc_in[MDATA][23] ), .D(n296), .E(dma_rp_new[7]), .F(n332), .Z(dma_wdata[39]) );
  HS65_LSS_XOR2X6 U402 ( .A(n91), .B(n624), .Z(dma_rp_new[7]) );
  HS65_LS_AO222X4 U403 ( .A(\add_545/A[8] ), .B(n327), .C(\proc_in[MDATA][24] ), .D(n296), .E(dma_rp_new[8]), .F(n332), .Z(dma_wdata[40]) );
  HS65_LSS_XOR2X6 U404 ( .A(n74), .B(\add_545/A[8] ), .Z(dma_rp_new[8]) );
  HS65_LS_AO222X4 U405 ( .A(\add_545/A[9] ), .B(n327), .C(\proc_in[MDATA][25] ), .D(n297), .E(dma_rp_new[9]), .F(n333), .Z(dma_wdata[41]) );
  HS65_LSS_XOR2X6 U406 ( .A(n79), .B(\add_545/A[9] ), .Z(dma_rp_new[9]) );
  HS65_LS_AO222X4 U407 ( .A(\add_545/A[10] ), .B(n327), .C(
        \proc_in[MDATA][26] ), .D(n297), .E(dma_rp_new[10]), .F(n333), .Z(
        dma_wdata[42]) );
  HS65_LSS_XOR2X6 U408 ( .A(n80), .B(\add_545/A[10] ), .Z(dma_rp_new[10]) );
  HS65_LS_AO222X4 U409 ( .A(\add_545/A[11] ), .B(n327), .C(
        \proc_in[MDATA][27] ), .D(n297), .E(dma_rp_new[11]), .F(n333), .Z(
        dma_wdata[43]) );
  HS65_LSS_XOR2X6 U410 ( .A(n84), .B(\add_545/A[11] ), .Z(dma_rp_new[11]) );
  HS65_LS_AO222X4 U411 ( .A(\add_545/A[12] ), .B(n327), .C(
        \proc_in[MDATA][28] ), .D(n297), .E(dma_rp_new[12]), .F(n333), .Z(
        dma_wdata[44]) );
  HS65_LSS_XOR2X6 U412 ( .A(n87), .B(\add_545/A[12] ), .Z(dma_rp_new[12]) );
  HS65_LS_AO222X4 U413 ( .A(\add_545/A[13] ), .B(n327), .C(
        \proc_in[MDATA][29] ), .D(n297), .E(dma_rp_new[13]), .F(n333), .Z(
        dma_wdata[45]) );
  HS65_LSS_XOR2X6 U414 ( .A(n88), .B(\add_545/A[13] ), .Z(dma_rp_new[13]) );
  HS65_LS_AO222X4 U415 ( .A(\add_545/A[14] ), .B(n326), .C(
        \proc_in[MDATA][30] ), .D(n297), .E(dma_rp_new[14]), .F(n333), .Z(
        dma_wdata[46]) );
  HS65_LSS_XOR2X6 U416 ( .A(n89), .B(\add_545/A[14] ), .Z(dma_rp_new[14]) );
  HS65_LS_AO222X4 U417 ( .A(dma_rp_new[0]), .B(n327), .C(\proc_in[MDATA][16] ), 
        .D(n296), .E(dma_rp_new[0]), .F(n332), .Z(dma_wdata[32]) );
  HS65_LS_NOR2AX3 U418 ( .A(dma_rdata[32]), .B(n856), .Z(dma_rp_new[0]) );
  HS65_LS_AO222X4 U419 ( .A(\add_545/A[15] ), .B(n327), .C(
        \proc_in[MDATA][31] ), .D(n297), .E(dma_rp_new[15]), .F(n333), .Z(
        dma_wdata[47]) );
  HS65_LSS_XOR2X6 U420 ( .A(\add_545/A[15] ), .B(n3), .Z(dma_rp_new[15]) );
  HS65_LS_IVX9 U421 ( .A(n880), .Z(\add_545/A[15] ) );
  HS65_LS_AOI312X4 U422 ( .A(n465), .B(n466), .C(n467), .D(n464), .E(n27), .F(
        n463), .Z(n125) );
  HS65_LS_NAND2X7 U423 ( .A(dma_rdata[51]), .B(n144), .Z(n842) );
  HS65_LS_NAND2X7 U424 ( .A(dma_rdata[52]), .B(n144), .Z(n843) );
  HS65_LS_NAND2X7 U425 ( .A(dma_rdata[55]), .B(n144), .Z(n844) );
  HS65_LS_NAND2X7 U426 ( .A(dma_rdata[56]), .B(n144), .Z(n845) );
  HS65_LS_NAND2X7 U427 ( .A(dma_rdata[58]), .B(n144), .Z(n846) );
  HS65_LS_NAND2X7 U428 ( .A(dma_rdata[49]), .B(n149), .Z(n867) );
  HS65_LS_NAND2X7 U429 ( .A(dma_rdata[50]), .B(n149), .Z(n866) );
  HS65_LS_NAND2X7 U430 ( .A(dma_rdata[53]), .B(n149), .Z(n865) );
  HS65_LS_NAND2X7 U431 ( .A(dma_rdata[54]), .B(n149), .Z(n864) );
  HS65_LS_NAND2X7 U432 ( .A(dma_rdata[57]), .B(n149), .Z(n863) );
  HS65_LS_NAND2X7 U433 ( .A(dma_rdata[59]), .B(n149), .Z(n862) );
  HS65_LH_OAI12X2 U434 ( .A(state_cnt[1]), .B(n689), .C(n325), .Z(
        phit_togo[34]) );
  HS65_LS_IVX9 U435 ( .A(dma_rdata[62]), .Z(n649) );
  HS65_LS_IVX18 U436 ( .A(state_cnt[0]), .Z(n448) );
  HS65_LS_AOI22X6 U437 ( .A(\proc_in[MADDR][0] ), .B(n656), .C(
        \proc_in[MADDR][1] ), .D(n839), .Z(n837) );
  HS65_LS_NAND3AX6 U438 ( .A(phitIn[33]), .B(phitIn[32]), .C(phitIn[34]), .Z(
        n870) );
  HS65_LS_NAND2X7 U439 ( .A(phitIn[33]), .B(phitIn[34]), .Z(n868) );
  HS65_LS_NAND2X7 U440 ( .A(dma_rdata[48]), .B(n144), .Z(n841) );
  HS65_LS_NAND2X7 U441 ( .A(dma_rdata[60]), .B(n144), .Z(n847) );
  HS65_LS_NAND2X7 U442 ( .A(dma_rdata[61]), .B(n144), .Z(n848) );
  HS65_LS_BFX9 U443 ( .A(n869), .Z(n298) );
  HS65_LS_NOR3AX2 U444 ( .A(phitIn[34]), .B(phitIn[32]), .C(phitIn[33]), .Z(
        n869) );
  HS65_LS_AO22X9 U445 ( .A(n868), .B(address[0]), .C(phitIn[17]), .D(n653), 
        .Z(n743) );
  HS65_LS_AO22X9 U446 ( .A(n868), .B(address[1]), .C(phitIn[18]), .D(n653), 
        .Z(n741) );
  HS65_LS_AO22X9 U447 ( .A(n868), .B(address[2]), .C(phitIn[19]), .D(n653), 
        .Z(n739) );
  HS65_LS_AO22X9 U448 ( .A(n868), .B(address[3]), .C(phitIn[20]), .D(n653), 
        .Z(n737) );
  HS65_LS_AO22X9 U449 ( .A(n868), .B(address[4]), .C(phitIn[21]), .D(n653), 
        .Z(n735) );
  HS65_LS_AO22X9 U450 ( .A(n868), .B(address[5]), .C(phitIn[22]), .D(n653), 
        .Z(n733) );
  HS65_LS_AO22X9 U451 ( .A(n868), .B(address[6]), .C(phitIn[23]), .D(n653), 
        .Z(n731) );
  HS65_LS_IVX9 U452 ( .A(slt_entry[3]), .Z(n650) );
  HS65_LS_IVX9 U453 ( .A(slt_entry[2]), .Z(n651) );
  HS65_LS_AO22X9 U454 ( .A(phitIn[0]), .B(n312), .C(\spm_out[MDATA][0] ), .D(
        n306), .Z(n832) );
  HS65_LS_AO22X9 U455 ( .A(phitIn[1]), .B(n323), .C(\spm_out[MDATA][1] ), .D(
        n306), .Z(n831) );
  HS65_LS_AO22X9 U456 ( .A(phitIn[2]), .B(n323), .C(\spm_out[MDATA][2] ), .D(
        n306), .Z(n830) );
  HS65_LS_AO22X9 U457 ( .A(phitIn[3]), .B(n323), .C(\spm_out[MDATA][3] ), .D(
        n305), .Z(n829) );
  HS65_LS_AO22X9 U458 ( .A(phitIn[4]), .B(n323), .C(\spm_out[MDATA][4] ), .D(
        n304), .Z(n828) );
  HS65_LS_AO22X9 U459 ( .A(phitIn[5]), .B(n323), .C(\spm_out[MDATA][5] ), .D(
        n870), .Z(n827) );
  HS65_LS_AO22X9 U460 ( .A(phitIn[6]), .B(n323), .C(\spm_out[MDATA][6] ), .D(
        n306), .Z(n826) );
  HS65_LS_AO22X9 U461 ( .A(phitIn[7]), .B(n323), .C(\spm_out[MDATA][7] ), .D(
        n870), .Z(n825) );
  HS65_LS_AO22X9 U462 ( .A(phitIn[8]), .B(n323), .C(\spm_out[MDATA][8] ), .D(
        n870), .Z(n824) );
  HS65_LS_AO22X9 U463 ( .A(phitIn[9]), .B(n323), .C(\spm_out[MDATA][9] ), .D(
        n870), .Z(n823) );
  HS65_LS_AO22X9 U464 ( .A(phitIn[10]), .B(n314), .C(\spm_out[MDATA][10] ), 
        .D(n870), .Z(n822) );
  HS65_LS_AO22X9 U465 ( .A(phitIn[11]), .B(n314), .C(\spm_out[MDATA][11] ), 
        .D(n870), .Z(n821) );
  HS65_LS_AO22X9 U466 ( .A(phitIn[12]), .B(n314), .C(\spm_out[MDATA][12] ), 
        .D(n870), .Z(n820) );
  HS65_LS_AO22X9 U467 ( .A(phitIn[13]), .B(n314), .C(\spm_out[MDATA][13] ), 
        .D(n870), .Z(n819) );
  HS65_LS_AO22X9 U468 ( .A(phitIn[14]), .B(n314), .C(\spm_out[MDATA][14] ), 
        .D(n870), .Z(n818) );
  HS65_LS_AO22X9 U469 ( .A(phitIn[15]), .B(n314), .C(\spm_out[MDATA][15] ), 
        .D(n870), .Z(n817) );
  HS65_LS_AO22X9 U470 ( .A(phitIn[16]), .B(n314), .C(\spm_out[MDATA][16] ), 
        .D(n870), .Z(n816) );
  HS65_LS_AO22X9 U471 ( .A(phitIn[17]), .B(n314), .C(\spm_out[MDATA][17] ), 
        .D(n870), .Z(n815) );
  HS65_LS_AO22X9 U472 ( .A(phitIn[18]), .B(n314), .C(\spm_out[MDATA][18] ), 
        .D(n870), .Z(n814) );
  HS65_LS_AO22X9 U473 ( .A(phitIn[19]), .B(n314), .C(\spm_out[MDATA][19] ), 
        .D(n306), .Z(n813) );
  HS65_LS_AO22X9 U474 ( .A(phitIn[20]), .B(n314), .C(\spm_out[MDATA][20] ), 
        .D(n306), .Z(n812) );
  HS65_LS_AO22X9 U475 ( .A(phitIn[21]), .B(n314), .C(\spm_out[MDATA][21] ), 
        .D(n306), .Z(n811) );
  HS65_LS_AO22X9 U476 ( .A(phitIn[22]), .B(n314), .C(\spm_out[MDATA][22] ), 
        .D(n306), .Z(n810) );
  HS65_LS_AO22X9 U477 ( .A(phitIn[23]), .B(n314), .C(\spm_out[MDATA][23] ), 
        .D(n306), .Z(n809) );
  HS65_LS_AO22X9 U478 ( .A(phitIn[24]), .B(n314), .C(\spm_out[MDATA][24] ), 
        .D(n306), .Z(n808) );
  HS65_LS_AO22X9 U479 ( .A(phitIn[25]), .B(n314), .C(\spm_out[MDATA][25] ), 
        .D(n306), .Z(n807) );
  HS65_LS_AO22X9 U480 ( .A(phitIn[26]), .B(n314), .C(\spm_out[MDATA][26] ), 
        .D(n306), .Z(n806) );
  HS65_LS_AO22X9 U481 ( .A(phitIn[27]), .B(n314), .C(\spm_out[MDATA][27] ), 
        .D(n306), .Z(n805) );
  HS65_LS_AO22X9 U482 ( .A(phitIn[28]), .B(n314), .C(\spm_out[MDATA][28] ), 
        .D(n306), .Z(n804) );
  HS65_LS_AO22X9 U483 ( .A(phitIn[29]), .B(n314), .C(\spm_out[MDATA][29] ), 
        .D(n306), .Z(n803) );
  HS65_LS_AO22X9 U484 ( .A(phitIn[30]), .B(n313), .C(\spm_out[MDATA][30] ), 
        .D(n306), .Z(n802) );
  HS65_LS_AO22X9 U485 ( .A(phitIn[31]), .B(n313), .C(\spm_out[MDATA][31] ), 
        .D(n306), .Z(n801) );
  HS65_LS_AO22X9 U486 ( .A(dIn_h[0]), .B(n313), .C(\spm_out[MDATA][32] ), .D(
        n305), .Z(n800) );
  HS65_LS_AO22X9 U487 ( .A(dIn_h[1]), .B(n313), .C(\spm_out[MDATA][33] ), .D(
        n305), .Z(n799) );
  HS65_LS_AO22X9 U488 ( .A(dIn_h[2]), .B(n313), .C(\spm_out[MDATA][34] ), .D(
        n305), .Z(n798) );
  HS65_LS_AO22X9 U489 ( .A(dIn_h[3]), .B(n313), .C(\spm_out[MDATA][35] ), .D(
        n305), .Z(n797) );
  HS65_LS_AO22X9 U490 ( .A(dIn_h[4]), .B(n313), .C(\spm_out[MDATA][36] ), .D(
        n305), .Z(n796) );
  HS65_LS_AO22X9 U491 ( .A(dIn_h[5]), .B(n313), .C(\spm_out[MDATA][37] ), .D(
        n305), .Z(n795) );
  HS65_LS_AO22X9 U492 ( .A(dIn_h[6]), .B(n313), .C(\spm_out[MDATA][38] ), .D(
        n305), .Z(n794) );
  HS65_LS_AO22X9 U493 ( .A(dIn_h[7]), .B(n313), .C(\spm_out[MDATA][39] ), .D(
        n305), .Z(n793) );
  HS65_LS_AO22X9 U494 ( .A(dIn_h[8]), .B(n313), .C(\spm_out[MDATA][40] ), .D(
        n305), .Z(n792) );
  HS65_LS_AO22X9 U495 ( .A(dIn_h[9]), .B(n313), .C(\spm_out[MDATA][41] ), .D(
        n305), .Z(n791) );
  HS65_LS_AO22X9 U496 ( .A(dIn_h[10]), .B(n313), .C(\spm_out[MDATA][42] ), .D(
        n305), .Z(n790) );
  HS65_LS_AO22X9 U497 ( .A(dIn_h[11]), .B(n313), .C(\spm_out[MDATA][43] ), .D(
        n305), .Z(n789) );
  HS65_LS_AO22X9 U498 ( .A(dIn_h[12]), .B(n313), .C(\spm_out[MDATA][44] ), .D(
        n304), .Z(n788) );
  HS65_LS_AO22X9 U499 ( .A(dIn_h[13]), .B(n313), .C(\spm_out[MDATA][45] ), .D(
        n304), .Z(n787) );
  HS65_LS_AO22X9 U500 ( .A(dIn_h[14]), .B(n313), .C(\spm_out[MDATA][46] ), .D(
        n304), .Z(n786) );
  HS65_LS_AO22X9 U501 ( .A(dIn_h[15]), .B(n313), .C(\spm_out[MDATA][47] ), .D(
        n304), .Z(n785) );
  HS65_LS_AO22X9 U502 ( .A(dIn_h[16]), .B(n313), .C(\spm_out[MDATA][48] ), .D(
        n304), .Z(n784) );
  HS65_LS_AO22X9 U503 ( .A(dIn_h[17]), .B(n312), .C(\spm_out[MDATA][49] ), .D(
        n304), .Z(n783) );
  HS65_LS_AO22X9 U504 ( .A(dIn_h[18]), .B(n312), .C(\spm_out[MDATA][50] ), .D(
        n304), .Z(n782) );
  HS65_LS_AO22X9 U505 ( .A(dIn_h[19]), .B(n312), .C(\spm_out[MDATA][51] ), .D(
        n304), .Z(n781) );
  HS65_LS_AO22X9 U506 ( .A(dIn_h[20]), .B(n313), .C(\spm_out[MDATA][52] ), .D(
        n304), .Z(n780) );
  HS65_LS_AO22X9 U507 ( .A(dIn_h[21]), .B(n312), .C(\spm_out[MDATA][53] ), .D(
        n305), .Z(n779) );
  HS65_LS_AO22X9 U508 ( .A(dIn_h[22]), .B(n312), .C(\spm_out[MDATA][54] ), .D(
        n304), .Z(n778) );
  HS65_LS_AO22X9 U509 ( .A(dIn_h[23]), .B(n312), .C(\spm_out[MDATA][55] ), .D(
        n304), .Z(n777) );
  HS65_LS_AO22X9 U510 ( .A(dIn_h[24]), .B(n312), .C(\spm_out[MDATA][56] ), .D(
        n304), .Z(n776) );
  HS65_LS_AO22X9 U511 ( .A(dIn_h[25]), .B(n312), .C(\spm_out[MDATA][57] ), .D(
        n304), .Z(n775) );
  HS65_LS_AO22X9 U512 ( .A(dIn_h[26]), .B(n312), .C(\spm_out[MDATA][58] ), .D(
        n304), .Z(n774) );
  HS65_LS_AO22X9 U513 ( .A(dIn_h[27]), .B(n312), .C(\spm_out[MDATA][59] ), .D(
        n305), .Z(n773) );
  HS65_LS_AO22X9 U514 ( .A(dIn_h[28]), .B(n312), .C(\spm_out[MDATA][60] ), .D(
        n304), .Z(n772) );
  HS65_LS_AO22X9 U515 ( .A(dIn_h[29]), .B(n312), .C(\spm_out[MDATA][61] ), .D(
        n305), .Z(n771) );
  HS65_LS_AO22X9 U516 ( .A(dIn_h[30]), .B(n312), .C(\spm_out[MDATA][62] ), .D(
        n304), .Z(n770) );
  HS65_LS_AO22X9 U517 ( .A(dIn_h[31]), .B(n312), .C(\spm_out[MDATA][63] ), .D(
        n306), .Z(n769) );
  HS65_LS_AO22X9 U518 ( .A(phitIn[17]), .B(n302), .C(n300), .D(dIn_h[17]), .Z(
        n744) );
  HS65_LS_AO22X9 U519 ( .A(phitIn[18]), .B(n302), .C(n300), .D(dIn_h[18]), .Z(
        n742) );
  HS65_LS_AO22X9 U520 ( .A(phitIn[19]), .B(n302), .C(n300), .D(dIn_h[19]), .Z(
        n740) );
  HS65_LS_AO22X9 U521 ( .A(phitIn[20]), .B(n302), .C(n300), .D(dIn_h[20]), .Z(
        n738) );
  HS65_LS_AO22X9 U522 ( .A(phitIn[21]), .B(n303), .C(n300), .D(dIn_h[21]), .Z(
        n736) );
  HS65_LS_AO22X9 U523 ( .A(phitIn[22]), .B(n303), .C(n300), .D(dIn_h[22]), .Z(
        n734) );
  HS65_LS_AO22X9 U524 ( .A(phitIn[23]), .B(n303), .C(n300), .D(dIn_h[23]), .Z(
        n732) );
  HS65_LS_AO22X9 U525 ( .A(phitIn[0]), .B(n301), .C(n299), .D(dIn_h[0]), .Z(
        n761) );
  HS65_LS_AO22X9 U526 ( .A(phitIn[1]), .B(n302), .C(n299), .D(dIn_h[1]), .Z(
        n760) );
  HS65_LS_AO22X9 U527 ( .A(phitIn[2]), .B(n302), .C(n299), .D(dIn_h[2]), .Z(
        n759) );
  HS65_LS_AO22X9 U528 ( .A(phitIn[3]), .B(n302), .C(n299), .D(dIn_h[3]), .Z(
        n758) );
  HS65_LS_AO22X9 U529 ( .A(phitIn[4]), .B(n302), .C(n299), .D(dIn_h[4]), .Z(
        n757) );
  HS65_LS_AO22X9 U530 ( .A(phitIn[5]), .B(n302), .C(n299), .D(dIn_h[5]), .Z(
        n756) );
  HS65_LS_AO22X9 U531 ( .A(phitIn[6]), .B(n302), .C(n299), .D(dIn_h[6]), .Z(
        n755) );
  HS65_LS_AO22X9 U532 ( .A(phitIn[7]), .B(n302), .C(n299), .D(dIn_h[7]), .Z(
        n754) );
  HS65_LS_AO22X9 U533 ( .A(phitIn[8]), .B(n302), .C(n299), .D(dIn_h[8]), .Z(
        n753) );
  HS65_LS_AO22X9 U534 ( .A(phitIn[9]), .B(n302), .C(n299), .D(dIn_h[9]), .Z(
        n752) );
  HS65_LS_AO22X9 U535 ( .A(phitIn[10]), .B(n302), .C(n299), .D(dIn_h[10]), .Z(
        n751) );
  HS65_LS_AO22X9 U536 ( .A(phitIn[11]), .B(n302), .C(n299), .D(dIn_h[11]), .Z(
        n750) );
  HS65_LS_AO22X9 U537 ( .A(phitIn[12]), .B(n302), .C(n299), .D(dIn_h[12]), .Z(
        n749) );
  HS65_LS_AO22X9 U538 ( .A(phitIn[13]), .B(n302), .C(n300), .D(dIn_h[13]), .Z(
        n748) );
  HS65_LS_AO22X9 U539 ( .A(phitIn[14]), .B(n302), .C(n300), .D(dIn_h[14]), .Z(
        n747) );
  HS65_LS_AO22X9 U540 ( .A(phitIn[15]), .B(n302), .C(n300), .D(dIn_h[15]), .Z(
        n746) );
  HS65_LS_AO22X9 U541 ( .A(phitIn[16]), .B(n302), .C(n300), .D(dIn_h[16]), .Z(
        n745) );
  HS65_LS_AO22X9 U542 ( .A(phitIn[24]), .B(n303), .C(n300), .D(dIn_h[24]), .Z(
        n730) );
  HS65_LS_AO22X9 U543 ( .A(phitIn[25]), .B(n303), .C(n300), .D(dIn_h[25]), .Z(
        n729) );
  HS65_LS_AO22X9 U544 ( .A(phitIn[26]), .B(n303), .C(n299), .D(dIn_h[26]), .Z(
        n728) );
  HS65_LS_AO22X9 U545 ( .A(phitIn[27]), .B(n303), .C(n300), .D(dIn_h[27]), .Z(
        n727) );
  HS65_LS_AO22X9 U546 ( .A(phitIn[28]), .B(n303), .C(n299), .D(dIn_h[28]), .Z(
        n726) );
  HS65_LS_AO22X9 U547 ( .A(phitIn[29]), .B(n303), .C(n300), .D(dIn_h[29]), .Z(
        n725) );
  HS65_LS_AO22X9 U548 ( .A(phitIn[30]), .B(n303), .C(n299), .D(dIn_h[30]), .Z(
        n724) );
  HS65_LS_AO22X9 U549 ( .A(phitIn[31]), .B(n303), .C(n300), .D(dIn_h[31]), .Z(
        n723) );
  HS65_LS_AO22X9 U550 ( .A(n312), .B(address[0]), .C(n305), .D(flit_buf[64]), 
        .Z(n768) );
  HS65_LS_AO22X9 U551 ( .A(n312), .B(address[1]), .C(n304), .D(flit_buf[65]), 
        .Z(n767) );
  HS65_LS_AO22X9 U552 ( .A(n312), .B(address[2]), .C(n305), .D(flit_buf[66]), 
        .Z(n766) );
  HS65_LS_AO22X9 U553 ( .A(n312), .B(address[3]), .C(n304), .D(flit_buf[67]), 
        .Z(n765) );
  HS65_LS_AO22X9 U554 ( .A(n311), .B(address[4]), .C(n305), .D(flit_buf[68]), 
        .Z(n764) );
  HS65_LS_AO22X9 U555 ( .A(n310), .B(address[5]), .C(n304), .D(flit_buf[69]), 
        .Z(n763) );
  HS65_LS_AO22X9 U556 ( .A(n312), .B(address[6]), .C(n305), .D(flit_buf[70]), 
        .Z(n762) );
  HS65_LS_OR2X9 U557 ( .A(vld_pkt), .B(n653), .Z(n684) );
  HS65_LS_NAND2X7 U558 ( .A(\proc_in[MADDR][0] ), .B(n836), .Z(n861) );
  HS65_LS_NOR4ABX2 U559 ( .A(n660), .B(n833), .C(\proc_in[MADDR][26] ), .D(
        \proc_in[MADDR][24] ), .Z(n860) );
  HS65_LS_IVX9 U560 ( .A(\proc_in[MADDR][25] ), .Z(n660) );
  HS65_LS_NOR3X4 U561 ( .A(\proc_in[MADDR][27] ), .B(\proc_in[MADDR][31] ), 
        .C(\proc_in[MADDR][30] ), .Z(n833) );
  HS65_LS_NAND4ABX3 U562 ( .A(\proc_in[MADDR][29] ), .B(\proc_in[MADDR][26] ), 
        .C(n835), .D(n834), .Z(n858) );
  HS65_LS_NOR2X6 U563 ( .A(\proc_in[MADDR][31] ), .B(\proc_in[MADDR][30] ), 
        .Z(n835) );
  HS65_LS_NOR4ABX2 U564 ( .A(\proc_in[MADDR][28] ), .B(\proc_in[MADDR][27] ), 
        .C(\proc_in[MADDR][25] ), .D(\proc_in[MADDR][24] ), .Z(n834) );
  HS65_LS_NOR3AX2 U565 ( .A(n860), .B(n659), .C(\proc_in[MADDR][29] ), .Z(n680) );
  HS65_LS_NAND4ABX3 U566 ( .A(config_reg[3]), .B(n874), .C(config_reg[4]), .D(
        n597), .Z(n875) );
  HS65_LS_OA32X4 U567 ( .A(config_reg[0]), .B(config_reg[1]), .C(n654), .D(
        n873), .E(config_reg[2]), .Z(n874) );
  HS65_LS_IVX9 U568 ( .A(config_reg[2]), .Z(n654) );
  HS65_LSS_XNOR2X6 U569 ( .A(config_reg[1]), .B(config_reg[0]), .Z(n873) );
  HS65_LS_BFX9 U570 ( .A(na_reset), .Z(n339) );
  HS65_LS_BFX9 U571 ( .A(na_reset), .Z(n340) );
  HS65_LS_NAND2X7 U572 ( .A(n680), .B(\proc_in[MCMD][0] ), .Z(n872) );
  HS65_LS_IVX9 U573 ( .A(\proc_in[MDATA][15] ), .Z(n664) );
  HS65_LS_IVX9 U574 ( .A(\proc_in[MDATA][6] ), .Z(n673) );
  HS65_LS_IVX9 U575 ( .A(\proc_in[MDATA][7] ), .Z(n672) );
  HS65_LS_IVX9 U576 ( .A(\proc_in[MDATA][8] ), .Z(n671) );
  HS65_LS_IVX9 U577 ( .A(\proc_in[MDATA][9] ), .Z(n670) );
  HS65_LS_IVX9 U578 ( .A(\proc_in[MADDR][28] ), .Z(n659) );
  HS65_LS_AND3X9 U579 ( .A(n860), .B(n659), .C(\proc_in[MADDR][29] ), .Z(n836)
         );
  HS65_LS_IVX9 U580 ( .A(\proc_in[MDATA][14] ), .Z(n665) );
  HS65_LS_IVX9 U581 ( .A(\proc_in[MDATA][0] ), .Z(n679) );
  HS65_LS_IVX9 U582 ( .A(\proc_in[MDATA][1] ), .Z(n678) );
  HS65_LS_IVX9 U583 ( .A(\proc_in[MDATA][2] ), .Z(n677) );
  HS65_LS_IVX9 U584 ( .A(\proc_in[MDATA][3] ), .Z(n676) );
  HS65_LS_IVX9 U585 ( .A(\proc_in[MDATA][4] ), .Z(n675) );
  HS65_LS_IVX9 U586 ( .A(\proc_in[MDATA][5] ), .Z(n674) );
  HS65_LS_IVX9 U587 ( .A(\proc_in[MDATA][10] ), .Z(n669) );
  HS65_LS_IVX9 U588 ( .A(\proc_in[MDATA][11] ), .Z(n668) );
  HS65_LS_IVX9 U589 ( .A(\proc_in[MDATA][12] ), .Z(n667) );
  HS65_LS_IVX9 U590 ( .A(\proc_in[MDATA][13] ), .Z(n666) );
  HS65_LS_IVX9 U591 ( .A(\proc_in[MADDR][0] ), .Z(n663) );
  HS65_LS_IVX9 U592 ( .A(\proc_in[MADDR][1] ), .Z(n662) );
  HS65_LS_IVX9 U593 ( .A(n17), .Z(n517) );
  HS65_LS_IVX18 U594 ( .A(n469), .Z(n471) );
  HS65_LH_MUX21I1X3 U595 ( .D0(n20), .D1(n455), .S0(n652), .Z(n687) );
  HS65_LS_IVX9 U596 ( .A(n142), .Z(n128) );
  HS65_LH_BFX2 U597 ( .A(n139), .Z(n142) );
  HS65_LS_NAND2X5 U598 ( .A(n448), .B(n19), .Z(n449) );
  HS65_LS_AOI33X5 U599 ( .A(phitOut2[34]), .B(n468), .C(n578), .D(n578), .E(
        n577), .F(phitOut0[34]), .Z(n579) );
  HS65_LS_NAND2X5 U600 ( .A(phitOut2[13]), .B(n25), .Z(n511) );
  HS65_LS_NAND2X5 U601 ( .A(phitOut2[17]), .B(n25), .Z(n524) );
  HS65_LS_NAND2X7 U602 ( .A(phitOut2[18]), .B(n517), .Z(n527) );
  HS65_LS_AND2X4 U603 ( .A(n27), .B(n415), .Z(phit_togo[32]) );
  HS65_LH_CBI4I1X3 U604 ( .A(n128), .B(n364), .C(n306), .D(n363), .Z(n685) );
  HS65_LS_AO33X9 U605 ( .A(n120), .B(n5), .C(n453), .D(\phase_next[1] ), .E(
        n451), .F(n450), .Z(n470) );
  HS65_LS_IVX9 U606 ( .A(n451), .Z(n652) );
  HS65_LS_IVX9 U607 ( .A(n856), .Z(n625) );
  HS65_LS_NAND2X7 U608 ( .A(dma_rdata[39]), .B(n149), .Z(n595) );
  HS65_LS_IVX9 U609 ( .A(n595), .Z(n624) );
  HS65_LS_NAND2X7 U610 ( .A(dma_rdata[38]), .B(n149), .Z(n593) );
  HS65_LS_IVX9 U611 ( .A(n593), .Z(n623) );
  HS65_LS_NAND2X7 U612 ( .A(dma_rdata[37]), .B(n293), .Z(n591) );
  HS65_LS_IVX9 U613 ( .A(n591), .Z(n622) );
  HS65_LS_NAND2X7 U614 ( .A(dma_rdata[36]), .B(n293), .Z(n589) );
  HS65_LS_IVX9 U615 ( .A(n589), .Z(n621) );
  HS65_LS_NAND2X7 U616 ( .A(dma_rdata[35]), .B(n293), .Z(n587) );
  HS65_LS_IVX9 U617 ( .A(n587), .Z(n620) );
  HS65_LS_NAND2X7 U618 ( .A(dma_rdata[34]), .B(n293), .Z(n585) );
  HS65_LS_IVX9 U619 ( .A(n585), .Z(n619) );
  HS65_LS_NAND2X7 U620 ( .A(dma_rdata[33]), .B(n293), .Z(n583) );
  HS65_LS_IVX9 U621 ( .A(n583), .Z(n618) );
  HS65_LS_NAND2X7 U622 ( .A(dma_rdata[31]), .B(n293), .Z(n413) );
  HS65_LS_IVX9 U623 ( .A(n413), .Z(n617) );
  HS65_LS_NAND2X7 U624 ( .A(dma_rdata[30]), .B(n293), .Z(n411) );
  HS65_LS_IVX9 U625 ( .A(n411), .Z(n616) );
  HS65_LS_NAND2X7 U626 ( .A(dma_rdata[29]), .B(n293), .Z(n409) );
  HS65_LS_IVX9 U627 ( .A(n409), .Z(n615) );
  HS65_LS_NAND2X7 U628 ( .A(dma_rdata[28]), .B(n293), .Z(n407) );
  HS65_LS_IVX9 U629 ( .A(n407), .Z(n614) );
  HS65_LS_NAND2X7 U630 ( .A(dma_rdata[27]), .B(n293), .Z(n405) );
  HS65_LS_IVX9 U631 ( .A(n405), .Z(n613) );
  HS65_LS_NAND2X7 U632 ( .A(dma_rdata[26]), .B(n293), .Z(n403) );
  HS65_LS_IVX9 U633 ( .A(n403), .Z(n612) );
  HS65_LS_NAND2X7 U634 ( .A(dma_rdata[25]), .B(n293), .Z(n401) );
  HS65_LS_IVX9 U635 ( .A(n401), .Z(n611) );
  HS65_LS_NAND2X7 U636 ( .A(dma_rdata[24]), .B(n293), .Z(n399) );
  HS65_LS_IVX9 U637 ( .A(n399), .Z(n610) );
  HS65_LS_NAND2X7 U638 ( .A(dma_rdata[23]), .B(n293), .Z(n397) );
  HS65_LS_IVX9 U639 ( .A(n397), .Z(n609) );
  HS65_LS_NAND2X7 U640 ( .A(dma_rdata[22]), .B(n293), .Z(n395) );
  HS65_LS_IVX9 U641 ( .A(n395), .Z(n608) );
  HS65_LS_NAND2X7 U642 ( .A(dma_rdata[21]), .B(n293), .Z(n393) );
  HS65_LS_IVX9 U643 ( .A(n393), .Z(n607) );
  HS65_LS_NAND2X7 U644 ( .A(dma_rdata[20]), .B(n293), .Z(n391) );
  HS65_LS_IVX9 U645 ( .A(n391), .Z(n606) );
  HS65_LS_NAND2X7 U646 ( .A(dma_rdata[19]), .B(n149), .Z(n389) );
  HS65_LS_IVX9 U647 ( .A(n389), .Z(n605) );
  HS65_LS_NAND2X7 U648 ( .A(dma_rdata[18]), .B(n149), .Z(n387) );
  HS65_LS_IVX9 U649 ( .A(n387), .Z(n604) );
  HS65_LS_NAND2X7 U650 ( .A(dma_rdata[17]), .B(n149), .Z(n385) );
  HS65_LS_IVX9 U651 ( .A(n385), .Z(n603) );
  HS65_LS_IVX9 U652 ( .A(\proc_in[MCMD][0] ), .Z(n360) );
  HS65_LS_IVX9 U653 ( .A(n362), .Z(n361) );
  HS65_LS_NAND2X7 U654 ( .A(n839), .B(n1), .Z(n857) );
  HS65_LS_OAI22X6 U655 ( .A(n650), .B(n365), .C(n838), .D(n362), .Z(
        dma_raddr[1]) );
  HS65_LS_OAI22X6 U656 ( .A(n651), .B(n365), .C(n837), .D(n362), .Z(
        dma_raddr[0]) );
  HS65_LS_NAND2X7 U657 ( .A(dma_rdata[16]), .B(n149), .Z(n383) );
  HS65_LS_IVX9 U658 ( .A(n383), .Z(n600) );
  HS65_LS_IVX9 U659 ( .A(n690), .Z(n455) );
  HS65_LS_IVX9 U660 ( .A(vld_pkt), .Z(n364) );
  HS65_LS_IVX9 U661 ( .A(n688), .Z(n581) );
  HS65_LS_IVX9 U662 ( .A(n365), .Z(n602) );
  HS65_LS_IVX9 U663 ( .A(n689), .Z(n415) );
  HS65_LS_NAND2X7 U664 ( .A(n602), .B(n415), .Z(n414) );
  HS65_LS_IVX9 U665 ( .A(dOut_l[0]), .Z(n416) );
  HS65_LS_NAND2X7 U666 ( .A(\spm_in[SDATA][32] ), .B(n130), .Z(n366) );
  HS65_LS_OAI212X5 U667 ( .A(n136), .B(n416), .C(n329), .D(n647), .E(n366), 
        .Z(mux_out[0]) );
  HS65_LS_IVX9 U668 ( .A(dOut_l[1]), .Z(n417) );
  HS65_LS_NAND2X7 U669 ( .A(\spm_in[SDATA][33] ), .B(n130), .Z(n367) );
  HS65_LS_OAI212X5 U670 ( .A(n136), .B(n417), .C(n329), .D(n646), .E(n367), 
        .Z(mux_out[1]) );
  HS65_LS_IVX9 U671 ( .A(dOut_l[2]), .Z(n418) );
  HS65_LS_NAND2X7 U672 ( .A(\spm_in[SDATA][34] ), .B(n130), .Z(n368) );
  HS65_LS_OAI212X5 U673 ( .A(n136), .B(n418), .C(n329), .D(n645), .E(n368), 
        .Z(mux_out[2]) );
  HS65_LS_IVX9 U674 ( .A(dOut_l[3]), .Z(n419) );
  HS65_LS_NAND2X7 U675 ( .A(\spm_in[SDATA][35] ), .B(n130), .Z(n369) );
  HS65_LS_OAI212X5 U676 ( .A(n136), .B(n419), .C(n329), .D(n644), .E(n369), 
        .Z(mux_out[3]) );
  HS65_LS_IVX9 U677 ( .A(dOut_l[4]), .Z(n420) );
  HS65_LS_NAND2X7 U678 ( .A(\spm_in[SDATA][36] ), .B(n130), .Z(n370) );
  HS65_LS_OAI212X5 U679 ( .A(n136), .B(n420), .C(n329), .D(n643), .E(n370), 
        .Z(mux_out[4]) );
  HS65_LS_IVX9 U680 ( .A(dOut_l[5]), .Z(n421) );
  HS65_LS_NAND2X7 U681 ( .A(\spm_in[SDATA][37] ), .B(n130), .Z(n371) );
  HS65_LS_OAI212X5 U682 ( .A(n136), .B(n421), .C(n329), .D(n642), .E(n371), 
        .Z(mux_out[5]) );
  HS65_LS_IVX9 U683 ( .A(dOut_l[6]), .Z(n422) );
  HS65_LS_NAND2X7 U684 ( .A(\spm_in[SDATA][38] ), .B(n130), .Z(n372) );
  HS65_LS_OAI212X5 U685 ( .A(n136), .B(n422), .C(n329), .D(n641), .E(n372), 
        .Z(mux_out[6]) );
  HS65_LS_IVX9 U686 ( .A(dOut_l[7]), .Z(n423) );
  HS65_LS_NAND2X7 U687 ( .A(\spm_in[SDATA][39] ), .B(n130), .Z(n373) );
  HS65_LS_OAI212X5 U688 ( .A(n136), .B(n423), .C(n329), .D(n640), .E(n373), 
        .Z(mux_out[7]) );
  HS65_LS_IVX9 U689 ( .A(dOut_l[8]), .Z(n424) );
  HS65_LS_NAND2X7 U690 ( .A(\spm_in[SDATA][40] ), .B(n130), .Z(n374) );
  HS65_LS_OAI212X5 U691 ( .A(n136), .B(n424), .C(n329), .D(n639), .E(n374), 
        .Z(mux_out[8]) );
  HS65_LS_IVX9 U692 ( .A(dOut_l[9]), .Z(n425) );
  HS65_LS_NAND2X7 U693 ( .A(\spm_in[SDATA][41] ), .B(n130), .Z(n375) );
  HS65_LS_OAI212X5 U694 ( .A(n136), .B(n425), .C(n328), .D(n638), .E(n375), 
        .Z(mux_out[9]) );
  HS65_LS_IVX9 U695 ( .A(dOut_l[10]), .Z(n426) );
  HS65_LS_NAND2X7 U696 ( .A(\spm_in[SDATA][42] ), .B(n130), .Z(n376) );
  HS65_LS_OAI212X5 U697 ( .A(n136), .B(n426), .C(n328), .D(n637), .E(n376), 
        .Z(mux_out[10]) );
  HS65_LS_IVX9 U698 ( .A(dOut_l[11]), .Z(n427) );
  HS65_LS_NAND2X7 U699 ( .A(\spm_in[SDATA][43] ), .B(n130), .Z(n377) );
  HS65_LS_OAI212X5 U700 ( .A(n136), .B(n427), .C(n328), .D(n636), .E(n377), 
        .Z(mux_out[11]) );
  HS65_LS_IVX9 U701 ( .A(dOut_l[12]), .Z(n428) );
  HS65_LS_NAND2X7 U702 ( .A(\spm_in[SDATA][44] ), .B(n132), .Z(n378) );
  HS65_LS_OAI212X5 U703 ( .A(n137), .B(n428), .C(n328), .D(n635), .E(n378), 
        .Z(mux_out[12]) );
  HS65_LS_IVX9 U704 ( .A(dOut_l[13]), .Z(n429) );
  HS65_LS_NAND2X7 U705 ( .A(\spm_in[SDATA][45] ), .B(n132), .Z(n379) );
  HS65_LS_OAI212X5 U706 ( .A(n137), .B(n429), .C(n328), .D(n634), .E(n379), 
        .Z(mux_out[13]) );
  HS65_LS_IVX9 U707 ( .A(dOut_l[14]), .Z(n430) );
  HS65_LS_NAND2X7 U708 ( .A(\spm_in[SDATA][46] ), .B(n132), .Z(n380) );
  HS65_LS_OAI212X5 U709 ( .A(n137), .B(n430), .C(n328), .D(n633), .E(n380), 
        .Z(mux_out[14]) );
  HS65_LS_IVX9 U710 ( .A(dOut_l[15]), .Z(n431) );
  HS65_LS_NAND2X7 U711 ( .A(\spm_in[SDATA][47] ), .B(n132), .Z(n381) );
  HS65_LS_OAI212X5 U712 ( .A(n137), .B(n431), .C(n328), .D(n632), .E(n381), 
        .Z(mux_out[15]) );
  HS65_LS_IVX9 U713 ( .A(dOut_l[16]), .Z(n432) );
  HS65_LS_NAND2X7 U714 ( .A(\spm_in[SDATA][48] ), .B(n132), .Z(n382) );
  HS65_LS_OAI212X5 U715 ( .A(n137), .B(n432), .C(n328), .D(n383), .E(n382), 
        .Z(mux_out[16]) );
  HS65_LS_IVX9 U716 ( .A(dOut_l[17]), .Z(n433) );
  HS65_LS_NAND2X7 U717 ( .A(\spm_in[SDATA][49] ), .B(n132), .Z(n384) );
  HS65_LS_OAI212X5 U718 ( .A(n137), .B(n433), .C(n328), .D(n385), .E(n384), 
        .Z(mux_out[17]) );
  HS65_LS_IVX9 U719 ( .A(dOut_l[18]), .Z(n434) );
  HS65_LS_NAND2X7 U720 ( .A(\spm_in[SDATA][50] ), .B(n132), .Z(n386) );
  HS65_LS_OAI212X5 U721 ( .A(n137), .B(n434), .C(n328), .D(n387), .E(n386), 
        .Z(mux_out[18]) );
  HS65_LS_IVX9 U722 ( .A(dOut_l[19]), .Z(n435) );
  HS65_LS_NAND2X7 U723 ( .A(\spm_in[SDATA][51] ), .B(n132), .Z(n388) );
  HS65_LS_OAI212X5 U724 ( .A(n137), .B(n435), .C(n328), .D(n389), .E(n388), 
        .Z(mux_out[19]) );
  HS65_LS_IVX9 U725 ( .A(dOut_l[20]), .Z(n436) );
  HS65_LS_NAND2X7 U726 ( .A(\spm_in[SDATA][52] ), .B(n132), .Z(n390) );
  HS65_LS_OAI212X5 U727 ( .A(n137), .B(n436), .C(n328), .D(n391), .E(n390), 
        .Z(mux_out[20]) );
  HS65_LS_IVX9 U728 ( .A(dOut_l[21]), .Z(n437) );
  HS65_LS_NAND2X7 U729 ( .A(\spm_in[SDATA][53] ), .B(n132), .Z(n392) );
  HS65_LS_OAI212X5 U730 ( .A(n137), .B(n437), .C(n328), .D(n393), .E(n392), 
        .Z(mux_out[21]) );
  HS65_LS_IVX9 U731 ( .A(dOut_l[22]), .Z(n438) );
  HS65_LS_NAND2X7 U732 ( .A(\spm_in[SDATA][54] ), .B(n132), .Z(n394) );
  HS65_LS_OAI212X5 U733 ( .A(n137), .B(n438), .C(n328), .D(n395), .E(n394), 
        .Z(mux_out[22]) );
  HS65_LS_IVX9 U734 ( .A(dOut_l[23]), .Z(n439) );
  HS65_LS_NAND2X7 U735 ( .A(\spm_in[SDATA][55] ), .B(n132), .Z(n396) );
  HS65_LS_OAI212X5 U736 ( .A(n137), .B(n439), .C(n328), .D(n397), .E(n396), 
        .Z(mux_out[23]) );
  HS65_LS_IVX9 U737 ( .A(dOut_l[24]), .Z(n440) );
  HS65_LS_NAND2X7 U738 ( .A(\spm_in[SDATA][56] ), .B(n133), .Z(n398) );
  HS65_LS_OAI212X5 U739 ( .A(n138), .B(n440), .C(n328), .D(n399), .E(n398), 
        .Z(mux_out[24]) );
  HS65_LS_IVX9 U740 ( .A(dOut_l[25]), .Z(n441) );
  HS65_LS_NAND2X7 U741 ( .A(\spm_in[SDATA][57] ), .B(n133), .Z(n400) );
  HS65_LS_OAI212X5 U742 ( .A(n138), .B(n441), .C(n328), .D(n401), .E(n400), 
        .Z(mux_out[25]) );
  HS65_LS_IVX9 U743 ( .A(dOut_l[26]), .Z(n442) );
  HS65_LS_NAND2X7 U744 ( .A(\spm_in[SDATA][58] ), .B(n133), .Z(n402) );
  HS65_LS_OAI212X5 U745 ( .A(n138), .B(n442), .C(n328), .D(n403), .E(n402), 
        .Z(mux_out[26]) );
  HS65_LS_IVX9 U746 ( .A(dOut_l[27]), .Z(n443) );
  HS65_LS_NAND2X7 U747 ( .A(\spm_in[SDATA][59] ), .B(n133), .Z(n404) );
  HS65_LS_OAI212X5 U748 ( .A(n138), .B(n443), .C(n327), .D(n405), .E(n404), 
        .Z(mux_out[27]) );
  HS65_LS_IVX9 U749 ( .A(dOut_l[28]), .Z(n444) );
  HS65_LS_NAND2X7 U750 ( .A(\spm_in[SDATA][60] ), .B(n133), .Z(n406) );
  HS65_LS_OAI212X5 U751 ( .A(n138), .B(n444), .C(n328), .D(n407), .E(n406), 
        .Z(mux_out[28]) );
  HS65_LS_IVX9 U752 ( .A(dOut_l[29]), .Z(n445) );
  HS65_LS_NAND2X7 U753 ( .A(\spm_in[SDATA][61] ), .B(n133), .Z(n408) );
  HS65_LS_OAI212X5 U754 ( .A(n138), .B(n445), .C(n327), .D(n409), .E(n408), 
        .Z(mux_out[29]) );
  HS65_LS_IVX9 U755 ( .A(dOut_l[30]), .Z(n446) );
  HS65_LS_NAND2X7 U756 ( .A(\spm_in[SDATA][62] ), .B(n133), .Z(n410) );
  HS65_LS_OAI212X5 U757 ( .A(n138), .B(n446), .C(n328), .D(n411), .E(n410), 
        .Z(mux_out[30]) );
  HS65_LS_IVX9 U758 ( .A(dOut_l[31]), .Z(n447) );
  HS65_LS_NAND2X7 U759 ( .A(\spm_in[SDATA][63] ), .B(n133), .Z(n412) );
  HS65_LS_OAI212X5 U760 ( .A(n138), .B(n447), .C(n327), .D(n413), .E(n412), 
        .Z(mux_out[31]) );
  HS65_LS_MUX21I1X6 U761 ( .D0(n416), .D1(\spm_in[SDATA][0] ), .S0(n140), .Z(
        n722) );
  HS65_LS_MUX21I1X6 U762 ( .D0(n417), .D1(\spm_in[SDATA][1] ), .S0(n140), .Z(
        n721) );
  HS65_LS_MUX21I1X6 U763 ( .D0(n418), .D1(\spm_in[SDATA][2] ), .S0(n140), .Z(
        n720) );
  HS65_LS_MUX21I1X6 U764 ( .D0(n419), .D1(\spm_in[SDATA][3] ), .S0(n142), .Z(
        n719) );
  HS65_LS_MUX21I1X6 U765 ( .D0(n420), .D1(\spm_in[SDATA][4] ), .S0(n140), .Z(
        n718) );
  HS65_LS_MUX21I1X6 U766 ( .D0(n421), .D1(\spm_in[SDATA][5] ), .S0(n142), .Z(
        n717) );
  HS65_LS_MUX21I1X6 U767 ( .D0(n422), .D1(\spm_in[SDATA][6] ), .S0(n34), .Z(
        n716) );
  HS65_LS_MUX21I1X6 U768 ( .D0(n423), .D1(\spm_in[SDATA][7] ), .S0(n140), .Z(
        n715) );
  HS65_LS_MUX21I1X6 U769 ( .D0(n424), .D1(\spm_in[SDATA][8] ), .S0(n140), .Z(
        n714) );
  HS65_LS_MUX21I1X6 U770 ( .D0(n425), .D1(\spm_in[SDATA][9] ), .S0(n140), .Z(
        n713) );
  HS65_LS_MUX21I1X6 U771 ( .D0(n426), .D1(\spm_in[SDATA][10] ), .S0(n34), .Z(
        n712) );
  HS65_LS_MUX21I1X6 U772 ( .D0(n427), .D1(\spm_in[SDATA][11] ), .S0(n140), .Z(
        n711) );
  HS65_LS_MUX21I1X6 U773 ( .D0(n428), .D1(\spm_in[SDATA][12] ), .S0(n34), .Z(
        n710) );
  HS65_LS_MUX21I1X6 U774 ( .D0(n429), .D1(\spm_in[SDATA][13] ), .S0(n34), .Z(
        n709) );
  HS65_LS_MUX21I1X6 U775 ( .D0(n430), .D1(\spm_in[SDATA][14] ), .S0(n34), .Z(
        n708) );
  HS65_LS_MUX21I1X6 U776 ( .D0(n431), .D1(\spm_in[SDATA][15] ), .S0(n34), .Z(
        n707) );
  HS65_LS_MUX21I1X6 U777 ( .D0(n432), .D1(\spm_in[SDATA][16] ), .S0(n34), .Z(
        n706) );
  HS65_LS_MUX21I1X6 U778 ( .D0(n433), .D1(\spm_in[SDATA][17] ), .S0(n140), .Z(
        n705) );
  HS65_LS_MUX21I1X6 U779 ( .D0(n434), .D1(\spm_in[SDATA][18] ), .S0(n34), .Z(
        n704) );
  HS65_LS_MUX21I1X6 U780 ( .D0(n435), .D1(\spm_in[SDATA][19] ), .S0(n140), .Z(
        n703) );
  HS65_LS_MUX21I1X6 U781 ( .D0(n436), .D1(\spm_in[SDATA][20] ), .S0(n34), .Z(
        n702) );
  HS65_LS_MUX21I1X6 U782 ( .D0(n437), .D1(\spm_in[SDATA][21] ), .S0(n140), .Z(
        n701) );
  HS65_LS_MUX21I1X6 U783 ( .D0(n438), .D1(\spm_in[SDATA][22] ), .S0(n142), .Z(
        n700) );
  HS65_LS_MUX21I1X6 U784 ( .D0(n439), .D1(\spm_in[SDATA][23] ), .S0(n34), .Z(
        n699) );
  HS65_LS_MUX21I1X6 U785 ( .D0(n440), .D1(\spm_in[SDATA][24] ), .S0(n140), .Z(
        n698) );
  HS65_LS_MUX21I1X6 U786 ( .D0(n441), .D1(\spm_in[SDATA][25] ), .S0(n34), .Z(
        n697) );
  HS65_LS_MUX21I1X6 U787 ( .D0(n442), .D1(\spm_in[SDATA][26] ), .S0(n34), .Z(
        n696) );
  HS65_LS_MUX21I1X6 U788 ( .D0(n443), .D1(\spm_in[SDATA][27] ), .S0(n140), .Z(
        n695) );
  HS65_LS_MUX21I1X6 U789 ( .D0(n444), .D1(\spm_in[SDATA][28] ), .S0(n34), .Z(
        n694) );
  HS65_LS_MUX21I1X6 U790 ( .D0(n445), .D1(\spm_in[SDATA][29] ), .S0(n140), .Z(
        n693) );
  HS65_LS_MUX21I1X6 U791 ( .D0(n446), .D1(\spm_in[SDATA][30] ), .S0(n34), .Z(
        n692) );
  HS65_LS_MUX21I1X6 U792 ( .D0(n447), .D1(\spm_in[SDATA][31] ), .S0(n140), .Z(
        n691) );
  HS65_LS_IVX9 U793 ( .A(\phase_next[1] ), .Z(n458) );
  HS65_LS_IVX9 U794 ( .A(n449), .Z(n465) );
  HS65_LS_NAND2X7 U795 ( .A(n27), .B(n461), .Z(n459) );
  HS65_LS_IVX9 U796 ( .A(n461), .Z(n464) );
  HS65_LS_IVX9 U797 ( .A(n462), .Z(n463) );
  HS65_LS_IVX9 U798 ( .A(phitOut1[0]), .Z(n475) );
  HS65_LS_IVX9 U799 ( .A(phitOut0[0]), .Z(n474) );
  HS65_LS_OAI212X5 U800 ( .A(n29), .B(n475), .C(n30), .D(n474), .E(n473), .Z(
        pkt_out[0]) );
  HS65_LS_IVX9 U801 ( .A(phitOut1[1]), .Z(n478) );
  HS65_LS_IVX9 U802 ( .A(phitOut0[1]), .Z(n477) );
  HS65_LS_OAI212X5 U803 ( .A(n22), .B(n478), .C(n30), .D(n477), .E(n476), .Z(
        pkt_out[1]) );
  HS65_LS_IVX9 U804 ( .A(phitOut1[2]), .Z(n480) );
  HS65_LS_IVX9 U805 ( .A(phitOut1[3]), .Z(n484) );
  HS65_LS_IVX9 U806 ( .A(phitOut0[3]), .Z(n483) );
  HS65_LS_NAND2X7 U807 ( .A(phitOut2[3]), .B(n572), .Z(n482) );
  HS65_LS_OAI212X5 U808 ( .A(n15), .B(n484), .C(n48), .D(n483), .E(n482), .Z(
        pkt_out[3]) );
  HS65_LS_IVX9 U809 ( .A(phitOut1[4]), .Z(n487) );
  HS65_LS_IVX9 U810 ( .A(phitOut0[4]), .Z(n486) );
  HS65_LS_OAI212X5 U811 ( .A(n22), .B(n487), .C(n48), .D(n486), .E(n485), .Z(
        pkt_out[4]) );
  HS65_LS_IVX9 U812 ( .A(phitOut1[5]), .Z(n490) );
  HS65_LS_IVX9 U813 ( .A(phitOut0[5]), .Z(n489) );
  HS65_LS_OAI212X5 U814 ( .A(n29), .B(n490), .C(n30), .D(n489), .E(n488), .Z(
        pkt_out[5]) );
  HS65_LS_IVX9 U815 ( .A(phitOut1[6]), .Z(n493) );
  HS65_LS_IVX9 U816 ( .A(phitOut0[6]), .Z(n492) );
  HS65_LS_NAND2X7 U817 ( .A(phitOut2[6]), .B(n572), .Z(n491) );
  HS65_LS_OAI212X5 U818 ( .A(n21), .B(n493), .C(n30), .D(n492), .E(n491), .Z(
        pkt_out[6]) );
  HS65_LS_IVX9 U819 ( .A(phitOut1[7]), .Z(n496) );
  HS65_LS_IVX9 U820 ( .A(phitOut0[7]), .Z(n495) );
  HS65_LS_OAI212X5 U821 ( .A(n29), .B(n496), .C(n30), .D(n495), .E(n494), .Z(
        pkt_out[7]) );
  HS65_LS_IVX9 U822 ( .A(phitOut1[8]), .Z(n499) );
  HS65_LS_IVX9 U823 ( .A(phitOut0[8]), .Z(n498) );
  HS65_LS_OAI212X5 U824 ( .A(n22), .B(n499), .C(n48), .D(n498), .E(n497), .Z(
        pkt_out[8]) );
  HS65_LS_IVX9 U825 ( .A(phitOut1[9]), .Z(n502) );
  HS65_LS_IVX9 U826 ( .A(phitOut0[9]), .Z(n501) );
  HS65_LS_NAND2X7 U827 ( .A(phitOut2[9]), .B(n572), .Z(n500) );
  HS65_LS_OAI212X5 U828 ( .A(n22), .B(n502), .C(n47), .D(n501), .E(n500), .Z(
        pkt_out[9]) );
  HS65_LS_IVX9 U829 ( .A(phitOut1[10]), .Z(n505) );
  HS65_LS_IVX9 U830 ( .A(phitOut0[10]), .Z(n504) );
  HS65_LS_NAND2X7 U831 ( .A(phitOut2[10]), .B(n572), .Z(n503) );
  HS65_LS_OAI212X5 U832 ( .A(n29), .B(n505), .C(n30), .D(n504), .E(n503), .Z(
        pkt_out[10]) );
  HS65_LS_IVX9 U833 ( .A(phitOut1[11]), .Z(n507) );
  HS65_LS_IVX9 U834 ( .A(phitOut1[12]), .Z(n510) );
  HS65_LS_IVX9 U835 ( .A(phitOut0[12]), .Z(n509) );
  HS65_LS_OAI212X5 U836 ( .A(n29), .B(n510), .C(n47), .D(n509), .E(n508), .Z(
        pkt_out[12]) );
  HS65_LS_IVX9 U837 ( .A(phitOut1[13]), .Z(n513) );
  HS65_LS_IVX9 U838 ( .A(phitOut0[13]), .Z(n512) );
  HS65_LS_OAI212X5 U839 ( .A(n22), .B(n513), .C(n48), .D(n512), .E(n511), .Z(
        pkt_out[13]) );
  HS65_LS_IVX9 U840 ( .A(phitOut1[14]), .Z(n516) );
  HS65_LS_IVX9 U841 ( .A(phitOut0[14]), .Z(n515) );
  HS65_LS_OAI212X5 U842 ( .A(n29), .B(n516), .C(n30), .D(n515), .E(n514), .Z(
        pkt_out[14]) );
  HS65_LS_IVX9 U843 ( .A(phitOut1[15]), .Z(n520) );
  HS65_LS_IVX9 U844 ( .A(phitOut0[15]), .Z(n519) );
  HS65_LS_OAI212X5 U845 ( .A(n22), .B(n520), .C(n30), .D(n519), .E(n518), .Z(
        pkt_out[15]) );
  HS65_LS_IVX9 U846 ( .A(phitOut1[16]), .Z(n523) );
  HS65_LS_IVX9 U847 ( .A(phitOut0[16]), .Z(n522) );
  HS65_LS_NAND2X7 U848 ( .A(phitOut2[16]), .B(n572), .Z(n521) );
  HS65_LS_OAI212X5 U849 ( .A(n29), .B(n523), .C(n47), .D(n522), .E(n521), .Z(
        pkt_out[16]) );
  HS65_LS_IVX9 U850 ( .A(phitOut1[17]), .Z(n526) );
  HS65_LS_IVX9 U851 ( .A(phitOut0[17]), .Z(n525) );
  HS65_LS_OAI212X5 U852 ( .A(n22), .B(n526), .C(n30), .D(n525), .E(n524), .Z(
        pkt_out[17]) );
  HS65_LS_IVX9 U853 ( .A(phitOut1[18]), .Z(n529) );
  HS65_LS_IVX9 U854 ( .A(phitOut0[18]), .Z(n528) );
  HS65_LS_OAI212X5 U855 ( .A(n22), .B(n529), .C(n47), .D(n528), .E(n527), .Z(
        pkt_out[18]) );
  HS65_LS_IVX9 U856 ( .A(phitOut1[19]), .Z(n532) );
  HS65_LS_IVX9 U857 ( .A(phitOut0[19]), .Z(n531) );
  HS65_LS_OAI212X5 U858 ( .A(n29), .B(n532), .C(n47), .D(n531), .E(n530), .Z(
        pkt_out[19]) );
  HS65_LS_IVX9 U859 ( .A(phitOut1[20]), .Z(n535) );
  HS65_LS_IVX9 U860 ( .A(phitOut0[20]), .Z(n534) );
  HS65_LS_NAND2X7 U861 ( .A(phitOut2[20]), .B(n572), .Z(n533) );
  HS65_LS_OAI212X5 U862 ( .A(n22), .B(n535), .C(n48), .D(n534), .E(n533), .Z(
        pkt_out[20]) );
  HS65_LS_IVX9 U863 ( .A(phitOut1[21]), .Z(n538) );
  HS65_LS_IVX9 U864 ( .A(phitOut0[21]), .Z(n537) );
  HS65_LS_OAI212X5 U865 ( .A(n15), .B(n538), .C(n48), .D(n537), .E(n536), .Z(
        pkt_out[21]) );
  HS65_LS_IVX9 U866 ( .A(phitOut1[22]), .Z(n541) );
  HS65_LS_IVX9 U867 ( .A(phitOut0[22]), .Z(n540) );
  HS65_LS_OAI212X5 U868 ( .A(n22), .B(n541), .C(n47), .D(n540), .E(n539), .Z(
        pkt_out[22]) );
  HS65_LS_IVX9 U869 ( .A(phitOut1[23]), .Z(n544) );
  HS65_LS_IVX9 U870 ( .A(phitOut0[23]), .Z(n543) );
  HS65_LS_OAI212X5 U871 ( .A(n22), .B(n544), .C(n47), .D(n543), .E(n542), .Z(
        pkt_out[23]) );
  HS65_LS_IVX9 U872 ( .A(phitOut1[24]), .Z(n547) );
  HS65_LS_IVX9 U873 ( .A(phitOut0[24]), .Z(n546) );
  HS65_LS_NAND2X7 U874 ( .A(phitOut2[24]), .B(n572), .Z(n545) );
  HS65_LS_OAI212X5 U875 ( .A(n22), .B(n547), .C(n47), .D(n546), .E(n545), .Z(
        pkt_out[24]) );
  HS65_LS_IVX9 U876 ( .A(phitOut1[25]), .Z(n550) );
  HS65_LS_IVX9 U877 ( .A(phitOut0[25]), .Z(n549) );
  HS65_LS_OAI212X5 U878 ( .A(n15), .B(n550), .C(n48), .D(n549), .E(n548), .Z(
        pkt_out[25]) );
  HS65_LS_IVX9 U879 ( .A(phitOut1[26]), .Z(n553) );
  HS65_LS_IVX9 U880 ( .A(phitOut0[26]), .Z(n552) );
  HS65_LS_NAND2X7 U881 ( .A(phitOut2[26]), .B(n517), .Z(n551) );
  HS65_LS_OAI212X5 U882 ( .A(n22), .B(n553), .C(n48), .D(n552), .E(n551), .Z(
        pkt_out[26]) );
  HS65_LS_IVX9 U883 ( .A(phitOut1[27]), .Z(n556) );
  HS65_LS_IVX9 U884 ( .A(phitOut0[27]), .Z(n555) );
  HS65_LS_OAI212X5 U885 ( .A(n15), .B(n556), .C(n48), .D(n555), .E(n554), .Z(
        pkt_out[27]) );
  HS65_LS_IVX9 U886 ( .A(phitOut1[28]), .Z(n559) );
  HS65_LS_IVX9 U887 ( .A(phitOut0[28]), .Z(n558) );
  HS65_LS_NAND2X7 U888 ( .A(phitOut2[28]), .B(n572), .Z(n557) );
  HS65_LS_OAI212X5 U889 ( .A(n15), .B(n559), .C(n48), .D(n558), .E(n557), .Z(
        pkt_out[28]) );
  HS65_LS_IVX9 U890 ( .A(phitOut1[29]), .Z(n562) );
  HS65_LS_IVX9 U891 ( .A(phitOut0[29]), .Z(n561) );
  HS65_LS_OAI212X5 U892 ( .A(n22), .B(n562), .C(n48), .D(n561), .E(n560), .Z(
        pkt_out[29]) );
  HS65_LS_IVX9 U893 ( .A(phitOut1[30]), .Z(n565) );
  HS65_LS_IVX9 U894 ( .A(phitOut0[30]), .Z(n564) );
  HS65_LS_NAND2X7 U895 ( .A(phitOut2[30]), .B(n572), .Z(n563) );
  HS65_LS_OAI212X5 U896 ( .A(n22), .B(n565), .C(n48), .D(n564), .E(n563), .Z(
        pkt_out[30]) );
  HS65_LS_IVX9 U897 ( .A(phitOut1[31]), .Z(n568) );
  HS65_LS_IVX9 U898 ( .A(phitOut0[31]), .Z(n567) );
  HS65_LS_NAND2X7 U899 ( .A(phitOut2[31]), .B(n572), .Z(n566) );
  HS65_LS_OAI212X5 U900 ( .A(n15), .B(n568), .C(n47), .D(n567), .E(n566), .Z(
        pkt_out[31]) );
  HS65_LS_IVX9 U901 ( .A(phitOut1[32]), .Z(n571) );
  HS65_LS_IVX9 U902 ( .A(phitOut0[32]), .Z(n570) );
  HS65_LS_NAND2X7 U903 ( .A(phitOut2[32]), .B(n572), .Z(n569) );
  HS65_LS_OAI212X5 U904 ( .A(n15), .B(n571), .C(n47), .D(n570), .E(n569), .Z(
        pkt_out[32]) );
  HS65_LS_IVX9 U905 ( .A(phitOut1[33]), .Z(n576) );
  HS65_LS_IVX9 U906 ( .A(phitOut0[33]), .Z(n574) );
  HS65_LS_OAI212X5 U907 ( .A(n22), .B(n576), .C(n48), .D(n574), .E(n573), .Z(
        pkt_out[33]) );
  HS65_LS_IVX9 U908 ( .A(phitOut1[34]), .Z(n580) );
  HS65_LS_IVX9 U909 ( .A(flit_buf[64]), .Z(n582) );
  HS65_LS_OAI22X6 U910 ( .A(n359), .B(n583), .C(n596), .D(n582), .Z(
        \spm_out[MADDR][0] ) );
  HS65_LS_IVX9 U911 ( .A(flit_buf[65]), .Z(n584) );
  HS65_LS_OAI22X6 U912 ( .A(n359), .B(n585), .C(n596), .D(n584), .Z(
        \spm_out[MADDR][1] ) );
  HS65_LS_IVX9 U913 ( .A(flit_buf[66]), .Z(n586) );
  HS65_LS_OAI22X6 U914 ( .A(n359), .B(n587), .C(n596), .D(n586), .Z(
        \spm_out[MADDR][2] ) );
  HS65_LS_IVX9 U915 ( .A(flit_buf[67]), .Z(n588) );
  HS65_LS_OAI22X6 U916 ( .A(n359), .B(n589), .C(n596), .D(n588), .Z(
        \spm_out[MADDR][3] ) );
  HS65_LS_IVX9 U917 ( .A(flit_buf[68]), .Z(n590) );
  HS65_LS_OAI22X6 U918 ( .A(n359), .B(n591), .C(n596), .D(n590), .Z(
        \spm_out[MADDR][4] ) );
  HS65_LS_IVX9 U919 ( .A(flit_buf[69]), .Z(n592) );
  HS65_LS_OAI22X6 U920 ( .A(n359), .B(n593), .C(n596), .D(n592), .Z(
        \spm_out[MADDR][5] ) );
  HS65_LS_IVX9 U921 ( .A(flit_buf[70]), .Z(n594) );
  HS65_LS_OAI22X6 U922 ( .A(n595), .B(n359), .C(n596), .D(n594), .Z(
        \spm_out[MADDR][6] ) );
  HS65_LS_IVX9 U923 ( .A(n596), .Z(\spm_out[MCMD][0] ) );
  HS65_LS_IVX9 U924 ( .A(n597), .Z(n599) );
  HS65_LS_OAI112X5 U925 ( .A(n872), .B(n599), .C(n871), .D(n598), .Z(
        \proc_out[SCMDACCEPT] ) );
endmodule


module latch_controller_1_30 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_30 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n3, n4, n5, n6;
  assign N0 = preset;

  latch_controller_1_30 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n4), .RN(n3), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n3), .Z(n5) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n6), .B(n5), .Z(N5) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_IVX9 U3 ( .A(lt_enable), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(N0), .Z(n3) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n4), .Z(lt_gated) );
endmodule


module latch_controller_1_29 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_29 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n3, n4, n5, n6;
  assign N0 = preset;

  latch_controller_1_29 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n4), .RN(n3), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n3), .Z(n5) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n6), .B(n5), .Z(N5) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_IVX9 U3 ( .A(lt_enable), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(N0), .Z(n3) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n4), .Z(lt_gated) );
endmodule


module latch_controller_1_28 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_28 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n3, n4, n5, n6;
  assign N0 = preset;

  latch_controller_1_28 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n4), .RN(n3), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n3), .Z(n5) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n6), .B(n5), .Z(N5) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_IVX9 U3 ( .A(lt_enable), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(N0), .Z(n3) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n4), .Z(lt_gated) );
endmodule


module latch_controller_1_27 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_27 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n3, n4, n5, n6;
  assign N0 = preset;

  latch_controller_1_27 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n4), .RN(n3), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n3), .Z(n5) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n6), .B(n5), .Z(N5) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_IVX9 U3 ( .A(lt_enable), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(N0), .Z(n3) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n4), .Z(lt_gated) );
endmodule


module latch_controller_1_26 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_NOR2AX3 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_26 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n3, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_26 controller ( .preset(n3), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLRQX18 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(n3), .Z(n7) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_LDHQX18 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX18 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX18 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX18 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX18 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX18 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX18 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX18 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX18 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX18 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX18 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX18 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX18 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX18 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX18 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX18 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX18 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX18 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX18 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX18 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX18 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX18 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX18 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX18 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX18 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX18 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX18 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX18 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX18 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX18 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX18 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX18 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX18 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX18 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_IVX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_IVX9 U5 ( .A(N0), .Z(n4) );
  HS65_LS_NAND2X7 U9 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_comb_0_0_2 ( data_valid, data_in, preset, data_out, sel );
  input [34:0] data_in;
  output [34:0] data_out;
  output [4:0] sel;
  input data_valid, preset;
  wire   data_in_34, data_in_33, data_in_32, \data_in[31] , \data_in[30] ,
         \data_in[29] , \data_in[28] , \data_in[27] , \data_in[26] ,
         \data_in[25] , \data_in[24] , \data_in[23] , \data_in[22] ,
         \data_in[21] , \data_in[20] , \data_in[19] , \data_in[18] ,
         \data_in[17] , \data_in[16] , N23, N25, N26, N27, N28, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n22,
         n23, n24;
  assign data_out[34] = data_in_34;
  assign data_in_34 = data_in[34];
  assign data_out[33] = data_in_33;
  assign data_in_33 = data_in[33];
  assign data_out[32] = data_in_32;
  assign data_in_32 = data_in[32];
  assign data_out[31] = \data_in[31] ;
  assign \data_in[31]  = data_in[31];
  assign data_out[30] = \data_in[30] ;
  assign \data_in[30]  = data_in[30];
  assign data_out[29] = \data_in[29] ;
  assign \data_in[29]  = data_in[29];
  assign data_out[28] = \data_in[28] ;
  assign \data_in[28]  = data_in[28];
  assign data_out[27] = \data_in[27] ;
  assign \data_in[27]  = data_in[27];
  assign data_out[26] = \data_in[26] ;
  assign \data_in[26]  = data_in[26];
  assign data_out[25] = \data_in[25] ;
  assign \data_in[25]  = data_in[25];
  assign data_out[24] = \data_in[24] ;
  assign \data_in[24]  = data_in[24];
  assign data_out[23] = \data_in[23] ;
  assign \data_in[23]  = data_in[23];
  assign data_out[22] = \data_in[22] ;
  assign \data_in[22]  = data_in[22];
  assign data_out[21] = \data_in[21] ;
  assign \data_in[21]  = data_in[21];
  assign data_out[20] = \data_in[20] ;
  assign \data_in[20]  = data_in[20];
  assign data_out[19] = \data_in[19] ;
  assign \data_in[19]  = data_in[19];
  assign data_out[18] = \data_in[18] ;
  assign \data_in[18]  = data_in[18];
  assign data_out[17] = \data_in[17] ;
  assign \data_in[17]  = data_in[17];
  assign data_out[16] = \data_in[16] ;
  assign \data_in[16]  = data_in[16];
  assign sel[0] = 1'b0;

  HS65_LS_LDHQX9 \sel_reg[4]  ( .G(N23), .D(N28), .Q(sel[4]) );
  HS65_LS_LDHQX9 \sel_reg[3]  ( .G(N23), .D(N27), .Q(sel[3]) );
  HS65_LS_LDHQX9 \sel_reg[2]  ( .G(N23), .D(N26), .Q(sel[2]) );
  HS65_LS_LDHQX9 \sel_reg[1]  ( .G(N23), .D(N25), .Q(sel[1]) );
  HS65_LS_NAND3AX6 U4 ( .A(preset), .B(n23), .C(n2), .Z(n22) );
  HS65_LS_OAI22X6 U5 ( .A(n9), .B(n24), .C(n2), .D(n11), .Z(data_out[7]) );
  HS65_LS_OAI22X6 U6 ( .A(n24), .B(n16), .C(n2), .D(n18), .Z(data_out[0]) );
  HS65_LS_OAI22X6 U7 ( .A(n24), .B(n15), .C(n2), .D(n17), .Z(data_out[1]) );
  HS65_LS_OAI22X6 U8 ( .A(n24), .B(n14), .C(n2), .D(n16), .Z(data_out[2]) );
  HS65_LS_OAI22X6 U9 ( .A(n24), .B(n13), .C(n2), .D(n15), .Z(data_out[3]) );
  HS65_LS_OAI22X6 U10 ( .A(n24), .B(n12), .C(n2), .D(n14), .Z(data_out[4]) );
  HS65_LS_OAI22X6 U11 ( .A(n24), .B(n11), .C(n2), .D(n13), .Z(data_out[5]) );
  HS65_LS_OAI22X6 U12 ( .A(n24), .B(n10), .C(n2), .D(n12), .Z(data_out[6]) );
  HS65_LS_OAI22X6 U13 ( .A(n24), .B(n8), .C(n2), .D(n10), .Z(data_out[8]) );
  HS65_LS_OAI22X6 U14 ( .A(n24), .B(n7), .C(n2), .D(n9), .Z(data_out[9]) );
  HS65_LS_OAI22X6 U15 ( .A(n24), .B(n6), .C(n2), .D(n8), .Z(data_out[10]) );
  HS65_LS_OAI22X6 U16 ( .A(n24), .B(n5), .C(n2), .D(n7), .Z(data_out[11]) );
  HS65_LS_OAI22X6 U17 ( .A(n24), .B(n4), .C(n2), .D(n6), .Z(data_out[12]) );
  HS65_LS_OAI22X6 U18 ( .A(n24), .B(n3), .C(n2), .D(n5), .Z(data_out[13]) );
  HS65_LS_IVX9 U19 ( .A(n24), .Z(n2) );
  HS65_LS_NOR3X4 U20 ( .A(n23), .B(preset), .C(n24), .Z(N28) );
  HS65_LS_NOR3X4 U21 ( .A(n22), .B(n17), .C(n18), .Z(N27) );
  HS65_LS_NAND2X7 U22 ( .A(n17), .B(n18), .Z(n23) );
  HS65_LS_NOR2X6 U23 ( .A(n2), .B(n4), .Z(data_out[14]) );
  HS65_LS_NOR2X6 U24 ( .A(n2), .B(n3), .Z(data_out[15]) );
  HS65_LS_NAND2X14 U25 ( .A(data_in_34), .B(data_in_33), .Z(n24) );
  HS65_LS_IVX9 U26 ( .A(data_in[1]), .Z(n17) );
  HS65_LS_IVX9 U27 ( .A(data_in[0]), .Z(n18) );
  HS65_LS_NOR2X6 U28 ( .A(data_in[1]), .B(n22), .Z(N25) );
  HS65_LS_NOR2X6 U29 ( .A(data_in[0]), .B(n22), .Z(N26) );
  HS65_LS_IVX9 U30 ( .A(data_in[9]), .Z(n9) );
  HS65_LS_IVX9 U31 ( .A(data_in[2]), .Z(n16) );
  HS65_LS_IVX9 U32 ( .A(data_in[3]), .Z(n15) );
  HS65_LS_IVX9 U33 ( .A(data_in[4]), .Z(n14) );
  HS65_LS_IVX9 U34 ( .A(data_in[5]), .Z(n13) );
  HS65_LS_IVX9 U35 ( .A(data_in[6]), .Z(n12) );
  HS65_LS_IVX9 U36 ( .A(data_in[7]), .Z(n11) );
  HS65_LS_IVX9 U37 ( .A(data_in[8]), .Z(n10) );
  HS65_LS_IVX9 U38 ( .A(data_in[10]), .Z(n8) );
  HS65_LS_IVX9 U39 ( .A(data_in[11]), .Z(n7) );
  HS65_LS_IVX9 U40 ( .A(data_in[12]), .Z(n6) );
  HS65_LS_IVX9 U41 ( .A(data_in[13]), .Z(n5) );
  HS65_LS_IVX9 U42 ( .A(data_in[14]), .Z(n4) );
  HS65_LS_IVX9 U43 ( .A(data_in[15]), .Z(n3) );
  HS65_LS_CB4I6X9 U44 ( .A(n2), .B(n1), .C(data_valid), .D(preset), .Z(N23) );
  HS65_LS_IVX9 U45 ( .A(data_in_34), .Z(n1) );
endmodule


module latch_controller_1_10 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_10 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_10 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n7) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_IVX9 U3 ( .A(N0), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_0_0_2 ( preset, .chan_in_f({\chan_in_f[REQ] , \chan_in_f[DATA][34] , 
        \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , 
        \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , 
        \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , 
        \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , 
        \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , 
        \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , 
        \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , 
        \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , 
        \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , 
        \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , 
        \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , 
        \chan_in_f[DATA][0] }), .chan_in_b(\chan_in_b[ACK] ), .chan_out_f({
        \chan_out_f[REQ] , \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , 
        \chan_out_f[DATA][32] , \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , 
        \chan_out_f[DATA][29] , \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , 
        \chan_out_f[DATA][26] , \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , 
        \chan_out_f[DATA][23] , \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , 
        \chan_out_f[DATA][20] , \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , 
        \chan_out_f[DATA][17] , \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , 
        \chan_out_f[DATA][14] , \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , 
        \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , 
        \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , 
        \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , 
        \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), 
    .chan_out_b(\chan_out_b[ACK] ), sel );
  output [4:0] sel;
  input preset, \chan_in_f[REQ] , \chan_in_f[DATA][34] , \chan_in_f[DATA][33] ,
         \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , \chan_in_f[DATA][30] ,
         \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , \chan_in_f[DATA][27] ,
         \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , \chan_in_f[DATA][24] ,
         \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , \chan_in_f[DATA][21] ,
         \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , \chan_in_f[DATA][18] ,
         \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , \chan_in_f[DATA][15] ,
         \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , \chan_in_f[DATA][12] ,
         \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , \chan_in_f[DATA][9] ,
         \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , \chan_in_f[DATA][6] ,
         \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , \chan_in_f[DATA][3] ,
         \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , \chan_in_f[DATA][0] ,
         \chan_out_b[ACK] ;
  output \chan_in_b[ACK] , \chan_out_f[REQ] , \chan_out_f[DATA][34] ,
         \chan_out_f[DATA][33] , \chan_out_f[DATA][32] ,
         \chan_out_f[DATA][31] , \chan_out_f[DATA][30] ,
         \chan_out_f[DATA][29] , \chan_out_f[DATA][28] ,
         \chan_out_f[DATA][27] , \chan_out_f[DATA][26] ,
         \chan_out_f[DATA][25] , \chan_out_f[DATA][24] ,
         \chan_out_f[DATA][23] , \chan_out_f[DATA][22] ,
         \chan_out_f[DATA][21] , \chan_out_f[DATA][20] ,
         \chan_out_f[DATA][19] , \chan_out_f[DATA][18] ,
         \chan_out_f[DATA][17] , \chan_out_f[DATA][16] ,
         \chan_out_f[DATA][15] , \chan_out_f[DATA][14] ,
         \chan_out_f[DATA][13] , \chan_out_f[DATA][12] ,
         \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] ,
         \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] ,
         \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] ,
         \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] ;
  wire   \chan_internal_f[REQ] , \chan_internal_f[DATA][34] ,
         \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] ,
         \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] ,
         \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] ,
         \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] ,
         \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] ,
         \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] ,
         \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] ,
         \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] ,
         \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] ,
         \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] ,
         \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] ,
         \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] ,
         \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] ,
         \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] ,
         \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] ,
         \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] ,
         \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] , req_n, lt_en,
         n1, n2, n3, n4, n5, n6, n7;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign sel[0] = 1'b0;

  hpu_comb_0_0_2 hpu_combinatorial ( .data_valid(lt_en), .data_in({
        \chan_in_f[DATA][34] , \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , 
        \chan_in_f[DATA][31] , \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , 
        \chan_in_f[DATA][28] , \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , 
        \chan_in_f[DATA][25] , \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , 
        \chan_in_f[DATA][22] , \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , 
        \chan_in_f[DATA][19] , \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , 
        \chan_in_f[DATA][16] , \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , 
        \chan_in_f[DATA][13] , \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , 
        \chan_in_f[DATA][10] , \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , 
        \chan_in_f[DATA][7] , \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , 
        \chan_in_f[DATA][4] , \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , 
        \chan_in_f[DATA][1] , \chan_in_f[DATA][0] }), .preset(n7), .data_out({
        \chan_internal_f[DATA][34] , \chan_internal_f[DATA][33] , 
        \chan_internal_f[DATA][32] , \chan_internal_f[DATA][31] , 
        \chan_internal_f[DATA][30] , \chan_internal_f[DATA][29] , 
        \chan_internal_f[DATA][28] , \chan_internal_f[DATA][27] , 
        \chan_internal_f[DATA][26] , \chan_internal_f[DATA][25] , 
        \chan_internal_f[DATA][24] , \chan_internal_f[DATA][23] , 
        \chan_internal_f[DATA][22] , \chan_internal_f[DATA][21] , 
        \chan_internal_f[DATA][20] , \chan_internal_f[DATA][19] , 
        \chan_internal_f[DATA][18] , \chan_internal_f[DATA][17] , 
        \chan_internal_f[DATA][16] , \chan_internal_f[DATA][15] , 
        \chan_internal_f[DATA][14] , \chan_internal_f[DATA][13] , 
        \chan_internal_f[DATA][12] , \chan_internal_f[DATA][11] , 
        \chan_internal_f[DATA][10] , \chan_internal_f[DATA][9] , 
        \chan_internal_f[DATA][8] , \chan_internal_f[DATA][7] , 
        \chan_internal_f[DATA][6] , \chan_internal_f[DATA][5] , 
        \chan_internal_f[DATA][4] , \chan_internal_f[DATA][3] , 
        \chan_internal_f[DATA][2] , \chan_internal_f[DATA][1] , 
        \chan_internal_f[DATA][0] }), .sel({sel[4:1], SYNOPSYS_UNCONNECTED__0}) );
  channel_latch_1_xxxxxxxxx_10 token_latch ( .preset(n7), .left_in({
        \chan_internal_f[REQ] , \chan_internal_f[DATA][34] , 
        \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] , 
        \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] , 
        \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] , 
        \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] , 
        \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] , 
        \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] , 
        \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] , 
        \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] , 
        \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] , 
        \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] , 
        \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] , 
        \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] , 
        \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] , 
        \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] , 
        \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] , 
        \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] , 
        \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] }), .left_out(
        \chan_in_b[ACK] ), .right_out({\chan_out_f[REQ] , 
        \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , \chan_out_f[DATA][32] , 
        \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , \chan_out_f[DATA][29] , 
        \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , \chan_out_f[DATA][26] , 
        \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , \chan_out_f[DATA][23] , 
        \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , \chan_out_f[DATA][20] , 
        \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , \chan_out_f[DATA][17] , 
        \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , \chan_out_f[DATA][14] , 
        \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , \chan_out_f[DATA][11] , 
        \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , \chan_out_f[DATA][8] , 
        \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , \chan_out_f[DATA][5] , 
        \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , \chan_out_f[DATA][2] , 
        \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), .right_in(
        \chan_out_b[ACK] ), .lt_enable(lt_en) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chan_internal_f[REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(\chan_in_f[REQ] ), .Z(req_n) );
  HS65_LS_BFX9 U1 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U2 ( .A(n3), .Z(n2) );
  HS65_LS_BFX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_BFX9 U4 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U6 ( .A(req_n), .Z(n6) );
  HS65_LS_BFX9 U7 ( .A(preset), .Z(n7) );
endmodule


module hpu_comb_0_2_2 ( data_valid, data_in, preset, data_out, sel );
  input [34:0] data_in;
  output [34:0] data_out;
  output [4:0] sel;
  input data_valid, preset;
  wire   data_in_34, data_in_33, data_in_32, \data_in[31] , \data_in[30] ,
         \data_in[29] , \data_in[28] , \data_in[27] , \data_in[26] ,
         \data_in[25] , \data_in[24] , \data_in[23] , \data_in[22] ,
         \data_in[21] , \data_in[20] , \data_in[19] , \data_in[18] ,
         \data_in[17] , \data_in[16] , N26, N27, N28, N30, N31, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n15, n16, n17, n18;
  assign data_out[34] = data_in_34;
  assign data_in_34 = data_in[34];
  assign data_out[33] = data_in_33;
  assign data_in_33 = data_in[33];
  assign data_out[32] = data_in_32;
  assign data_in_32 = data_in[32];
  assign data_out[31] = \data_in[31] ;
  assign \data_in[31]  = data_in[31];
  assign data_out[30] = \data_in[30] ;
  assign \data_in[30]  = data_in[30];
  assign data_out[29] = \data_in[29] ;
  assign \data_in[29]  = data_in[29];
  assign data_out[28] = \data_in[28] ;
  assign \data_in[28]  = data_in[28];
  assign data_out[27] = \data_in[27] ;
  assign \data_in[27]  = data_in[27];
  assign data_out[26] = \data_in[26] ;
  assign \data_in[26]  = data_in[26];
  assign data_out[25] = \data_in[25] ;
  assign \data_in[25]  = data_in[25];
  assign data_out[24] = \data_in[24] ;
  assign \data_in[24]  = data_in[24];
  assign data_out[23] = \data_in[23] ;
  assign \data_in[23]  = data_in[23];
  assign data_out[22] = \data_in[22] ;
  assign \data_in[22]  = data_in[22];
  assign data_out[21] = \data_in[21] ;
  assign \data_in[21]  = data_in[21];
  assign data_out[20] = \data_in[20] ;
  assign \data_in[20]  = data_in[20];
  assign data_out[19] = \data_in[19] ;
  assign \data_in[19]  = data_in[19];
  assign data_out[18] = \data_in[18] ;
  assign \data_in[18]  = data_in[18];
  assign data_out[17] = \data_in[17] ;
  assign \data_in[17]  = data_in[17];
  assign data_out[16] = \data_in[16] ;
  assign \data_in[16]  = data_in[16];
  assign sel[2] = 1'b0;

  HS65_LS_LDHQX9 \sel_reg[4]  ( .G(N26), .D(N31), .Q(sel[4]) );
  HS65_LS_LDHQX9 \sel_reg[3]  ( .G(N26), .D(N30), .Q(sel[3]) );
  HS65_LS_LDHQX9 \sel_reg[1]  ( .G(N26), .D(N28), .Q(sel[1]) );
  HS65_LS_LDHQX9 \sel_reg[0]  ( .G(N26), .D(N27), .Q(sel[0]) );
  HS65_LS_OAI22X6 U4 ( .A(n18), .B(n9), .C(n2), .D(n10), .Z(data_out[0]) );
  HS65_LS_OAI22X6 U5 ( .A(n18), .B(n8), .C(n2), .D(n9), .Z(data_out[2]) );
  HS65_LS_OAI22X6 U6 ( .A(n18), .B(n7), .C(n2), .D(n8), .Z(data_out[4]) );
  HS65_LS_OAI22X6 U7 ( .A(n18), .B(n6), .C(n2), .D(n7), .Z(data_out[6]) );
  HS65_LS_OAI22X6 U8 ( .A(n18), .B(n5), .C(n2), .D(n6), .Z(data_out[8]) );
  HS65_LS_OAI22X6 U9 ( .A(n18), .B(n4), .C(n2), .D(n5), .Z(data_out[10]) );
  HS65_LS_OAI22X6 U10 ( .A(n18), .B(n3), .C(n2), .D(n4), .Z(data_out[12]) );
  HS65_LS_NAND3AX6 U11 ( .A(preset), .B(n17), .C(n2), .Z(n16) );
  HS65_LS_NOR3X4 U12 ( .A(n17), .B(preset), .C(n18), .Z(N31) );
  HS65_LS_IVX9 U13 ( .A(n18), .Z(n2) );
  HS65_LS_NOR3X4 U14 ( .A(n16), .B(n10), .C(n15), .Z(N30) );
  HS65_LS_NOR2AX3 U15 ( .A(n15), .B(n16), .Z(N28) );
  HS65_LS_NOR2X6 U16 ( .A(n2), .B(n3), .Z(data_out[14]) );
  HS65_LS_NAND2X14 U17 ( .A(data_in_34), .B(data_in_33), .Z(n18) );
  HS65_LS_IVX9 U18 ( .A(data_in[0]), .Z(n10) );
  HS65_LS_NAND2X7 U19 ( .A(data_in[1]), .B(n10), .Z(n17) );
  HS65_LS_NOR2X6 U20 ( .A(n10), .B(data_in[1]), .Z(n15) );
  HS65_LS_NOR2X6 U21 ( .A(data_in[0]), .B(n16), .Z(N27) );
  HS65_LS_IVX9 U22 ( .A(data_in[2]), .Z(n9) );
  HS65_LS_IVX9 U23 ( .A(data_in[4]), .Z(n8) );
  HS65_LS_IVX9 U24 ( .A(data_in[6]), .Z(n7) );
  HS65_LS_IVX9 U25 ( .A(data_in[8]), .Z(n6) );
  HS65_LS_IVX9 U26 ( .A(data_in[10]), .Z(n5) );
  HS65_LS_IVX9 U27 ( .A(data_in[12]), .Z(n4) );
  HS65_LS_IVX9 U28 ( .A(data_in[14]), .Z(n3) );
  HS65_LS_AO22X9 U29 ( .A(n2), .B(data_in[3]), .C(n18), .D(data_in[1]), .Z(
        data_out[1]) );
  HS65_LS_AO22X9 U30 ( .A(n2), .B(data_in[5]), .C(n18), .D(data_in[3]), .Z(
        data_out[3]) );
  HS65_LS_AO22X9 U31 ( .A(n2), .B(data_in[7]), .C(n18), .D(data_in[5]), .Z(
        data_out[5]) );
  HS65_LS_AO22X9 U32 ( .A(data_in[9]), .B(n2), .C(n18), .D(data_in[7]), .Z(
        data_out[7]) );
  HS65_LS_AO22X9 U33 ( .A(n2), .B(data_in[11]), .C(n18), .D(data_in[9]), .Z(
        data_out[9]) );
  HS65_LS_AO22X9 U34 ( .A(n2), .B(data_in[13]), .C(n18), .D(data_in[11]), .Z(
        data_out[11]) );
  HS65_LS_AO22X9 U35 ( .A(n2), .B(data_in[15]), .C(n18), .D(data_in[13]), .Z(
        data_out[13]) );
  HS65_LS_AND2X4 U36 ( .A(data_in[15]), .B(n18), .Z(data_out[15]) );
  HS65_LS_CB4I6X9 U37 ( .A(n2), .B(n1), .C(data_valid), .D(preset), .Z(N26) );
  HS65_LS_IVX9 U38 ( .A(data_in_34), .Z(n1) );
endmodule


module latch_controller_1_9 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_9 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_9 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n7) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_IVX9 U3 ( .A(N0), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_0_2_2 ( preset, .chan_in_f({\chan_in_f[REQ] , \chan_in_f[DATA][34] , 
        \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , 
        \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , 
        \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , 
        \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , 
        \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , 
        \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , 
        \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , 
        \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , 
        \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , 
        \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , 
        \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , 
        \chan_in_f[DATA][0] }), .chan_in_b(\chan_in_b[ACK] ), .chan_out_f({
        \chan_out_f[REQ] , \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , 
        \chan_out_f[DATA][32] , \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , 
        \chan_out_f[DATA][29] , \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , 
        \chan_out_f[DATA][26] , \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , 
        \chan_out_f[DATA][23] , \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , 
        \chan_out_f[DATA][20] , \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , 
        \chan_out_f[DATA][17] , \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , 
        \chan_out_f[DATA][14] , \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , 
        \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , 
        \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , 
        \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , 
        \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), 
    .chan_out_b(\chan_out_b[ACK] ), sel );
  output [4:0] sel;
  input preset, \chan_in_f[REQ] , \chan_in_f[DATA][34] , \chan_in_f[DATA][33] ,
         \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , \chan_in_f[DATA][30] ,
         \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , \chan_in_f[DATA][27] ,
         \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , \chan_in_f[DATA][24] ,
         \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , \chan_in_f[DATA][21] ,
         \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , \chan_in_f[DATA][18] ,
         \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , \chan_in_f[DATA][15] ,
         \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , \chan_in_f[DATA][12] ,
         \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , \chan_in_f[DATA][9] ,
         \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , \chan_in_f[DATA][6] ,
         \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , \chan_in_f[DATA][3] ,
         \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , \chan_in_f[DATA][0] ,
         \chan_out_b[ACK] ;
  output \chan_in_b[ACK] , \chan_out_f[REQ] , \chan_out_f[DATA][34] ,
         \chan_out_f[DATA][33] , \chan_out_f[DATA][32] ,
         \chan_out_f[DATA][31] , \chan_out_f[DATA][30] ,
         \chan_out_f[DATA][29] , \chan_out_f[DATA][28] ,
         \chan_out_f[DATA][27] , \chan_out_f[DATA][26] ,
         \chan_out_f[DATA][25] , \chan_out_f[DATA][24] ,
         \chan_out_f[DATA][23] , \chan_out_f[DATA][22] ,
         \chan_out_f[DATA][21] , \chan_out_f[DATA][20] ,
         \chan_out_f[DATA][19] , \chan_out_f[DATA][18] ,
         \chan_out_f[DATA][17] , \chan_out_f[DATA][16] ,
         \chan_out_f[DATA][15] , \chan_out_f[DATA][14] ,
         \chan_out_f[DATA][13] , \chan_out_f[DATA][12] ,
         \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] ,
         \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] ,
         \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] ,
         \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] ;
  wire   \chan_internal_f[REQ] , \chan_internal_f[DATA][34] ,
         \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] ,
         \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] ,
         \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] ,
         \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] ,
         \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] ,
         \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] ,
         \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] ,
         \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] ,
         \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] ,
         \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] ,
         \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] ,
         \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] ,
         \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] ,
         \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] ,
         \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] ,
         \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] ,
         \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] , req_n, lt_en,
         n1, n2, n3, n4, n5, n6, n7;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign sel[2] = 1'b0;

  hpu_comb_0_2_2 hpu_combinatorial ( .data_valid(lt_en), .data_in({
        \chan_in_f[DATA][34] , \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , 
        \chan_in_f[DATA][31] , \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , 
        \chan_in_f[DATA][28] , \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , 
        \chan_in_f[DATA][25] , \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , 
        \chan_in_f[DATA][22] , \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , 
        \chan_in_f[DATA][19] , \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , 
        \chan_in_f[DATA][16] , \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , 
        \chan_in_f[DATA][13] , \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , 
        \chan_in_f[DATA][10] , \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , 
        \chan_in_f[DATA][7] , \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , 
        \chan_in_f[DATA][4] , \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , 
        \chan_in_f[DATA][1] , \chan_in_f[DATA][0] }), .preset(n7), .data_out({
        \chan_internal_f[DATA][34] , \chan_internal_f[DATA][33] , 
        \chan_internal_f[DATA][32] , \chan_internal_f[DATA][31] , 
        \chan_internal_f[DATA][30] , \chan_internal_f[DATA][29] , 
        \chan_internal_f[DATA][28] , \chan_internal_f[DATA][27] , 
        \chan_internal_f[DATA][26] , \chan_internal_f[DATA][25] , 
        \chan_internal_f[DATA][24] , \chan_internal_f[DATA][23] , 
        \chan_internal_f[DATA][22] , \chan_internal_f[DATA][21] , 
        \chan_internal_f[DATA][20] , \chan_internal_f[DATA][19] , 
        \chan_internal_f[DATA][18] , \chan_internal_f[DATA][17] , 
        \chan_internal_f[DATA][16] , \chan_internal_f[DATA][15] , 
        \chan_internal_f[DATA][14] , \chan_internal_f[DATA][13] , 
        \chan_internal_f[DATA][12] , \chan_internal_f[DATA][11] , 
        \chan_internal_f[DATA][10] , \chan_internal_f[DATA][9] , 
        \chan_internal_f[DATA][8] , \chan_internal_f[DATA][7] , 
        \chan_internal_f[DATA][6] , \chan_internal_f[DATA][5] , 
        \chan_internal_f[DATA][4] , \chan_internal_f[DATA][3] , 
        \chan_internal_f[DATA][2] , \chan_internal_f[DATA][1] , 
        \chan_internal_f[DATA][0] }), .sel({sel[4:3], SYNOPSYS_UNCONNECTED__0, 
        sel[1:0]}) );
  channel_latch_1_xxxxxxxxx_9 token_latch ( .preset(n7), .left_in({
        \chan_internal_f[REQ] , \chan_internal_f[DATA][34] , 
        \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] , 
        \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] , 
        \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] , 
        \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] , 
        \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] , 
        \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] , 
        \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] , 
        \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] , 
        \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] , 
        \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] , 
        \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] , 
        \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] , 
        \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] , 
        \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] , 
        \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] , 
        \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] , 
        \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] }), .left_out(
        \chan_in_b[ACK] ), .right_out({\chan_out_f[REQ] , 
        \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , \chan_out_f[DATA][32] , 
        \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , \chan_out_f[DATA][29] , 
        \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , \chan_out_f[DATA][26] , 
        \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , \chan_out_f[DATA][23] , 
        \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , \chan_out_f[DATA][20] , 
        \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , \chan_out_f[DATA][17] , 
        \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , \chan_out_f[DATA][14] , 
        \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , \chan_out_f[DATA][11] , 
        \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , \chan_out_f[DATA][8] , 
        \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , \chan_out_f[DATA][5] , 
        \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , \chan_out_f[DATA][2] , 
        \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), .right_in(
        \chan_out_b[ACK] ), .lt_enable(lt_en) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chan_internal_f[REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(\chan_in_f[REQ] ), .Z(req_n) );
  HS65_LS_BFX9 U1 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U2 ( .A(n3), .Z(n2) );
  HS65_LS_BFX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_BFX9 U4 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U6 ( .A(req_n), .Z(n6) );
  HS65_LS_BFX9 U7 ( .A(preset), .Z(n7) );
endmodule


module hpu_comb_0_1_2 ( data_valid, data_in, preset, data_out, sel );
  input [34:0] data_in;
  output [34:0] data_out;
  output [4:0] sel;
  input data_valid, preset;
  wire   data_in_34, data_in_33, data_in_32, \data_in[31] , \data_in[30] ,
         \data_in[29] , \data_in[28] , \data_in[27] , \data_in[26] ,
         \data_in[25] , \data_in[24] , \data_in[23] , \data_in[22] ,
         \data_in[21] , \data_in[20] , \data_in[19] , \data_in[18] ,
         \data_in[17] , \data_in[16] , N23, N24, N26, N27, N28, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n15, n16, n17, n18;
  assign data_out[34] = data_in_34;
  assign data_in_34 = data_in[34];
  assign data_out[33] = data_in_33;
  assign data_in_33 = data_in[33];
  assign data_out[32] = data_in_32;
  assign data_in_32 = data_in[32];
  assign data_out[31] = \data_in[31] ;
  assign \data_in[31]  = data_in[31];
  assign data_out[30] = \data_in[30] ;
  assign \data_in[30]  = data_in[30];
  assign data_out[29] = \data_in[29] ;
  assign \data_in[29]  = data_in[29];
  assign data_out[28] = \data_in[28] ;
  assign \data_in[28]  = data_in[28];
  assign data_out[27] = \data_in[27] ;
  assign \data_in[27]  = data_in[27];
  assign data_out[26] = \data_in[26] ;
  assign \data_in[26]  = data_in[26];
  assign data_out[25] = \data_in[25] ;
  assign \data_in[25]  = data_in[25];
  assign data_out[24] = \data_in[24] ;
  assign \data_in[24]  = data_in[24];
  assign data_out[23] = \data_in[23] ;
  assign \data_in[23]  = data_in[23];
  assign data_out[22] = \data_in[22] ;
  assign \data_in[22]  = data_in[22];
  assign data_out[21] = \data_in[21] ;
  assign \data_in[21]  = data_in[21];
  assign data_out[20] = \data_in[20] ;
  assign \data_in[20]  = data_in[20];
  assign data_out[19] = \data_in[19] ;
  assign \data_in[19]  = data_in[19];
  assign data_out[18] = \data_in[18] ;
  assign \data_in[18]  = data_in[18];
  assign data_out[17] = \data_in[17] ;
  assign \data_in[17]  = data_in[17];
  assign data_out[16] = \data_in[16] ;
  assign \data_in[16]  = data_in[16];
  assign sel[1] = 1'b0;

  HS65_LS_LDHQX9 \sel_reg[4]  ( .G(N23), .D(N28), .Q(sel[4]) );
  HS65_LS_LDHQX9 \sel_reg[3]  ( .G(N23), .D(N27), .Q(sel[3]) );
  HS65_LS_LDHQX9 \sel_reg[2]  ( .G(N23), .D(N26), .Q(sel[2]) );
  HS65_LS_LDHQX9 \sel_reg[0]  ( .G(N23), .D(N24), .Q(sel[0]) );
  HS65_LS_OAI22X6 U4 ( .A(n6), .B(n18), .C(n2), .D(n7), .Z(data_out[7]) );
  HS65_LS_OAI22X6 U5 ( .A(n18), .B(n9), .C(n2), .D(n10), .Z(data_out[1]) );
  HS65_LS_OAI22X6 U6 ( .A(n18), .B(n8), .C(n2), .D(n9), .Z(data_out[3]) );
  HS65_LS_OAI22X6 U7 ( .A(n18), .B(n7), .C(n2), .D(n8), .Z(data_out[5]) );
  HS65_LS_OAI22X6 U8 ( .A(n18), .B(n5), .C(n2), .D(n6), .Z(data_out[9]) );
  HS65_LS_OAI22X6 U9 ( .A(n18), .B(n4), .C(n2), .D(n5), .Z(data_out[11]) );
  HS65_LS_OAI22X6 U10 ( .A(n18), .B(n3), .C(n2), .D(n4), .Z(data_out[13]) );
  HS65_LS_NAND3AX6 U11 ( .A(preset), .B(n17), .C(n2), .Z(n16) );
  HS65_LS_NOR3X4 U12 ( .A(n17), .B(preset), .C(n18), .Z(N28) );
  HS65_LS_IVX9 U13 ( .A(n18), .Z(n2) );
  HS65_LS_NOR3X4 U14 ( .A(n16), .B(n10), .C(n15), .Z(N27) );
  HS65_LS_NOR2AX3 U15 ( .A(n15), .B(n16), .Z(N26) );
  HS65_LS_NOR2X6 U16 ( .A(n2), .B(n3), .Z(data_out[15]) );
  HS65_LS_NAND2X14 U17 ( .A(data_in_34), .B(data_in_33), .Z(n18) );
  HS65_LS_IVX9 U18 ( .A(data_in[1]), .Z(n10) );
  HS65_LS_NAND2X7 U19 ( .A(data_in[0]), .B(n10), .Z(n17) );
  HS65_LS_NOR2X6 U20 ( .A(n10), .B(data_in[0]), .Z(n15) );
  HS65_LS_NOR2X6 U21 ( .A(data_in[1]), .B(n16), .Z(N24) );
  HS65_LS_IVX9 U22 ( .A(data_in[9]), .Z(n6) );
  HS65_LS_IVX9 U23 ( .A(data_in[3]), .Z(n9) );
  HS65_LS_IVX9 U24 ( .A(data_in[5]), .Z(n8) );
  HS65_LS_IVX9 U25 ( .A(data_in[7]), .Z(n7) );
  HS65_LS_IVX9 U26 ( .A(data_in[11]), .Z(n5) );
  HS65_LS_IVX9 U27 ( .A(data_in[13]), .Z(n4) );
  HS65_LS_IVX9 U28 ( .A(data_in[15]), .Z(n3) );
  HS65_LS_AO22X9 U29 ( .A(n2), .B(data_in[2]), .C(n18), .D(data_in[0]), .Z(
        data_out[0]) );
  HS65_LS_AO22X9 U30 ( .A(n2), .B(data_in[4]), .C(n18), .D(data_in[2]), .Z(
        data_out[2]) );
  HS65_LS_AO22X9 U31 ( .A(n2), .B(data_in[6]), .C(n18), .D(data_in[4]), .Z(
        data_out[4]) );
  HS65_LS_AO22X9 U32 ( .A(n2), .B(data_in[8]), .C(n18), .D(data_in[6]), .Z(
        data_out[6]) );
  HS65_LS_AO22X9 U33 ( .A(n2), .B(data_in[10]), .C(n18), .D(data_in[8]), .Z(
        data_out[8]) );
  HS65_LS_AO22X9 U34 ( .A(n2), .B(data_in[12]), .C(n18), .D(data_in[10]), .Z(
        data_out[10]) );
  HS65_LS_AO22X9 U35 ( .A(n2), .B(data_in[14]), .C(n18), .D(data_in[12]), .Z(
        data_out[12]) );
  HS65_LS_AND2X4 U36 ( .A(data_in[14]), .B(n18), .Z(data_out[14]) );
  HS65_LS_CB4I6X9 U37 ( .A(n2), .B(n1), .C(data_valid), .D(preset), .Z(N23) );
  HS65_LS_IVX9 U38 ( .A(data_in_34), .Z(n1) );
endmodule


module latch_controller_1_8 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_8 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_8 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n7) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_IVX9 U3 ( .A(N0), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_0_1_2 ( preset, .chan_in_f({\chan_in_f[REQ] , \chan_in_f[DATA][34] , 
        \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , 
        \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , 
        \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , 
        \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , 
        \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , 
        \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , 
        \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , 
        \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , 
        \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , 
        \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , 
        \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , 
        \chan_in_f[DATA][0] }), .chan_in_b(\chan_in_b[ACK] ), .chan_out_f({
        \chan_out_f[REQ] , \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , 
        \chan_out_f[DATA][32] , \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , 
        \chan_out_f[DATA][29] , \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , 
        \chan_out_f[DATA][26] , \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , 
        \chan_out_f[DATA][23] , \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , 
        \chan_out_f[DATA][20] , \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , 
        \chan_out_f[DATA][17] , \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , 
        \chan_out_f[DATA][14] , \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , 
        \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , 
        \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , 
        \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , 
        \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), 
    .chan_out_b(\chan_out_b[ACK] ), sel );
  output [4:0] sel;
  input preset, \chan_in_f[REQ] , \chan_in_f[DATA][34] , \chan_in_f[DATA][33] ,
         \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , \chan_in_f[DATA][30] ,
         \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , \chan_in_f[DATA][27] ,
         \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , \chan_in_f[DATA][24] ,
         \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , \chan_in_f[DATA][21] ,
         \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , \chan_in_f[DATA][18] ,
         \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , \chan_in_f[DATA][15] ,
         \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , \chan_in_f[DATA][12] ,
         \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , \chan_in_f[DATA][9] ,
         \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , \chan_in_f[DATA][6] ,
         \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , \chan_in_f[DATA][3] ,
         \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , \chan_in_f[DATA][0] ,
         \chan_out_b[ACK] ;
  output \chan_in_b[ACK] , \chan_out_f[REQ] , \chan_out_f[DATA][34] ,
         \chan_out_f[DATA][33] , \chan_out_f[DATA][32] ,
         \chan_out_f[DATA][31] , \chan_out_f[DATA][30] ,
         \chan_out_f[DATA][29] , \chan_out_f[DATA][28] ,
         \chan_out_f[DATA][27] , \chan_out_f[DATA][26] ,
         \chan_out_f[DATA][25] , \chan_out_f[DATA][24] ,
         \chan_out_f[DATA][23] , \chan_out_f[DATA][22] ,
         \chan_out_f[DATA][21] , \chan_out_f[DATA][20] ,
         \chan_out_f[DATA][19] , \chan_out_f[DATA][18] ,
         \chan_out_f[DATA][17] , \chan_out_f[DATA][16] ,
         \chan_out_f[DATA][15] , \chan_out_f[DATA][14] ,
         \chan_out_f[DATA][13] , \chan_out_f[DATA][12] ,
         \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] ,
         \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] ,
         \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] ,
         \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] ;
  wire   \chan_internal_f[REQ] , \chan_internal_f[DATA][34] ,
         \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] ,
         \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] ,
         \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] ,
         \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] ,
         \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] ,
         \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] ,
         \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] ,
         \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] ,
         \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] ,
         \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] ,
         \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] ,
         \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] ,
         \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] ,
         \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] ,
         \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] ,
         \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] ,
         \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] , req_n, lt_en,
         n1, n2, n3, n4, n5, n6, n7;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign sel[1] = 1'b0;

  hpu_comb_0_1_2 hpu_combinatorial ( .data_valid(lt_en), .data_in({
        \chan_in_f[DATA][34] , \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , 
        \chan_in_f[DATA][31] , \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , 
        \chan_in_f[DATA][28] , \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , 
        \chan_in_f[DATA][25] , \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , 
        \chan_in_f[DATA][22] , \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , 
        \chan_in_f[DATA][19] , \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , 
        \chan_in_f[DATA][16] , \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , 
        \chan_in_f[DATA][13] , \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , 
        \chan_in_f[DATA][10] , \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , 
        \chan_in_f[DATA][7] , \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , 
        \chan_in_f[DATA][4] , \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , 
        \chan_in_f[DATA][1] , \chan_in_f[DATA][0] }), .preset(n7), .data_out({
        \chan_internal_f[DATA][34] , \chan_internal_f[DATA][33] , 
        \chan_internal_f[DATA][32] , \chan_internal_f[DATA][31] , 
        \chan_internal_f[DATA][30] , \chan_internal_f[DATA][29] , 
        \chan_internal_f[DATA][28] , \chan_internal_f[DATA][27] , 
        \chan_internal_f[DATA][26] , \chan_internal_f[DATA][25] , 
        \chan_internal_f[DATA][24] , \chan_internal_f[DATA][23] , 
        \chan_internal_f[DATA][22] , \chan_internal_f[DATA][21] , 
        \chan_internal_f[DATA][20] , \chan_internal_f[DATA][19] , 
        \chan_internal_f[DATA][18] , \chan_internal_f[DATA][17] , 
        \chan_internal_f[DATA][16] , \chan_internal_f[DATA][15] , 
        \chan_internal_f[DATA][14] , \chan_internal_f[DATA][13] , 
        \chan_internal_f[DATA][12] , \chan_internal_f[DATA][11] , 
        \chan_internal_f[DATA][10] , \chan_internal_f[DATA][9] , 
        \chan_internal_f[DATA][8] , \chan_internal_f[DATA][7] , 
        \chan_internal_f[DATA][6] , \chan_internal_f[DATA][5] , 
        \chan_internal_f[DATA][4] , \chan_internal_f[DATA][3] , 
        \chan_internal_f[DATA][2] , \chan_internal_f[DATA][1] , 
        \chan_internal_f[DATA][0] }), .sel({sel[4:2], SYNOPSYS_UNCONNECTED__0, 
        sel[0]}) );
  channel_latch_1_xxxxxxxxx_8 token_latch ( .preset(n7), .left_in({
        \chan_internal_f[REQ] , \chan_internal_f[DATA][34] , 
        \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] , 
        \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] , 
        \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] , 
        \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] , 
        \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] , 
        \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] , 
        \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] , 
        \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] , 
        \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] , 
        \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] , 
        \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] , 
        \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] , 
        \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] , 
        \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] , 
        \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] , 
        \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] , 
        \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] }), .left_out(
        \chan_in_b[ACK] ), .right_out({\chan_out_f[REQ] , 
        \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , \chan_out_f[DATA][32] , 
        \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , \chan_out_f[DATA][29] , 
        \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , \chan_out_f[DATA][26] , 
        \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , \chan_out_f[DATA][23] , 
        \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , \chan_out_f[DATA][20] , 
        \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , \chan_out_f[DATA][17] , 
        \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , \chan_out_f[DATA][14] , 
        \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , \chan_out_f[DATA][11] , 
        \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , \chan_out_f[DATA][8] , 
        \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , \chan_out_f[DATA][5] , 
        \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , \chan_out_f[DATA][2] , 
        \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), .right_in(
        \chan_out_b[ACK] ), .lt_enable(lt_en) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chan_internal_f[REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(\chan_in_f[REQ] ), .Z(req_n) );
  HS65_LS_BFX9 U1 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U2 ( .A(n3), .Z(n2) );
  HS65_LS_BFX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_BFX9 U4 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U6 ( .A(req_n), .Z(n6) );
  HS65_LS_BFX9 U7 ( .A(preset), .Z(n7) );
endmodule


module hpu_comb_0_3_2 ( data_valid, data_in, preset, data_out, sel );
  input [34:0] data_in;
  output [34:0] data_out;
  output [4:0] sel;
  input data_valid, preset;
  wire   data_in_34, data_in_33, data_in_32, \data_in[31] , \data_in[30] ,
         \data_in[29] , \data_in[28] , \data_in[27] , \data_in[26] ,
         \data_in[25] , \data_in[24] , \data_in[23] , \data_in[22] ,
         \data_in[21] , \data_in[20] , \data_in[19] , \data_in[18] ,
         \data_in[17] , \data_in[16] , N25, N26, N27, N28, N30, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n15, n16, n17, n18;
  assign data_out[34] = data_in_34;
  assign data_in_34 = data_in[34];
  assign data_out[33] = data_in_33;
  assign data_in_33 = data_in[33];
  assign data_out[32] = data_in_32;
  assign data_in_32 = data_in[32];
  assign data_out[31] = \data_in[31] ;
  assign \data_in[31]  = data_in[31];
  assign data_out[30] = \data_in[30] ;
  assign \data_in[30]  = data_in[30];
  assign data_out[29] = \data_in[29] ;
  assign \data_in[29]  = data_in[29];
  assign data_out[28] = \data_in[28] ;
  assign \data_in[28]  = data_in[28];
  assign data_out[27] = \data_in[27] ;
  assign \data_in[27]  = data_in[27];
  assign data_out[26] = \data_in[26] ;
  assign \data_in[26]  = data_in[26];
  assign data_out[25] = \data_in[25] ;
  assign \data_in[25]  = data_in[25];
  assign data_out[24] = \data_in[24] ;
  assign \data_in[24]  = data_in[24];
  assign data_out[23] = \data_in[23] ;
  assign \data_in[23]  = data_in[23];
  assign data_out[22] = \data_in[22] ;
  assign \data_in[22]  = data_in[22];
  assign data_out[21] = \data_in[21] ;
  assign \data_in[21]  = data_in[21];
  assign data_out[20] = \data_in[20] ;
  assign \data_in[20]  = data_in[20];
  assign data_out[19] = \data_in[19] ;
  assign \data_in[19]  = data_in[19];
  assign data_out[18] = \data_in[18] ;
  assign \data_in[18]  = data_in[18];
  assign data_out[17] = \data_in[17] ;
  assign \data_in[17]  = data_in[17];
  assign data_out[16] = \data_in[16] ;
  assign \data_in[16]  = data_in[16];
  assign sel[3] = 1'b0;

  HS65_LS_LDHQX9 \sel_reg[4]  ( .G(N25), .D(N30), .Q(sel[4]) );
  HS65_LS_LDHQX9 \sel_reg[2]  ( .G(N25), .D(N28), .Q(sel[2]) );
  HS65_LS_LDHQX9 \sel_reg[1]  ( .G(N25), .D(N27), .Q(sel[1]) );
  HS65_LS_LDHQX9 \sel_reg[0]  ( .G(N25), .D(N26), .Q(sel[0]) );
  HS65_LS_OAI22X6 U4 ( .A(n18), .B(n9), .C(n2), .D(n10), .Z(data_out[0]) );
  HS65_LS_OAI22X6 U5 ( .A(n18), .B(n8), .C(n2), .D(n9), .Z(data_out[2]) );
  HS65_LS_OAI22X6 U6 ( .A(n18), .B(n7), .C(n2), .D(n8), .Z(data_out[4]) );
  HS65_LS_OAI22X6 U7 ( .A(n18), .B(n6), .C(n2), .D(n7), .Z(data_out[6]) );
  HS65_LS_OAI22X6 U8 ( .A(n18), .B(n5), .C(n2), .D(n6), .Z(data_out[8]) );
  HS65_LS_OAI22X6 U9 ( .A(n18), .B(n4), .C(n2), .D(n5), .Z(data_out[10]) );
  HS65_LS_OAI22X6 U10 ( .A(n18), .B(n3), .C(n2), .D(n4), .Z(data_out[12]) );
  HS65_LS_NAND3AX6 U11 ( .A(preset), .B(n17), .C(n2), .Z(n16) );
  HS65_LS_NOR3X4 U12 ( .A(n17), .B(preset), .C(n18), .Z(N30) );
  HS65_LS_IVX9 U13 ( .A(n18), .Z(n2) );
  HS65_LS_NOR2X6 U14 ( .A(n10), .B(n16), .Z(N27) );
  HS65_LS_NOR2AX3 U15 ( .A(n15), .B(n16), .Z(N26) );
  HS65_LS_NOR2X6 U16 ( .A(n2), .B(n3), .Z(data_out[14]) );
  HS65_LS_NAND2X14 U17 ( .A(data_in_34), .B(data_in_33), .Z(n18) );
  HS65_LS_NOR3X4 U18 ( .A(n16), .B(data_in[0]), .C(n15), .Z(N28) );
  HS65_LS_NAND2X7 U19 ( .A(data_in[0]), .B(data_in[1]), .Z(n17) );
  HS65_LS_NOR2X6 U20 ( .A(data_in[1]), .B(data_in[0]), .Z(n15) );
  HS65_LS_IVX9 U21 ( .A(data_in[0]), .Z(n10) );
  HS65_LS_IVX9 U22 ( .A(data_in[2]), .Z(n9) );
  HS65_LS_IVX9 U23 ( .A(data_in[4]), .Z(n8) );
  HS65_LS_IVX9 U24 ( .A(data_in[6]), .Z(n7) );
  HS65_LS_IVX9 U25 ( .A(data_in[8]), .Z(n6) );
  HS65_LS_IVX9 U26 ( .A(data_in[10]), .Z(n5) );
  HS65_LS_IVX9 U27 ( .A(data_in[12]), .Z(n4) );
  HS65_LS_IVX9 U28 ( .A(data_in[14]), .Z(n3) );
  HS65_LS_AO22X9 U29 ( .A(n2), .B(data_in[3]), .C(n18), .D(data_in[1]), .Z(
        data_out[1]) );
  HS65_LS_AO22X9 U30 ( .A(n2), .B(data_in[5]), .C(n18), .D(data_in[3]), .Z(
        data_out[3]) );
  HS65_LS_AO22X9 U31 ( .A(n2), .B(data_in[7]), .C(n18), .D(data_in[5]), .Z(
        data_out[5]) );
  HS65_LS_AO22X9 U32 ( .A(data_in[9]), .B(n2), .C(n18), .D(data_in[7]), .Z(
        data_out[7]) );
  HS65_LS_AO22X9 U33 ( .A(n2), .B(data_in[11]), .C(n18), .D(data_in[9]), .Z(
        data_out[9]) );
  HS65_LS_AO22X9 U34 ( .A(n2), .B(data_in[13]), .C(n18), .D(data_in[11]), .Z(
        data_out[11]) );
  HS65_LS_AO22X9 U35 ( .A(n2), .B(data_in[15]), .C(n18), .D(data_in[13]), .Z(
        data_out[13]) );
  HS65_LS_AND2X4 U36 ( .A(data_in[15]), .B(n18), .Z(data_out[15]) );
  HS65_LS_CB4I6X9 U37 ( .A(n2), .B(n1), .C(data_valid), .D(preset), .Z(N25) );
  HS65_LS_IVX9 U38 ( .A(data_in_34), .Z(n1) );
endmodule


module latch_controller_1_7 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_7 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_7 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n7) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_IVX9 U3 ( .A(N0), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_0_3_2 ( preset, .chan_in_f({\chan_in_f[REQ] , \chan_in_f[DATA][34] , 
        \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , 
        \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , 
        \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , 
        \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , 
        \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , 
        \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , 
        \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , 
        \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , 
        \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , 
        \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , 
        \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , 
        \chan_in_f[DATA][0] }), .chan_in_b(\chan_in_b[ACK] ), .chan_out_f({
        \chan_out_f[REQ] , \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , 
        \chan_out_f[DATA][32] , \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , 
        \chan_out_f[DATA][29] , \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , 
        \chan_out_f[DATA][26] , \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , 
        \chan_out_f[DATA][23] , \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , 
        \chan_out_f[DATA][20] , \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , 
        \chan_out_f[DATA][17] , \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , 
        \chan_out_f[DATA][14] , \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , 
        \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , 
        \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , 
        \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , 
        \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), 
    .chan_out_b(\chan_out_b[ACK] ), sel );
  output [4:0] sel;
  input preset, \chan_in_f[REQ] , \chan_in_f[DATA][34] , \chan_in_f[DATA][33] ,
         \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , \chan_in_f[DATA][30] ,
         \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , \chan_in_f[DATA][27] ,
         \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , \chan_in_f[DATA][24] ,
         \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , \chan_in_f[DATA][21] ,
         \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , \chan_in_f[DATA][18] ,
         \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , \chan_in_f[DATA][15] ,
         \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , \chan_in_f[DATA][12] ,
         \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , \chan_in_f[DATA][9] ,
         \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , \chan_in_f[DATA][6] ,
         \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , \chan_in_f[DATA][3] ,
         \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , \chan_in_f[DATA][0] ,
         \chan_out_b[ACK] ;
  output \chan_in_b[ACK] , \chan_out_f[REQ] , \chan_out_f[DATA][34] ,
         \chan_out_f[DATA][33] , \chan_out_f[DATA][32] ,
         \chan_out_f[DATA][31] , \chan_out_f[DATA][30] ,
         \chan_out_f[DATA][29] , \chan_out_f[DATA][28] ,
         \chan_out_f[DATA][27] , \chan_out_f[DATA][26] ,
         \chan_out_f[DATA][25] , \chan_out_f[DATA][24] ,
         \chan_out_f[DATA][23] , \chan_out_f[DATA][22] ,
         \chan_out_f[DATA][21] , \chan_out_f[DATA][20] ,
         \chan_out_f[DATA][19] , \chan_out_f[DATA][18] ,
         \chan_out_f[DATA][17] , \chan_out_f[DATA][16] ,
         \chan_out_f[DATA][15] , \chan_out_f[DATA][14] ,
         \chan_out_f[DATA][13] , \chan_out_f[DATA][12] ,
         \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] ,
         \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] ,
         \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] ,
         \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] ;
  wire   \chan_internal_f[REQ] , \chan_internal_f[DATA][34] ,
         \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] ,
         \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] ,
         \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] ,
         \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] ,
         \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] ,
         \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] ,
         \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] ,
         \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] ,
         \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] ,
         \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] ,
         \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] ,
         \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] ,
         \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] ,
         \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] ,
         \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] ,
         \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] ,
         \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] , req_n, lt_en,
         n1, n2, n3, n4, n5, n6, n7;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign sel[3] = 1'b0;

  hpu_comb_0_3_2 hpu_combinatorial ( .data_valid(lt_en), .data_in({
        \chan_in_f[DATA][34] , \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , 
        \chan_in_f[DATA][31] , \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , 
        \chan_in_f[DATA][28] , \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , 
        \chan_in_f[DATA][25] , \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , 
        \chan_in_f[DATA][22] , \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , 
        \chan_in_f[DATA][19] , \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , 
        \chan_in_f[DATA][16] , \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , 
        \chan_in_f[DATA][13] , \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , 
        \chan_in_f[DATA][10] , \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , 
        \chan_in_f[DATA][7] , \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , 
        \chan_in_f[DATA][4] , \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , 
        \chan_in_f[DATA][1] , \chan_in_f[DATA][0] }), .preset(n7), .data_out({
        \chan_internal_f[DATA][34] , \chan_internal_f[DATA][33] , 
        \chan_internal_f[DATA][32] , \chan_internal_f[DATA][31] , 
        \chan_internal_f[DATA][30] , \chan_internal_f[DATA][29] , 
        \chan_internal_f[DATA][28] , \chan_internal_f[DATA][27] , 
        \chan_internal_f[DATA][26] , \chan_internal_f[DATA][25] , 
        \chan_internal_f[DATA][24] , \chan_internal_f[DATA][23] , 
        \chan_internal_f[DATA][22] , \chan_internal_f[DATA][21] , 
        \chan_internal_f[DATA][20] , \chan_internal_f[DATA][19] , 
        \chan_internal_f[DATA][18] , \chan_internal_f[DATA][17] , 
        \chan_internal_f[DATA][16] , \chan_internal_f[DATA][15] , 
        \chan_internal_f[DATA][14] , \chan_internal_f[DATA][13] , 
        \chan_internal_f[DATA][12] , \chan_internal_f[DATA][11] , 
        \chan_internal_f[DATA][10] , \chan_internal_f[DATA][9] , 
        \chan_internal_f[DATA][8] , \chan_internal_f[DATA][7] , 
        \chan_internal_f[DATA][6] , \chan_internal_f[DATA][5] , 
        \chan_internal_f[DATA][4] , \chan_internal_f[DATA][3] , 
        \chan_internal_f[DATA][2] , \chan_internal_f[DATA][1] , 
        \chan_internal_f[DATA][0] }), .sel({sel[4], SYNOPSYS_UNCONNECTED__0, 
        sel[2:0]}) );
  channel_latch_1_xxxxxxxxx_7 token_latch ( .preset(n7), .left_in({
        \chan_internal_f[REQ] , \chan_internal_f[DATA][34] , 
        \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] , 
        \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] , 
        \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] , 
        \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] , 
        \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] , 
        \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] , 
        \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] , 
        \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] , 
        \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] , 
        \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] , 
        \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] , 
        \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] , 
        \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] , 
        \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] , 
        \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] , 
        \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] , 
        \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] }), .left_out(
        \chan_in_b[ACK] ), .right_out({\chan_out_f[REQ] , 
        \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , \chan_out_f[DATA][32] , 
        \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , \chan_out_f[DATA][29] , 
        \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , \chan_out_f[DATA][26] , 
        \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , \chan_out_f[DATA][23] , 
        \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , \chan_out_f[DATA][20] , 
        \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , \chan_out_f[DATA][17] , 
        \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , \chan_out_f[DATA][14] , 
        \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , \chan_out_f[DATA][11] , 
        \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , \chan_out_f[DATA][8] , 
        \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , \chan_out_f[DATA][5] , 
        \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , \chan_out_f[DATA][2] , 
        \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), .right_in(
        \chan_out_b[ACK] ), .lt_enable(lt_en) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chan_internal_f[REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(\chan_in_f[REQ] ), .Z(req_n) );
  HS65_LS_BFX9 U1 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U2 ( .A(n3), .Z(n2) );
  HS65_LS_BFX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_BFX9 U4 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U6 ( .A(req_n), .Z(n6) );
  HS65_LS_BFX9 U7 ( .A(preset), .Z(n7) );
endmodule


module hpu_comb_1_x_2 ( data_valid, data_in, preset, data_out, sel );
  input [34:0] data_in;
  output [34:0] data_out;
  output [4:0] sel;
  input data_valid, preset;
  wire   data_in_34, data_in_33, data_in_32, \data_in[31] , \data_in[30] ,
         \data_in[29] , \data_in[28] , \data_in[27] , \data_in[26] ,
         \data_in[25] , \data_in[24] , \data_in[23] , \data_in[22] ,
         \data_in[21] , \data_in[20] , \data_in[19] , \data_in[18] ,
         \data_in[17] , \data_in[16] , N19, N20, N21, N22, N23, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n22,
         n23, n24;
  assign data_out[34] = data_in_34;
  assign data_in_34 = data_in[34];
  assign data_out[33] = data_in_33;
  assign data_in_33 = data_in[33];
  assign data_out[32] = data_in_32;
  assign data_in_32 = data_in[32];
  assign data_out[31] = \data_in[31] ;
  assign \data_in[31]  = data_in[31];
  assign data_out[30] = \data_in[30] ;
  assign \data_in[30]  = data_in[30];
  assign data_out[29] = \data_in[29] ;
  assign \data_in[29]  = data_in[29];
  assign data_out[28] = \data_in[28] ;
  assign \data_in[28]  = data_in[28];
  assign data_out[27] = \data_in[27] ;
  assign \data_in[27]  = data_in[27];
  assign data_out[26] = \data_in[26] ;
  assign \data_in[26]  = data_in[26];
  assign data_out[25] = \data_in[25] ;
  assign \data_in[25]  = data_in[25];
  assign data_out[24] = \data_in[24] ;
  assign \data_in[24]  = data_in[24];
  assign data_out[23] = \data_in[23] ;
  assign \data_in[23]  = data_in[23];
  assign data_out[22] = \data_in[22] ;
  assign \data_in[22]  = data_in[22];
  assign data_out[21] = \data_in[21] ;
  assign \data_in[21]  = data_in[21];
  assign data_out[20] = \data_in[20] ;
  assign \data_in[20]  = data_in[20];
  assign data_out[19] = \data_in[19] ;
  assign \data_in[19]  = data_in[19];
  assign data_out[18] = \data_in[18] ;
  assign \data_in[18]  = data_in[18];
  assign data_out[17] = \data_in[17] ;
  assign \data_in[17]  = data_in[17];
  assign data_out[16] = \data_in[16] ;
  assign \data_in[16]  = data_in[16];
  assign sel[4] = 1'b0;

  HS65_LS_LDHQX9 \sel_reg[0]  ( .G(N19), .D(N20), .Q(sel[0]) );
  HS65_LS_LDHQX9 \sel_reg[3]  ( .G(N19), .D(N23), .Q(sel[3]) );
  HS65_LS_LDHQX9 \sel_reg[2]  ( .G(N19), .D(N22), .Q(sel[2]) );
  HS65_LS_LDHQX9 \sel_reg[1]  ( .G(N19), .D(N21), .Q(sel[1]) );
  HS65_LS_NAND2X21 U4 ( .A(data_in_34), .B(data_in_33), .Z(n24) );
  HS65_LS_NAND3AX6 U5 ( .A(preset), .B(n22), .C(n2), .Z(n23) );
  HS65_LS_OAI22X6 U6 ( .A(n9), .B(n24), .C(n2), .D(n11), .Z(data_out[7]) );
  HS65_LS_OAI22X6 U7 ( .A(n24), .B(n16), .C(n2), .D(n18), .Z(data_out[0]) );
  HS65_LS_OAI22X6 U8 ( .A(n24), .B(n15), .C(n2), .D(n17), .Z(data_out[1]) );
  HS65_LS_OAI22X6 U9 ( .A(n24), .B(n14), .C(n2), .D(n16), .Z(data_out[2]) );
  HS65_LS_OAI22X6 U10 ( .A(n24), .B(n13), .C(n2), .D(n15), .Z(data_out[3]) );
  HS65_LS_OAI22X6 U11 ( .A(n24), .B(n12), .C(n2), .D(n14), .Z(data_out[4]) );
  HS65_LS_OAI22X6 U12 ( .A(n24), .B(n11), .C(n2), .D(n13), .Z(data_out[5]) );
  HS65_LS_OAI22X6 U13 ( .A(n24), .B(n10), .C(n2), .D(n12), .Z(data_out[6]) );
  HS65_LS_OAI22X6 U14 ( .A(n24), .B(n8), .C(n2), .D(n10), .Z(data_out[8]) );
  HS65_LS_OAI22X6 U15 ( .A(n24), .B(n7), .C(n2), .D(n9), .Z(data_out[9]) );
  HS65_LS_OAI22X6 U16 ( .A(n24), .B(n6), .C(n2), .D(n8), .Z(data_out[10]) );
  HS65_LS_OAI22X6 U17 ( .A(n24), .B(n5), .C(n2), .D(n7), .Z(data_out[11]) );
  HS65_LS_OAI22X6 U18 ( .A(n24), .B(n4), .C(n2), .D(n6), .Z(data_out[12]) );
  HS65_LS_OAI22X6 U19 ( .A(n24), .B(n3), .C(n2), .D(n5), .Z(data_out[13]) );
  HS65_LS_IVX9 U20 ( .A(n24), .Z(n2) );
  HS65_LS_NOR3X4 U21 ( .A(n22), .B(preset), .C(n24), .Z(N20) );
  HS65_LS_NOR3X4 U22 ( .A(n23), .B(n17), .C(n18), .Z(N23) );
  HS65_LS_NAND2X7 U23 ( .A(n17), .B(n18), .Z(n22) );
  HS65_LS_NOR2X6 U24 ( .A(n2), .B(n4), .Z(data_out[14]) );
  HS65_LS_NOR2X6 U25 ( .A(n2), .B(n3), .Z(data_out[15]) );
  HS65_LS_IVX9 U26 ( .A(data_in[1]), .Z(n17) );
  HS65_LS_IVX9 U27 ( .A(data_in[0]), .Z(n18) );
  HS65_LS_NOR2X6 U28 ( .A(data_in[1]), .B(n23), .Z(N21) );
  HS65_LS_NOR2X6 U29 ( .A(data_in[0]), .B(n23), .Z(N22) );
  HS65_LS_IVX9 U30 ( .A(data_in[9]), .Z(n9) );
  HS65_LS_IVX9 U31 ( .A(data_in[2]), .Z(n16) );
  HS65_LS_IVX9 U32 ( .A(data_in[4]), .Z(n14) );
  HS65_LS_IVX9 U33 ( .A(data_in[5]), .Z(n13) );
  HS65_LS_IVX9 U34 ( .A(data_in[6]), .Z(n12) );
  HS65_LS_IVX9 U35 ( .A(data_in[8]), .Z(n10) );
  HS65_LS_IVX9 U36 ( .A(data_in[10]), .Z(n8) );
  HS65_LS_IVX9 U37 ( .A(data_in[12]), .Z(n6) );
  HS65_LS_IVX9 U38 ( .A(data_in[13]), .Z(n5) );
  HS65_LS_IVX9 U39 ( .A(data_in[14]), .Z(n4) );
  HS65_LS_IVX9 U40 ( .A(data_in[15]), .Z(n3) );
  HS65_LS_IVX9 U41 ( .A(data_in[3]), .Z(n15) );
  HS65_LS_IVX9 U42 ( .A(data_in[7]), .Z(n11) );
  HS65_LS_IVX9 U43 ( .A(data_in[11]), .Z(n7) );
  HS65_LS_CB4I6X9 U44 ( .A(n2), .B(n1), .C(data_valid), .D(preset), .Z(N19) );
  HS65_LS_IVX9 U45 ( .A(data_in_34), .Z(n1) );
endmodule


module latch_controller_1_6 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_6 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_6 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n7) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_IVX9 U3 ( .A(N0), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_1_x_2 ( preset, .chan_in_f({\chan_in_f[REQ] , \chan_in_f[DATA][34] , 
        \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , 
        \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , 
        \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , 
        \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , 
        \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , 
        \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , 
        \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , 
        \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , 
        \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , 
        \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , 
        \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , 
        \chan_in_f[DATA][0] }), .chan_in_b(\chan_in_b[ACK] ), .chan_out_f({
        \chan_out_f[REQ] , \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , 
        \chan_out_f[DATA][32] , \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , 
        \chan_out_f[DATA][29] , \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , 
        \chan_out_f[DATA][26] , \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , 
        \chan_out_f[DATA][23] , \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , 
        \chan_out_f[DATA][20] , \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , 
        \chan_out_f[DATA][17] , \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , 
        \chan_out_f[DATA][14] , \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , 
        \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , 
        \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , 
        \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , 
        \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), 
    .chan_out_b(\chan_out_b[ACK] ), sel );
  output [4:0] sel;
  input preset, \chan_in_f[REQ] , \chan_in_f[DATA][34] , \chan_in_f[DATA][33] ,
         \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , \chan_in_f[DATA][30] ,
         \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , \chan_in_f[DATA][27] ,
         \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , \chan_in_f[DATA][24] ,
         \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , \chan_in_f[DATA][21] ,
         \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , \chan_in_f[DATA][18] ,
         \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , \chan_in_f[DATA][15] ,
         \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , \chan_in_f[DATA][12] ,
         \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , \chan_in_f[DATA][9] ,
         \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , \chan_in_f[DATA][6] ,
         \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , \chan_in_f[DATA][3] ,
         \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , \chan_in_f[DATA][0] ,
         \chan_out_b[ACK] ;
  output \chan_in_b[ACK] , \chan_out_f[REQ] , \chan_out_f[DATA][34] ,
         \chan_out_f[DATA][33] , \chan_out_f[DATA][32] ,
         \chan_out_f[DATA][31] , \chan_out_f[DATA][30] ,
         \chan_out_f[DATA][29] , \chan_out_f[DATA][28] ,
         \chan_out_f[DATA][27] , \chan_out_f[DATA][26] ,
         \chan_out_f[DATA][25] , \chan_out_f[DATA][24] ,
         \chan_out_f[DATA][23] , \chan_out_f[DATA][22] ,
         \chan_out_f[DATA][21] , \chan_out_f[DATA][20] ,
         \chan_out_f[DATA][19] , \chan_out_f[DATA][18] ,
         \chan_out_f[DATA][17] , \chan_out_f[DATA][16] ,
         \chan_out_f[DATA][15] , \chan_out_f[DATA][14] ,
         \chan_out_f[DATA][13] , \chan_out_f[DATA][12] ,
         \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] ,
         \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] ,
         \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] ,
         \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] ;
  wire   \chan_internal_f[REQ] , \chan_internal_f[DATA][34] ,
         \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] ,
         \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] ,
         \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] ,
         \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] ,
         \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] ,
         \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] ,
         \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] ,
         \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] ,
         \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] ,
         \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] ,
         \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] ,
         \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] ,
         \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] ,
         \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] ,
         \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] ,
         \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] ,
         \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] , req_n, lt_en,
         n1, n2, n3, n4, n5, n6, n7;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign sel[4] = 1'b0;

  hpu_comb_1_x_2 hpu_combinatorial ( .data_valid(lt_en), .data_in({
        \chan_in_f[DATA][34] , \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , 
        \chan_in_f[DATA][31] , \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , 
        \chan_in_f[DATA][28] , \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , 
        \chan_in_f[DATA][25] , \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , 
        \chan_in_f[DATA][22] , \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , 
        \chan_in_f[DATA][19] , \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , 
        \chan_in_f[DATA][16] , \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , 
        \chan_in_f[DATA][13] , \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , 
        \chan_in_f[DATA][10] , \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , 
        \chan_in_f[DATA][7] , \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , 
        \chan_in_f[DATA][4] , \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , 
        \chan_in_f[DATA][1] , \chan_in_f[DATA][0] }), .preset(n7), .data_out({
        \chan_internal_f[DATA][34] , \chan_internal_f[DATA][33] , 
        \chan_internal_f[DATA][32] , \chan_internal_f[DATA][31] , 
        \chan_internal_f[DATA][30] , \chan_internal_f[DATA][29] , 
        \chan_internal_f[DATA][28] , \chan_internal_f[DATA][27] , 
        \chan_internal_f[DATA][26] , \chan_internal_f[DATA][25] , 
        \chan_internal_f[DATA][24] , \chan_internal_f[DATA][23] , 
        \chan_internal_f[DATA][22] , \chan_internal_f[DATA][21] , 
        \chan_internal_f[DATA][20] , \chan_internal_f[DATA][19] , 
        \chan_internal_f[DATA][18] , \chan_internal_f[DATA][17] , 
        \chan_internal_f[DATA][16] , \chan_internal_f[DATA][15] , 
        \chan_internal_f[DATA][14] , \chan_internal_f[DATA][13] , 
        \chan_internal_f[DATA][12] , \chan_internal_f[DATA][11] , 
        \chan_internal_f[DATA][10] , \chan_internal_f[DATA][9] , 
        \chan_internal_f[DATA][8] , \chan_internal_f[DATA][7] , 
        \chan_internal_f[DATA][6] , \chan_internal_f[DATA][5] , 
        \chan_internal_f[DATA][4] , \chan_internal_f[DATA][3] , 
        \chan_internal_f[DATA][2] , \chan_internal_f[DATA][1] , 
        \chan_internal_f[DATA][0] }), .sel({SYNOPSYS_UNCONNECTED__0, sel[3:0]}) );
  channel_latch_1_xxxxxxxxx_6 token_latch ( .preset(n7), .left_in({
        \chan_internal_f[REQ] , \chan_internal_f[DATA][34] , 
        \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] , 
        \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] , 
        \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] , 
        \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] , 
        \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] , 
        \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] , 
        \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] , 
        \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] , 
        \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] , 
        \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] , 
        \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] , 
        \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] , 
        \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] , 
        \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] , 
        \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] , 
        \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] , 
        \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] }), .left_out(
        \chan_in_b[ACK] ), .right_out({\chan_out_f[REQ] , 
        \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , \chan_out_f[DATA][32] , 
        \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , \chan_out_f[DATA][29] , 
        \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , \chan_out_f[DATA][26] , 
        \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , \chan_out_f[DATA][23] , 
        \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , \chan_out_f[DATA][20] , 
        \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , \chan_out_f[DATA][17] , 
        \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , \chan_out_f[DATA][14] , 
        \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , \chan_out_f[DATA][11] , 
        \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , \chan_out_f[DATA][8] , 
        \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , \chan_out_f[DATA][5] , 
        \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , \chan_out_f[DATA][2] , 
        \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), .right_in(
        \chan_out_b[ACK] ), .lt_enable(lt_en) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chan_internal_f[REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(\chan_in_f[REQ] ), .Z(req_n) );
  HS65_LS_BFX9 U1 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U2 ( .A(n3), .Z(n2) );
  HS65_LS_BFX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_BFX9 U4 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U6 ( .A(req_n), .Z(n6) );
  HS65_LS_BFX9 U7 ( .A(preset), .Z(n7) );
endmodule


module sr_latch_1_4 ( s, r, q, qn );
  input s, r;
  output q, qn;
  wire   N3, n1;

  HS65_LS_AND2X4 C9 ( .A(n1), .B(N3), .Z(qn) );
  HS65_LH_NOR2X3 U1 ( .A(r), .B(qn), .Z(q) );
  HS65_LS_IVX9 U2 ( .A(q), .Z(N3) );
  HS65_LS_IVX9 U3 ( .A(s), .Z(n1) );
endmodule


module c_gate_generic_1_5_4 ( preset, \input , \output  );
  input [4:0] \input ;
  input preset;
  output \output ;
  wire   set, reset, n1, n4, n5;

  sr_latch_1_4 latch ( .s(set), .r(reset), .q(\output ) );
  HS65_LS_NOR3X4 U3 ( .A(\input [3]), .B(preset), .C(\input [4]), .Z(n4) );
  HS65_LS_NOR4ABX2 U4 ( .A(n1), .B(n4), .C(\input [2]), .D(\input [1]), .Z(
        reset) );
  HS65_LS_AO31X9 U5 ( .A(n5), .B(\input [3]), .C(\input [4]), .D(preset), .Z(
        set) );
  HS65_LS_IVX9 U6 ( .A(\input [0]), .Z(n1) );
  HS65_LS_AND3X9 U7 ( .A(\input [1]), .B(\input [0]), .C(\input [2]), .Z(n5)
         );
endmodule


module sr_latch_1_3 ( s, r, q, qn );
  input s, r;
  output q, qn;
  wire   N3, n1;

  HS65_LS_AND2X4 C9 ( .A(n1), .B(N3), .Z(qn) );
  HS65_LS_IVX9 U1 ( .A(q), .Z(N3) );
  HS65_LS_IVX9 U2 ( .A(s), .Z(n1) );
  HS65_LS_NOR2X6 U3 ( .A(r), .B(qn), .Z(q) );
endmodule


module c_gate_generic_1_5_3 ( preset, \input , \output  );
  input [4:0] \input ;
  input preset;
  output \output ;
  wire   set, reset, n1, n4, n5;

  sr_latch_1_3 latch ( .s(set), .r(reset), .q(\output ) );
  HS65_LS_NOR3X4 U3 ( .A(\input [3]), .B(preset), .C(\input [4]), .Z(n4) );
  HS65_LS_NOR4ABX2 U4 ( .A(n1), .B(n4), .C(\input [2]), .D(\input [1]), .Z(
        reset) );
  HS65_LS_AO31X9 U5 ( .A(n5), .B(\input [3]), .C(\input [4]), .D(preset), .Z(
        set) );
  HS65_LS_IVX9 U6 ( .A(\input [0]), .Z(n1) );
  HS65_LS_AND3X9 U7 ( .A(\input [1]), .B(\input [0]), .C(\input [2]), .Z(n5)
         );
endmodule


module crossbar_2 ( preset, .switch_sel({\switch_sel[4][4] , 
        \switch_sel[4][3] , \switch_sel[4][2] , \switch_sel[4][1] , 
        \switch_sel[4][0] , \switch_sel[3][4] , \switch_sel[3][3] , 
        \switch_sel[3][2] , \switch_sel[3][1] , \switch_sel[3][0] , 
        \switch_sel[2][4] , \switch_sel[2][3] , \switch_sel[2][2] , 
        \switch_sel[2][1] , \switch_sel[2][0] , \switch_sel[1][4] , 
        \switch_sel[1][3] , \switch_sel[1][2] , \switch_sel[1][1] , 
        \switch_sel[1][0] , \switch_sel[0][4] , \switch_sel[0][3] , 
        \switch_sel[0][2] , \switch_sel[0][1] , \switch_sel[0][0] }), 
    .chs_in_f({\chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] , 
        \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] , 
        \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] , 
        \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] , 
        \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] , 
        \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] , 
        \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] , 
        \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] , 
        \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] , 
        \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] , 
        \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] , 
        \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] , 
        \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] , 
        \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] , \chs_in_f[4][DATA][7] , 
        \chs_in_f[4][DATA][6] , \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] , 
        \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] , \chs_in_f[4][DATA][1] , 
        \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] , \chs_in_f[3][DATA][34] , 
        \chs_in_f[3][DATA][33] , \chs_in_f[3][DATA][32] , 
        \chs_in_f[3][DATA][31] , \chs_in_f[3][DATA][30] , 
        \chs_in_f[3][DATA][29] , \chs_in_f[3][DATA][28] , 
        \chs_in_f[3][DATA][27] , \chs_in_f[3][DATA][26] , 
        \chs_in_f[3][DATA][25] , \chs_in_f[3][DATA][24] , 
        \chs_in_f[3][DATA][23] , \chs_in_f[3][DATA][22] , 
        \chs_in_f[3][DATA][21] , \chs_in_f[3][DATA][20] , 
        \chs_in_f[3][DATA][19] , \chs_in_f[3][DATA][18] , 
        \chs_in_f[3][DATA][17] , \chs_in_f[3][DATA][16] , 
        \chs_in_f[3][DATA][15] , \chs_in_f[3][DATA][14] , 
        \chs_in_f[3][DATA][13] , \chs_in_f[3][DATA][12] , 
        \chs_in_f[3][DATA][11] , \chs_in_f[3][DATA][10] , 
        \chs_in_f[3][DATA][9] , \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] , 
        \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] , \chs_in_f[3][DATA][4] , 
        \chs_in_f[3][DATA][3] , \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] , 
        \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] , 
        \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] , 
        \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] , 
        \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] , 
        \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] , 
        \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] , 
        \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] , 
        \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] , 
        \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] , 
        \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] , 
        \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] , 
        \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] , 
        \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] , 
        \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] , \chs_in_f[2][DATA][7] , 
        \chs_in_f[2][DATA][6] , \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] , 
        \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] , \chs_in_f[2][DATA][1] , 
        \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] , \chs_in_f[1][DATA][34] , 
        \chs_in_f[1][DATA][33] , \chs_in_f[1][DATA][32] , 
        \chs_in_f[1][DATA][31] , \chs_in_f[1][DATA][30] , 
        \chs_in_f[1][DATA][29] , \chs_in_f[1][DATA][28] , 
        \chs_in_f[1][DATA][27] , \chs_in_f[1][DATA][26] , 
        \chs_in_f[1][DATA][25] , \chs_in_f[1][DATA][24] , 
        \chs_in_f[1][DATA][23] , \chs_in_f[1][DATA][22] , 
        \chs_in_f[1][DATA][21] , \chs_in_f[1][DATA][20] , 
        \chs_in_f[1][DATA][19] , \chs_in_f[1][DATA][18] , 
        \chs_in_f[1][DATA][17] , \chs_in_f[1][DATA][16] , 
        \chs_in_f[1][DATA][15] , \chs_in_f[1][DATA][14] , 
        \chs_in_f[1][DATA][13] , \chs_in_f[1][DATA][12] , 
        \chs_in_f[1][DATA][11] , \chs_in_f[1][DATA][10] , 
        \chs_in_f[1][DATA][9] , \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] , 
        \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] , \chs_in_f[1][DATA][4] , 
        \chs_in_f[1][DATA][3] , \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] , 
        \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] , 
        \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] , 
        \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] , 
        \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] , 
        \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] , 
        \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] , 
        \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] , 
        \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] , 
        \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] , 
        \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] , 
        \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] , 
        \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] , 
        \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] , 
        \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] , \chs_in_f[0][DATA][7] , 
        \chs_in_f[0][DATA][6] , \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] , 
        \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] , \chs_in_f[0][DATA][1] , 
        \chs_in_f[0][DATA][0] }), .chs_in_b({\chs_in_b[4][ACK] , 
        \chs_in_b[3][ACK] , \chs_in_b[2][ACK] , \chs_in_b[1][ACK] , 
        \chs_in_b[0][ACK] }), .chs_out_f({\chs_out_f[4][REQ] , 
        \chs_out_f[4][DATA][34] , \chs_out_f[4][DATA][33] , 
        \chs_out_f[4][DATA][32] , \chs_out_f[4][DATA][31] , 
        \chs_out_f[4][DATA][30] , \chs_out_f[4][DATA][29] , 
        \chs_out_f[4][DATA][28] , \chs_out_f[4][DATA][27] , 
        \chs_out_f[4][DATA][26] , \chs_out_f[4][DATA][25] , 
        \chs_out_f[4][DATA][24] , \chs_out_f[4][DATA][23] , 
        \chs_out_f[4][DATA][22] , \chs_out_f[4][DATA][21] , 
        \chs_out_f[4][DATA][20] , \chs_out_f[4][DATA][19] , 
        \chs_out_f[4][DATA][18] , \chs_out_f[4][DATA][17] , 
        \chs_out_f[4][DATA][16] , \chs_out_f[4][DATA][15] , 
        \chs_out_f[4][DATA][14] , \chs_out_f[4][DATA][13] , 
        \chs_out_f[4][DATA][12] , \chs_out_f[4][DATA][11] , 
        \chs_out_f[4][DATA][10] , \chs_out_f[4][DATA][9] , 
        \chs_out_f[4][DATA][8] , \chs_out_f[4][DATA][7] , 
        \chs_out_f[4][DATA][6] , \chs_out_f[4][DATA][5] , 
        \chs_out_f[4][DATA][4] , \chs_out_f[4][DATA][3] , 
        \chs_out_f[4][DATA][2] , \chs_out_f[4][DATA][1] , 
        \chs_out_f[4][DATA][0] , \chs_out_f[3][REQ] , \chs_out_f[3][DATA][34] , 
        \chs_out_f[3][DATA][33] , \chs_out_f[3][DATA][32] , 
        \chs_out_f[3][DATA][31] , \chs_out_f[3][DATA][30] , 
        \chs_out_f[3][DATA][29] , \chs_out_f[3][DATA][28] , 
        \chs_out_f[3][DATA][27] , \chs_out_f[3][DATA][26] , 
        \chs_out_f[3][DATA][25] , \chs_out_f[3][DATA][24] , 
        \chs_out_f[3][DATA][23] , \chs_out_f[3][DATA][22] , 
        \chs_out_f[3][DATA][21] , \chs_out_f[3][DATA][20] , 
        \chs_out_f[3][DATA][19] , \chs_out_f[3][DATA][18] , 
        \chs_out_f[3][DATA][17] , \chs_out_f[3][DATA][16] , 
        \chs_out_f[3][DATA][15] , \chs_out_f[3][DATA][14] , 
        \chs_out_f[3][DATA][13] , \chs_out_f[3][DATA][12] , 
        \chs_out_f[3][DATA][11] , \chs_out_f[3][DATA][10] , 
        \chs_out_f[3][DATA][9] , \chs_out_f[3][DATA][8] , 
        \chs_out_f[3][DATA][7] , \chs_out_f[3][DATA][6] , 
        \chs_out_f[3][DATA][5] , \chs_out_f[3][DATA][4] , 
        \chs_out_f[3][DATA][3] , \chs_out_f[3][DATA][2] , 
        \chs_out_f[3][DATA][1] , \chs_out_f[3][DATA][0] , \chs_out_f[2][REQ] , 
        \chs_out_f[2][DATA][34] , \chs_out_f[2][DATA][33] , 
        \chs_out_f[2][DATA][32] , \chs_out_f[2][DATA][31] , 
        \chs_out_f[2][DATA][30] , \chs_out_f[2][DATA][29] , 
        \chs_out_f[2][DATA][28] , \chs_out_f[2][DATA][27] , 
        \chs_out_f[2][DATA][26] , \chs_out_f[2][DATA][25] , 
        \chs_out_f[2][DATA][24] , \chs_out_f[2][DATA][23] , 
        \chs_out_f[2][DATA][22] , \chs_out_f[2][DATA][21] , 
        \chs_out_f[2][DATA][20] , \chs_out_f[2][DATA][19] , 
        \chs_out_f[2][DATA][18] , \chs_out_f[2][DATA][17] , 
        \chs_out_f[2][DATA][16] , \chs_out_f[2][DATA][15] , 
        \chs_out_f[2][DATA][14] , \chs_out_f[2][DATA][13] , 
        \chs_out_f[2][DATA][12] , \chs_out_f[2][DATA][11] , 
        \chs_out_f[2][DATA][10] , \chs_out_f[2][DATA][9] , 
        \chs_out_f[2][DATA][8] , \chs_out_f[2][DATA][7] , 
        \chs_out_f[2][DATA][6] , \chs_out_f[2][DATA][5] , 
        \chs_out_f[2][DATA][4] , \chs_out_f[2][DATA][3] , 
        \chs_out_f[2][DATA][2] , \chs_out_f[2][DATA][1] , 
        \chs_out_f[2][DATA][0] , \chs_out_f[1][REQ] , \chs_out_f[1][DATA][34] , 
        \chs_out_f[1][DATA][33] , \chs_out_f[1][DATA][32] , 
        \chs_out_f[1][DATA][31] , \chs_out_f[1][DATA][30] , 
        \chs_out_f[1][DATA][29] , \chs_out_f[1][DATA][28] , 
        \chs_out_f[1][DATA][27] , \chs_out_f[1][DATA][26] , 
        \chs_out_f[1][DATA][25] , \chs_out_f[1][DATA][24] , 
        \chs_out_f[1][DATA][23] , \chs_out_f[1][DATA][22] , 
        \chs_out_f[1][DATA][21] , \chs_out_f[1][DATA][20] , 
        \chs_out_f[1][DATA][19] , \chs_out_f[1][DATA][18] , 
        \chs_out_f[1][DATA][17] , \chs_out_f[1][DATA][16] , 
        \chs_out_f[1][DATA][15] , \chs_out_f[1][DATA][14] , 
        \chs_out_f[1][DATA][13] , \chs_out_f[1][DATA][12] , 
        \chs_out_f[1][DATA][11] , \chs_out_f[1][DATA][10] , 
        \chs_out_f[1][DATA][9] , \chs_out_f[1][DATA][8] , 
        \chs_out_f[1][DATA][7] , \chs_out_f[1][DATA][6] , 
        \chs_out_f[1][DATA][5] , \chs_out_f[1][DATA][4] , 
        \chs_out_f[1][DATA][3] , \chs_out_f[1][DATA][2] , 
        \chs_out_f[1][DATA][1] , \chs_out_f[1][DATA][0] , \chs_out_f[0][REQ] , 
        \chs_out_f[0][DATA][34] , \chs_out_f[0][DATA][33] , 
        \chs_out_f[0][DATA][32] , \chs_out_f[0][DATA][31] , 
        \chs_out_f[0][DATA][30] , \chs_out_f[0][DATA][29] , 
        \chs_out_f[0][DATA][28] , \chs_out_f[0][DATA][27] , 
        \chs_out_f[0][DATA][26] , \chs_out_f[0][DATA][25] , 
        \chs_out_f[0][DATA][24] , \chs_out_f[0][DATA][23] , 
        \chs_out_f[0][DATA][22] , \chs_out_f[0][DATA][21] , 
        \chs_out_f[0][DATA][20] , \chs_out_f[0][DATA][19] , 
        \chs_out_f[0][DATA][18] , \chs_out_f[0][DATA][17] , 
        \chs_out_f[0][DATA][16] , \chs_out_f[0][DATA][15] , 
        \chs_out_f[0][DATA][14] , \chs_out_f[0][DATA][13] , 
        \chs_out_f[0][DATA][12] , \chs_out_f[0][DATA][11] , 
        \chs_out_f[0][DATA][10] , \chs_out_f[0][DATA][9] , 
        \chs_out_f[0][DATA][8] , \chs_out_f[0][DATA][7] , 
        \chs_out_f[0][DATA][6] , \chs_out_f[0][DATA][5] , 
        \chs_out_f[0][DATA][4] , \chs_out_f[0][DATA][3] , 
        \chs_out_f[0][DATA][2] , \chs_out_f[0][DATA][1] , 
        \chs_out_f[0][DATA][0] }), .chs_out_b({\chs_out_b[4][ACK] , 
        \chs_out_b[3][ACK] , \chs_out_b[2][ACK] , \chs_out_b[1][ACK] , 
        \chs_out_b[0][ACK] }) );
  input preset, \switch_sel[4][4] , \switch_sel[4][3] , \switch_sel[4][2] ,
         \switch_sel[4][1] , \switch_sel[4][0] , \switch_sel[3][4] ,
         \switch_sel[3][3] , \switch_sel[3][2] , \switch_sel[3][1] ,
         \switch_sel[3][0] , \switch_sel[2][4] , \switch_sel[2][3] ,
         \switch_sel[2][2] , \switch_sel[2][1] , \switch_sel[2][0] ,
         \switch_sel[1][4] , \switch_sel[1][3] , \switch_sel[1][2] ,
         \switch_sel[1][1] , \switch_sel[1][0] , \switch_sel[0][4] ,
         \switch_sel[0][3] , \switch_sel[0][2] , \switch_sel[0][1] ,
         \switch_sel[0][0] , \chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] ,
         \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] ,
         \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] ,
         \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] ,
         \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] ,
         \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] ,
         \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] ,
         \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] ,
         \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] ,
         \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] ,
         \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] ,
         \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] ,
         \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] ,
         \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] ,
         \chs_in_f[4][DATA][7] , \chs_in_f[4][DATA][6] ,
         \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] ,
         \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] ,
         \chs_in_f[4][DATA][1] , \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] ,
         \chs_in_f[3][DATA][34] , \chs_in_f[3][DATA][33] ,
         \chs_in_f[3][DATA][32] , \chs_in_f[3][DATA][31] ,
         \chs_in_f[3][DATA][30] , \chs_in_f[3][DATA][29] ,
         \chs_in_f[3][DATA][28] , \chs_in_f[3][DATA][27] ,
         \chs_in_f[3][DATA][26] , \chs_in_f[3][DATA][25] ,
         \chs_in_f[3][DATA][24] , \chs_in_f[3][DATA][23] ,
         \chs_in_f[3][DATA][22] , \chs_in_f[3][DATA][21] ,
         \chs_in_f[3][DATA][20] , \chs_in_f[3][DATA][19] ,
         \chs_in_f[3][DATA][18] , \chs_in_f[3][DATA][17] ,
         \chs_in_f[3][DATA][16] , \chs_in_f[3][DATA][15] ,
         \chs_in_f[3][DATA][14] , \chs_in_f[3][DATA][13] ,
         \chs_in_f[3][DATA][12] , \chs_in_f[3][DATA][11] ,
         \chs_in_f[3][DATA][10] , \chs_in_f[3][DATA][9] ,
         \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] ,
         \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] ,
         \chs_in_f[3][DATA][4] , \chs_in_f[3][DATA][3] ,
         \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] ,
         \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] ,
         \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] ,
         \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] ,
         \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] ,
         \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] ,
         \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] ,
         \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] ,
         \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] ,
         \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] ,
         \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] ,
         \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] ,
         \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] ,
         \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] ,
         \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] ,
         \chs_in_f[2][DATA][7] , \chs_in_f[2][DATA][6] ,
         \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] ,
         \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] ,
         \chs_in_f[2][DATA][1] , \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] ,
         \chs_in_f[1][DATA][34] , \chs_in_f[1][DATA][33] ,
         \chs_in_f[1][DATA][32] , \chs_in_f[1][DATA][31] ,
         \chs_in_f[1][DATA][30] , \chs_in_f[1][DATA][29] ,
         \chs_in_f[1][DATA][28] , \chs_in_f[1][DATA][27] ,
         \chs_in_f[1][DATA][26] , \chs_in_f[1][DATA][25] ,
         \chs_in_f[1][DATA][24] , \chs_in_f[1][DATA][23] ,
         \chs_in_f[1][DATA][22] , \chs_in_f[1][DATA][21] ,
         \chs_in_f[1][DATA][20] , \chs_in_f[1][DATA][19] ,
         \chs_in_f[1][DATA][18] , \chs_in_f[1][DATA][17] ,
         \chs_in_f[1][DATA][16] , \chs_in_f[1][DATA][15] ,
         \chs_in_f[1][DATA][14] , \chs_in_f[1][DATA][13] ,
         \chs_in_f[1][DATA][12] , \chs_in_f[1][DATA][11] ,
         \chs_in_f[1][DATA][10] , \chs_in_f[1][DATA][9] ,
         \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] ,
         \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] ,
         \chs_in_f[1][DATA][4] , \chs_in_f[1][DATA][3] ,
         \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] ,
         \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] ,
         \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] ,
         \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] ,
         \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] ,
         \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] ,
         \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] ,
         \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] ,
         \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] ,
         \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] ,
         \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] ,
         \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] ,
         \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] ,
         \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] ,
         \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] ,
         \chs_in_f[0][DATA][7] , \chs_in_f[0][DATA][6] ,
         \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] ,
         \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] ,
         \chs_in_f[0][DATA][1] , \chs_in_f[0][DATA][0] , \chs_out_b[4][ACK] ,
         \chs_out_b[3][ACK] , \chs_out_b[2][ACK] , \chs_out_b[1][ACK] ,
         \chs_out_b[0][ACK] ;
  output \chs_in_b[4][ACK] , \chs_in_b[3][ACK] , \chs_in_b[2][ACK] ,
         \chs_in_b[1][ACK] , \chs_in_b[0][ACK] , \chs_out_f[4][REQ] ,
         \chs_out_f[4][DATA][34] , \chs_out_f[4][DATA][33] ,
         \chs_out_f[4][DATA][32] , \chs_out_f[4][DATA][31] ,
         \chs_out_f[4][DATA][30] , \chs_out_f[4][DATA][29] ,
         \chs_out_f[4][DATA][28] , \chs_out_f[4][DATA][27] ,
         \chs_out_f[4][DATA][26] , \chs_out_f[4][DATA][25] ,
         \chs_out_f[4][DATA][24] , \chs_out_f[4][DATA][23] ,
         \chs_out_f[4][DATA][22] , \chs_out_f[4][DATA][21] ,
         \chs_out_f[4][DATA][20] , \chs_out_f[4][DATA][19] ,
         \chs_out_f[4][DATA][18] , \chs_out_f[4][DATA][17] ,
         \chs_out_f[4][DATA][16] , \chs_out_f[4][DATA][15] ,
         \chs_out_f[4][DATA][14] , \chs_out_f[4][DATA][13] ,
         \chs_out_f[4][DATA][12] , \chs_out_f[4][DATA][11] ,
         \chs_out_f[4][DATA][10] , \chs_out_f[4][DATA][9] ,
         \chs_out_f[4][DATA][8] , \chs_out_f[4][DATA][7] ,
         \chs_out_f[4][DATA][6] , \chs_out_f[4][DATA][5] ,
         \chs_out_f[4][DATA][4] , \chs_out_f[4][DATA][3] ,
         \chs_out_f[4][DATA][2] , \chs_out_f[4][DATA][1] ,
         \chs_out_f[4][DATA][0] , \chs_out_f[3][REQ] ,
         \chs_out_f[3][DATA][34] , \chs_out_f[3][DATA][33] ,
         \chs_out_f[3][DATA][32] , \chs_out_f[3][DATA][31] ,
         \chs_out_f[3][DATA][30] , \chs_out_f[3][DATA][29] ,
         \chs_out_f[3][DATA][28] , \chs_out_f[3][DATA][27] ,
         \chs_out_f[3][DATA][26] , \chs_out_f[3][DATA][25] ,
         \chs_out_f[3][DATA][24] , \chs_out_f[3][DATA][23] ,
         \chs_out_f[3][DATA][22] , \chs_out_f[3][DATA][21] ,
         \chs_out_f[3][DATA][20] , \chs_out_f[3][DATA][19] ,
         \chs_out_f[3][DATA][18] , \chs_out_f[3][DATA][17] ,
         \chs_out_f[3][DATA][16] , \chs_out_f[3][DATA][15] ,
         \chs_out_f[3][DATA][14] , \chs_out_f[3][DATA][13] ,
         \chs_out_f[3][DATA][12] , \chs_out_f[3][DATA][11] ,
         \chs_out_f[3][DATA][10] , \chs_out_f[3][DATA][9] ,
         \chs_out_f[3][DATA][8] , \chs_out_f[3][DATA][7] ,
         \chs_out_f[3][DATA][6] , \chs_out_f[3][DATA][5] ,
         \chs_out_f[3][DATA][4] , \chs_out_f[3][DATA][3] ,
         \chs_out_f[3][DATA][2] , \chs_out_f[3][DATA][1] ,
         \chs_out_f[3][DATA][0] , \chs_out_f[2][REQ] ,
         \chs_out_f[2][DATA][34] , \chs_out_f[2][DATA][33] ,
         \chs_out_f[2][DATA][32] , \chs_out_f[2][DATA][31] ,
         \chs_out_f[2][DATA][30] , \chs_out_f[2][DATA][29] ,
         \chs_out_f[2][DATA][28] , \chs_out_f[2][DATA][27] ,
         \chs_out_f[2][DATA][26] , \chs_out_f[2][DATA][25] ,
         \chs_out_f[2][DATA][24] , \chs_out_f[2][DATA][23] ,
         \chs_out_f[2][DATA][22] , \chs_out_f[2][DATA][21] ,
         \chs_out_f[2][DATA][20] , \chs_out_f[2][DATA][19] ,
         \chs_out_f[2][DATA][18] , \chs_out_f[2][DATA][17] ,
         \chs_out_f[2][DATA][16] , \chs_out_f[2][DATA][15] ,
         \chs_out_f[2][DATA][14] , \chs_out_f[2][DATA][13] ,
         \chs_out_f[2][DATA][12] , \chs_out_f[2][DATA][11] ,
         \chs_out_f[2][DATA][10] , \chs_out_f[2][DATA][9] ,
         \chs_out_f[2][DATA][8] , \chs_out_f[2][DATA][7] ,
         \chs_out_f[2][DATA][6] , \chs_out_f[2][DATA][5] ,
         \chs_out_f[2][DATA][4] , \chs_out_f[2][DATA][3] ,
         \chs_out_f[2][DATA][2] , \chs_out_f[2][DATA][1] ,
         \chs_out_f[2][DATA][0] , \chs_out_f[1][REQ] ,
         \chs_out_f[1][DATA][34] , \chs_out_f[1][DATA][33] ,
         \chs_out_f[1][DATA][32] , \chs_out_f[1][DATA][31] ,
         \chs_out_f[1][DATA][30] , \chs_out_f[1][DATA][29] ,
         \chs_out_f[1][DATA][28] , \chs_out_f[1][DATA][27] ,
         \chs_out_f[1][DATA][26] , \chs_out_f[1][DATA][25] ,
         \chs_out_f[1][DATA][24] , \chs_out_f[1][DATA][23] ,
         \chs_out_f[1][DATA][22] , \chs_out_f[1][DATA][21] ,
         \chs_out_f[1][DATA][20] , \chs_out_f[1][DATA][19] ,
         \chs_out_f[1][DATA][18] , \chs_out_f[1][DATA][17] ,
         \chs_out_f[1][DATA][16] , \chs_out_f[1][DATA][15] ,
         \chs_out_f[1][DATA][14] , \chs_out_f[1][DATA][13] ,
         \chs_out_f[1][DATA][12] , \chs_out_f[1][DATA][11] ,
         \chs_out_f[1][DATA][10] , \chs_out_f[1][DATA][9] ,
         \chs_out_f[1][DATA][8] , \chs_out_f[1][DATA][7] ,
         \chs_out_f[1][DATA][6] , \chs_out_f[1][DATA][5] ,
         \chs_out_f[1][DATA][4] , \chs_out_f[1][DATA][3] ,
         \chs_out_f[1][DATA][2] , \chs_out_f[1][DATA][1] ,
         \chs_out_f[1][DATA][0] , \chs_out_f[0][REQ] ,
         \chs_out_f[0][DATA][34] , \chs_out_f[0][DATA][33] ,
         \chs_out_f[0][DATA][32] , \chs_out_f[0][DATA][31] ,
         \chs_out_f[0][DATA][30] , \chs_out_f[0][DATA][29] ,
         \chs_out_f[0][DATA][28] , \chs_out_f[0][DATA][27] ,
         \chs_out_f[0][DATA][26] , \chs_out_f[0][DATA][25] ,
         \chs_out_f[0][DATA][24] , \chs_out_f[0][DATA][23] ,
         \chs_out_f[0][DATA][22] , \chs_out_f[0][DATA][21] ,
         \chs_out_f[0][DATA][20] , \chs_out_f[0][DATA][19] ,
         \chs_out_f[0][DATA][18] , \chs_out_f[0][DATA][17] ,
         \chs_out_f[0][DATA][16] , \chs_out_f[0][DATA][15] ,
         \chs_out_f[0][DATA][14] , \chs_out_f[0][DATA][13] ,
         \chs_out_f[0][DATA][12] , \chs_out_f[0][DATA][11] ,
         \chs_out_f[0][DATA][10] , \chs_out_f[0][DATA][9] ,
         \chs_out_f[0][DATA][8] , \chs_out_f[0][DATA][7] ,
         \chs_out_f[0][DATA][6] , \chs_out_f[0][DATA][5] ,
         \chs_out_f[0][DATA][4] , \chs_out_f[0][DATA][3] ,
         \chs_out_f[0][DATA][2] , \chs_out_f[0][DATA][1] ,
         \chs_out_f[0][DATA][0] ;
  wire   \chs_in_b[4][ACK] , \chs_out_f[4][REQ] , synced_req, del, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510;
  assign \chs_in_b[0][ACK]  = \chs_in_b[4][ACK] ;
  assign \chs_in_b[1][ACK]  = \chs_in_b[4][ACK] ;
  assign \chs_in_b[2][ACK]  = \chs_in_b[4][ACK] ;
  assign \chs_in_b[3][ACK]  = \chs_in_b[4][ACK] ;
  assign \chs_out_f[0][REQ]  = \chs_out_f[4][REQ] ;
  assign \chs_out_f[1][REQ]  = \chs_out_f[4][REQ] ;
  assign \chs_out_f[2][REQ]  = \chs_out_f[4][REQ] ;
  assign \chs_out_f[3][REQ]  = \chs_out_f[4][REQ] ;

  c_gate_generic_1_5_4 c_sync_req ( .preset(preset), .\input ({
        \chs_in_f[4][REQ] , \chs_in_f[3][REQ] , \chs_in_f[2][REQ] , 
        \chs_in_f[1][REQ] , \chs_in_f[0][REQ] }), .\output (synced_req) );
  c_gate_generic_1_5_3 c_sync_ack ( .preset(preset), .\input ({
        \chs_out_b[4][ACK] , \chs_out_b[3][ACK] , \chs_out_b[2][ACK] , 
        \chs_out_b[1][ACK] , \chs_out_b[0][ACK] }), .\output (
        \chs_in_b[4][ACK] ) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chs_out_f[4][REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(synced_req), .Z(del) );
  HS65_LS_IVX9 U2 ( .A(\switch_sel[3][4] ), .Z(n261) );
  HS65_LS_IVX9 U3 ( .A(\switch_sel[3][2] ), .Z(n262) );
  HS65_LS_IVX9 U4 ( .A(\switch_sel[3][1] ), .Z(n263) );
  HS65_LS_IVX9 U5 ( .A(\switch_sel[3][0] ), .Z(n264) );
  HS65_LS_BFX9 U6 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U7 ( .A(del), .Z(n2) );
  HS65_LS_BFX9 U8 ( .A(n256), .Z(n5) );
  HS65_LS_BFX7 U9 ( .A(n259), .Z(n12) );
  HS65_LS_BFX7 U10 ( .A(n259), .Z(n13) );
  HS65_LS_BFX7 U11 ( .A(n257), .Z(n8) );
  HS65_LS_OAI212X3 U12 ( .A(n20), .B(n296), .C(n17), .D(n331), .E(n505), .Z(
        \chs_out_f[4][DATA][4] ) );
  HS65_LS_OAI212X3 U13 ( .A(n18), .B(n290), .C(n15), .D(n325), .E(n477), .Z(
        \chs_out_f[4][DATA][10] ) );
  HS65_LS_OAI212X3 U14 ( .A(n18), .B(n289), .C(n15), .D(n324), .E(n478), .Z(
        \chs_out_f[4][DATA][11] ) );
  HS65_LS_OAI212X3 U15 ( .A(n18), .B(n288), .C(n15), .D(n323), .E(n479), .Z(
        \chs_out_f[4][DATA][12] ) );
  HS65_LS_OAI212X3 U16 ( .A(n18), .B(n287), .C(n15), .D(n322), .E(n480), .Z(
        \chs_out_f[4][DATA][13] ) );
  HS65_LS_OAI212X3 U17 ( .A(n18), .B(n300), .C(n15), .D(n335), .E(n476), .Z(
        \chs_out_f[4][DATA][0] ) );
  HS65_LS_OAI212X3 U18 ( .A(n18), .B(n299), .C(n15), .D(n334), .E(n487), .Z(
        \chs_out_f[4][DATA][1] ) );
  HS65_LS_OAI212X3 U19 ( .A(n19), .B(n298), .C(n16), .D(n333), .E(n498), .Z(
        \chs_out_f[4][DATA][2] ) );
  HS65_LS_OAI212X3 U20 ( .A(n20), .B(n297), .C(n17), .D(n332), .E(n504), .Z(
        \chs_out_f[4][DATA][3] ) );
  HS65_LS_BFX9 U21 ( .A(\switch_sel[0][4] ), .Z(n45) );
  HS65_LS_BFX9 U22 ( .A(\switch_sel[1][4] ), .Z(n61) );
  HS65_LS_BFX9 U23 ( .A(\switch_sel[0][3] ), .Z(n41) );
  HS65_LS_BFX9 U24 ( .A(\switch_sel[1][3] ), .Z(n57) );
  HS65_LS_BFX9 U25 ( .A(\switch_sel[1][2] ), .Z(n53) );
  HS65_LS_BFX9 U26 ( .A(\switch_sel[0][1] ), .Z(n33) );
  HS65_LS_BFX9 U27 ( .A(\switch_sel[1][0] ), .Z(n49) );
  HS65_LS_BFX9 U28 ( .A(n261), .Z(n18) );
  HS65_LS_BFX9 U29 ( .A(n261), .Z(n19) );
  HS65_LS_BFX9 U30 ( .A(n61), .Z(n62) );
  HS65_LS_BFX9 U31 ( .A(n61), .Z(n63) );
  HS65_LS_BFX9 U32 ( .A(n77), .Z(n78) );
  HS65_LS_BFX9 U33 ( .A(n77), .Z(n79) );
  HS65_LS_BFX9 U34 ( .A(n45), .Z(n46) );
  HS65_LS_BFX9 U35 ( .A(n45), .Z(n47) );
  HS65_LS_BFX9 U36 ( .A(n262), .Z(n21) );
  HS65_LS_BFX9 U37 ( .A(n262), .Z(n22) );
  HS65_LS_BFX9 U38 ( .A(n263), .Z(n24) );
  HS65_LS_BFX9 U39 ( .A(n263), .Z(n25) );
  HS65_LS_BFX9 U40 ( .A(n264), .Z(n27) );
  HS65_LS_BFX9 U41 ( .A(n264), .Z(n28) );
  HS65_LS_BFX9 U42 ( .A(n57), .Z(n58) );
  HS65_LS_BFX9 U43 ( .A(n57), .Z(n59) );
  HS65_LS_BFX9 U44 ( .A(n53), .Z(n54) );
  HS65_LS_BFX9 U45 ( .A(n53), .Z(n55) );
  HS65_LS_BFX9 U46 ( .A(n49), .Z(n50) );
  HS65_LS_BFX9 U47 ( .A(n49), .Z(n51) );
  HS65_LS_BFX9 U48 ( .A(n73), .Z(n74) );
  HS65_LS_BFX9 U49 ( .A(n73), .Z(n75) );
  HS65_LS_BFX9 U50 ( .A(n69), .Z(n70) );
  HS65_LS_BFX9 U51 ( .A(n69), .Z(n71) );
  HS65_LS_BFX9 U52 ( .A(n65), .Z(n66) );
  HS65_LS_BFX9 U53 ( .A(n65), .Z(n67) );
  HS65_LS_BFX9 U54 ( .A(n261), .Z(n20) );
  HS65_LS_BFX9 U55 ( .A(n41), .Z(n42) );
  HS65_LS_BFX9 U56 ( .A(n41), .Z(n43) );
  HS65_LS_BFX9 U57 ( .A(n37), .Z(n38) );
  HS65_LS_BFX9 U58 ( .A(n37), .Z(n39) );
  HS65_LS_BFX9 U59 ( .A(n33), .Z(n34) );
  HS65_LS_BFX9 U60 ( .A(n33), .Z(n35) );
  HS65_LS_BFX9 U61 ( .A(n45), .Z(n48) );
  HS65_LS_BFX9 U62 ( .A(n257), .Z(n6) );
  HS65_LS_BFX9 U63 ( .A(n257), .Z(n7) );
  HS65_LS_BFX9 U64 ( .A(n258), .Z(n9) );
  HS65_LS_BFX9 U65 ( .A(n258), .Z(n10) );
  HS65_LS_BFX9 U66 ( .A(n256), .Z(n3) );
  HS65_LS_BFX9 U67 ( .A(n256), .Z(n4) );
  HS65_LS_BFX9 U68 ( .A(n57), .Z(n60) );
  HS65_LS_BFX9 U69 ( .A(n53), .Z(n56) );
  HS65_LS_BFX9 U70 ( .A(n49), .Z(n52) );
  HS65_LS_BFX9 U71 ( .A(n73), .Z(n76) );
  HS65_LS_BFX9 U72 ( .A(n69), .Z(n72) );
  HS65_LS_BFX9 U73 ( .A(n65), .Z(n68) );
  HS65_LS_BFX9 U74 ( .A(n41), .Z(n44) );
  HS65_LS_BFX9 U75 ( .A(n37), .Z(n40) );
  HS65_LS_BFX9 U76 ( .A(n33), .Z(n36) );
  HS65_LS_BFX9 U77 ( .A(n259), .Z(n14) );
  HS65_LS_BFX9 U78 ( .A(n258), .Z(n11) );
  HS65_LS_BFX9 U79 ( .A(n262), .Z(n23) );
  HS65_LS_BFX9 U80 ( .A(n263), .Z(n26) );
  HS65_LS_BFX9 U81 ( .A(n264), .Z(n29) );
  HS65_LS_BFX9 U82 ( .A(n61), .Z(n64) );
  HS65_LS_BFX9 U83 ( .A(n77), .Z(n80) );
  HS65_LS_BFX9 U84 ( .A(n260), .Z(n15) );
  HS65_LS_BFX9 U85 ( .A(n260), .Z(n16) );
  HS65_LS_BFX9 U86 ( .A(n265), .Z(n30) );
  HS65_LS_BFX9 U87 ( .A(n265), .Z(n31) );
  HS65_LS_BFX9 U88 ( .A(n260), .Z(n17) );
  HS65_LS_BFX9 U89 ( .A(n265), .Z(n32) );
  HS65_LS_IVX9 U90 ( .A(\switch_sel[4][2] ), .Z(n257) );
  HS65_LS_IVX9 U91 ( .A(\switch_sel[4][1] ), .Z(n258) );
  HS65_LS_IVX9 U92 ( .A(\switch_sel[4][3] ), .Z(n256) );
  HS65_LS_IVX9 U93 ( .A(\switch_sel[4][0] ), .Z(n259) );
  HS65_LS_AOI222X2 U94 ( .A(\chs_in_f[2][DATA][34] ), .B(n78), .C(
        \chs_in_f[0][DATA][34] ), .D(n48), .E(\chs_in_f[1][DATA][34] ), .F(n62), .Z(n503) );
  HS65_LS_OAI212X5 U95 ( .A(n291), .B(n20), .C(n326), .D(n17), .E(n510), .Z(
        \chs_out_f[4][DATA][9] ) );
  HS65_LS_AOI222X2 U96 ( .A(n78), .B(\chs_in_f[2][DATA][9] ), .C(n48), .D(
        \chs_in_f[0][DATA][9] ), .E(n62), .F(\chs_in_f[1][DATA][9] ), .Z(n510)
         );
  HS65_LS_AOI222X2 U97 ( .A(n76), .B(\chs_in_f[2][DATA][34] ), .C(n44), .D(
        \chs_in_f[0][DATA][34] ), .E(n60), .F(\chs_in_f[1][DATA][34] ), .Z(
        n468) );
  HS65_LS_AOI222X2 U98 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][34] ), 
        .C(n40), .D(\chs_in_f[0][DATA][34] ), .E(n56), .F(
        \chs_in_f[1][DATA][34] ), .Z(n433) );
  HS65_LS_AOI222X2 U99 ( .A(n72), .B(\chs_in_f[2][DATA][34] ), .C(n36), .D(
        \chs_in_f[0][DATA][34] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][34] ), .Z(n398) );
  HS65_LS_AOI222X2 U100 ( .A(n68), .B(\chs_in_f[2][DATA][34] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][34] ), .E(n52), .F(
        \chs_in_f[1][DATA][34] ), .Z(n363) );
  HS65_LS_OAI212X5 U101 ( .A(n300), .B(n21), .C(n335), .D(n6), .E(n406), .Z(
        \chs_out_f[2][DATA][0] ) );
  HS65_LS_AOI222X2 U102 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][0] ), 
        .C(n38), .D(\chs_in_f[0][DATA][0] ), .E(n54), .F(
        \chs_in_f[1][DATA][0] ), .Z(n406) );
  HS65_LS_OAI212X5 U103 ( .A(n299), .B(n21), .C(n334), .D(n6), .E(n417), .Z(
        \chs_out_f[2][DATA][1] ) );
  HS65_LS_AOI222X2 U104 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][1] ), 
        .C(n38), .D(\chs_in_f[0][DATA][1] ), .E(n54), .F(
        \chs_in_f[1][DATA][1] ), .Z(n417) );
  HS65_LS_OAI212X5 U105 ( .A(n298), .B(n22), .C(n333), .D(n7), .E(n428), .Z(
        \chs_out_f[2][DATA][2] ) );
  HS65_LS_AOI222X2 U106 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][2] ), 
        .C(n39), .D(\chs_in_f[0][DATA][2] ), .E(n55), .F(
        \chs_in_f[1][DATA][2] ), .Z(n428) );
  HS65_LS_OAI212X5 U107 ( .A(n290), .B(n21), .C(n325), .D(n6), .E(n407), .Z(
        \chs_out_f[2][DATA][10] ) );
  HS65_LS_AOI222X2 U108 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][10] ), 
        .C(n38), .D(\chs_in_f[0][DATA][10] ), .E(n54), .F(
        \chs_in_f[1][DATA][10] ), .Z(n407) );
  HS65_LS_OAI212X5 U109 ( .A(n289), .B(n21), .C(n324), .D(n6), .E(n408), .Z(
        \chs_out_f[2][DATA][11] ) );
  HS65_LS_AOI222X2 U110 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][11] ), 
        .C(n38), .D(\chs_in_f[0][DATA][11] ), .E(n54), .F(
        \chs_in_f[1][DATA][11] ), .Z(n408) );
  HS65_LS_OAI212X5 U111 ( .A(n288), .B(n21), .C(n323), .D(n6), .E(n409), .Z(
        \chs_out_f[2][DATA][12] ) );
  HS65_LS_AOI222X2 U112 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][12] ), 
        .C(n38), .D(\chs_in_f[0][DATA][12] ), .E(n54), .F(
        \chs_in_f[1][DATA][12] ), .Z(n409) );
  HS65_LS_OAI212X5 U113 ( .A(n287), .B(n21), .C(n322), .D(n6), .E(n410), .Z(
        \chs_out_f[2][DATA][13] ) );
  HS65_LS_AOI222X2 U114 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][13] ), 
        .C(n38), .D(\chs_in_f[0][DATA][13] ), .E(n54), .F(
        \chs_in_f[1][DATA][13] ), .Z(n410) );
  HS65_LS_OAI212X5 U115 ( .A(n286), .B(n21), .C(n321), .D(n6), .E(n411), .Z(
        \chs_out_f[2][DATA][14] ) );
  HS65_LS_AOI222X2 U116 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][14] ), 
        .C(n38), .D(\chs_in_f[0][DATA][14] ), .E(n54), .F(
        \chs_in_f[1][DATA][14] ), .Z(n411) );
  HS65_LS_OAI212X5 U117 ( .A(n285), .B(n21), .C(n320), .D(n6), .E(n412), .Z(
        \chs_out_f[2][DATA][15] ) );
  HS65_LS_AOI222X2 U118 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][15] ), 
        .C(n38), .D(\chs_in_f[0][DATA][15] ), .E(n54), .F(
        \chs_in_f[1][DATA][15] ), .Z(n412) );
  HS65_LS_OAI212X5 U119 ( .A(n284), .B(n21), .C(n319), .D(n6), .E(n413), .Z(
        \chs_out_f[2][DATA][16] ) );
  HS65_LS_AOI222X2 U120 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][16] ), 
        .C(n38), .D(\chs_in_f[0][DATA][16] ), .E(n54), .F(
        \chs_in_f[1][DATA][16] ), .Z(n413) );
  HS65_LS_OAI212X5 U121 ( .A(n283), .B(n21), .C(n318), .D(n6), .E(n414), .Z(
        \chs_out_f[2][DATA][17] ) );
  HS65_LS_AOI222X2 U122 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][17] ), 
        .C(n38), .D(\chs_in_f[0][DATA][17] ), .E(n54), .F(
        \chs_in_f[1][DATA][17] ), .Z(n414) );
  HS65_LS_OAI212X5 U123 ( .A(n282), .B(n21), .C(n317), .D(n6), .E(n415), .Z(
        \chs_out_f[2][DATA][18] ) );
  HS65_LS_AOI222X2 U124 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][18] ), 
        .C(n38), .D(\chs_in_f[0][DATA][18] ), .E(n54), .F(
        \chs_in_f[1][DATA][18] ), .Z(n415) );
  HS65_LS_OAI212X5 U125 ( .A(n281), .B(n21), .C(n316), .D(n6), .E(n416), .Z(
        \chs_out_f[2][DATA][19] ) );
  HS65_LS_AOI222X2 U126 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][19] ), 
        .C(n38), .D(\chs_in_f[0][DATA][19] ), .E(n54), .F(
        \chs_in_f[1][DATA][19] ), .Z(n416) );
  HS65_LS_OAI212X5 U127 ( .A(n280), .B(n21), .C(n315), .D(n7), .E(n418), .Z(
        \chs_out_f[2][DATA][20] ) );
  HS65_LS_AOI222X2 U128 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][20] ), 
        .C(n39), .D(\chs_in_f[0][DATA][20] ), .E(n55), .F(
        \chs_in_f[1][DATA][20] ), .Z(n418) );
  HS65_LS_OAI212X5 U129 ( .A(n279), .B(n22), .C(n314), .D(n7), .E(n419), .Z(
        \chs_out_f[2][DATA][21] ) );
  HS65_LS_AOI222X2 U130 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][21] ), 
        .C(n39), .D(\chs_in_f[0][DATA][21] ), .E(n55), .F(
        \chs_in_f[1][DATA][21] ), .Z(n419) );
  HS65_LS_OAI212X5 U131 ( .A(n278), .B(n22), .C(n313), .D(n7), .E(n420), .Z(
        \chs_out_f[2][DATA][22] ) );
  HS65_LS_AOI222X2 U132 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][22] ), 
        .C(n39), .D(\chs_in_f[0][DATA][22] ), .E(n55), .F(
        \chs_in_f[1][DATA][22] ), .Z(n420) );
  HS65_LS_OAI212X5 U133 ( .A(n277), .B(n22), .C(n312), .D(n7), .E(n421), .Z(
        \chs_out_f[2][DATA][23] ) );
  HS65_LS_AOI222X2 U134 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][23] ), 
        .C(n39), .D(\chs_in_f[0][DATA][23] ), .E(n55), .F(
        \chs_in_f[1][DATA][23] ), .Z(n421) );
  HS65_LS_OAI212X5 U135 ( .A(n276), .B(n22), .C(n311), .D(n7), .E(n422), .Z(
        \chs_out_f[2][DATA][24] ) );
  HS65_LS_AOI222X2 U136 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][24] ), 
        .C(n39), .D(\chs_in_f[0][DATA][24] ), .E(n55), .F(
        \chs_in_f[1][DATA][24] ), .Z(n422) );
  HS65_LS_OAI212X5 U137 ( .A(n275), .B(n22), .C(n310), .D(n7), .E(n423), .Z(
        \chs_out_f[2][DATA][25] ) );
  HS65_LS_AOI222X2 U138 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][25] ), 
        .C(n39), .D(\chs_in_f[0][DATA][25] ), .E(n55), .F(
        \chs_in_f[1][DATA][25] ), .Z(n423) );
  HS65_LS_OAI212X5 U139 ( .A(n274), .B(n22), .C(n309), .D(n7), .E(n424), .Z(
        \chs_out_f[2][DATA][26] ) );
  HS65_LS_AOI222X2 U140 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][26] ), 
        .C(n39), .D(\chs_in_f[0][DATA][26] ), .E(n55), .F(
        \chs_in_f[1][DATA][26] ), .Z(n424) );
  HS65_LS_OAI212X5 U141 ( .A(n273), .B(n22), .C(n308), .D(n7), .E(n425), .Z(
        \chs_out_f[2][DATA][27] ) );
  HS65_LS_AOI222X2 U142 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][27] ), 
        .C(n39), .D(\chs_in_f[0][DATA][27] ), .E(n55), .F(
        \chs_in_f[1][DATA][27] ), .Z(n425) );
  HS65_LS_OAI212X5 U143 ( .A(n272), .B(n22), .C(n307), .D(n7), .E(n426), .Z(
        \chs_out_f[2][DATA][28] ) );
  HS65_LS_AOI222X2 U144 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][28] ), 
        .C(n39), .D(\chs_in_f[0][DATA][28] ), .E(n55), .F(
        \chs_in_f[1][DATA][28] ), .Z(n426) );
  HS65_LS_OAI212X5 U145 ( .A(n271), .B(n22), .C(n306), .D(n7), .E(n427), .Z(
        \chs_out_f[2][DATA][29] ) );
  HS65_LS_AOI222X2 U146 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][29] ), 
        .C(n39), .D(\chs_in_f[0][DATA][29] ), .E(n55), .F(
        \chs_in_f[1][DATA][29] ), .Z(n427) );
  HS65_LS_OAI212X5 U147 ( .A(n270), .B(n22), .C(n305), .D(n7), .E(n429), .Z(
        \chs_out_f[2][DATA][30] ) );
  HS65_LS_AOI222X2 U148 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][30] ), 
        .C(n39), .D(\chs_in_f[0][DATA][30] ), .E(n55), .F(
        \chs_in_f[1][DATA][30] ), .Z(n429) );
  HS65_LS_OAI212X5 U149 ( .A(n300), .B(n24), .C(n335), .D(n9), .E(n371), .Z(
        \chs_out_f[1][DATA][0] ) );
  HS65_LS_AOI222X2 U150 ( .A(n70), .B(\chs_in_f[2][DATA][0] ), .C(n34), .D(
        \chs_in_f[0][DATA][0] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][0] ), .Z(n371) );
  HS65_LS_OAI212X5 U151 ( .A(n299), .B(n24), .C(n334), .D(n9), .E(n382), .Z(
        \chs_out_f[1][DATA][1] ) );
  HS65_LS_AOI222X2 U152 ( .A(n70), .B(\chs_in_f[2][DATA][1] ), .C(n34), .D(
        \chs_in_f[0][DATA][1] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][1] ), .Z(n382) );
  HS65_LS_OAI212X5 U153 ( .A(n298), .B(n25), .C(n333), .D(n10), .E(n393), .Z(
        \chs_out_f[1][DATA][2] ) );
  HS65_LS_AOI222X2 U154 ( .A(n71), .B(\chs_in_f[2][DATA][2] ), .C(n35), .D(
        \chs_in_f[0][DATA][2] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][2] ), .Z(n393) );
  HS65_LS_OAI212X5 U155 ( .A(n290), .B(n24), .C(n325), .D(n9), .E(n372), .Z(
        \chs_out_f[1][DATA][10] ) );
  HS65_LS_AOI222X2 U156 ( .A(n70), .B(\chs_in_f[2][DATA][10] ), .C(n34), .D(
        \chs_in_f[0][DATA][10] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][10] ), .Z(n372) );
  HS65_LS_OAI212X5 U157 ( .A(n289), .B(n24), .C(n324), .D(n9), .E(n373), .Z(
        \chs_out_f[1][DATA][11] ) );
  HS65_LS_AOI222X2 U158 ( .A(n70), .B(\chs_in_f[2][DATA][11] ), .C(n34), .D(
        \chs_in_f[0][DATA][11] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][11] ), .Z(n373) );
  HS65_LS_OAI212X5 U159 ( .A(n288), .B(n24), .C(n323), .D(n9), .E(n374), .Z(
        \chs_out_f[1][DATA][12] ) );
  HS65_LS_AOI222X2 U160 ( .A(n70), .B(\chs_in_f[2][DATA][12] ), .C(n34), .D(
        \chs_in_f[0][DATA][12] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][12] ), .Z(n374) );
  HS65_LS_OAI212X5 U161 ( .A(n287), .B(n24), .C(n322), .D(n9), .E(n375), .Z(
        \chs_out_f[1][DATA][13] ) );
  HS65_LS_AOI222X2 U162 ( .A(n70), .B(\chs_in_f[2][DATA][13] ), .C(n34), .D(
        \chs_in_f[0][DATA][13] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][13] ), .Z(n375) );
  HS65_LS_OAI212X5 U163 ( .A(n286), .B(n24), .C(n321), .D(n9), .E(n376), .Z(
        \chs_out_f[1][DATA][14] ) );
  HS65_LS_AOI222X2 U164 ( .A(n70), .B(\chs_in_f[2][DATA][14] ), .C(n34), .D(
        \chs_in_f[0][DATA][14] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][14] ), .Z(n376) );
  HS65_LS_OAI212X5 U165 ( .A(n285), .B(n24), .C(n320), .D(n9), .E(n377), .Z(
        \chs_out_f[1][DATA][15] ) );
  HS65_LS_AOI222X2 U166 ( .A(n70), .B(\chs_in_f[2][DATA][15] ), .C(n34), .D(
        \chs_in_f[0][DATA][15] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][15] ), .Z(n377) );
  HS65_LS_OAI212X5 U167 ( .A(n284), .B(n24), .C(n319), .D(n9), .E(n378), .Z(
        \chs_out_f[1][DATA][16] ) );
  HS65_LS_AOI222X2 U168 ( .A(n70), .B(\chs_in_f[2][DATA][16] ), .C(n34), .D(
        \chs_in_f[0][DATA][16] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][16] ), .Z(n378) );
  HS65_LS_OAI212X5 U169 ( .A(n283), .B(n24), .C(n318), .D(n9), .E(n379), .Z(
        \chs_out_f[1][DATA][17] ) );
  HS65_LS_AOI222X2 U170 ( .A(n70), .B(\chs_in_f[2][DATA][17] ), .C(n34), .D(
        \chs_in_f[0][DATA][17] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][17] ), .Z(n379) );
  HS65_LS_OAI212X5 U171 ( .A(n282), .B(n24), .C(n317), .D(n9), .E(n380), .Z(
        \chs_out_f[1][DATA][18] ) );
  HS65_LS_AOI222X2 U172 ( .A(n70), .B(\chs_in_f[2][DATA][18] ), .C(n34), .D(
        \chs_in_f[0][DATA][18] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][18] ), .Z(n380) );
  HS65_LS_OAI212X5 U173 ( .A(n281), .B(n24), .C(n316), .D(n9), .E(n381), .Z(
        \chs_out_f[1][DATA][19] ) );
  HS65_LS_AOI222X2 U174 ( .A(n70), .B(\chs_in_f[2][DATA][19] ), .C(n34), .D(
        \chs_in_f[0][DATA][19] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][19] ), .Z(n381) );
  HS65_LS_OAI212X5 U175 ( .A(n280), .B(n24), .C(n315), .D(n10), .E(n383), .Z(
        \chs_out_f[1][DATA][20] ) );
  HS65_LS_AOI222X2 U176 ( .A(n71), .B(\chs_in_f[2][DATA][20] ), .C(n35), .D(
        \chs_in_f[0][DATA][20] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][20] ), .Z(n383) );
  HS65_LS_OAI212X5 U177 ( .A(n279), .B(n25), .C(n314), .D(n10), .E(n384), .Z(
        \chs_out_f[1][DATA][21] ) );
  HS65_LS_AOI222X2 U178 ( .A(n71), .B(\chs_in_f[2][DATA][21] ), .C(n35), .D(
        \chs_in_f[0][DATA][21] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][21] ), .Z(n384) );
  HS65_LS_OAI212X5 U179 ( .A(n278), .B(n25), .C(n313), .D(n10), .E(n385), .Z(
        \chs_out_f[1][DATA][22] ) );
  HS65_LS_AOI222X2 U180 ( .A(n71), .B(\chs_in_f[2][DATA][22] ), .C(n35), .D(
        \chs_in_f[0][DATA][22] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][22] ), .Z(n385) );
  HS65_LS_OAI212X5 U181 ( .A(n277), .B(n25), .C(n312), .D(n10), .E(n386), .Z(
        \chs_out_f[1][DATA][23] ) );
  HS65_LS_AOI222X2 U182 ( .A(n71), .B(\chs_in_f[2][DATA][23] ), .C(n35), .D(
        \chs_in_f[0][DATA][23] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][23] ), .Z(n386) );
  HS65_LS_OAI212X5 U183 ( .A(n276), .B(n25), .C(n311), .D(n10), .E(n387), .Z(
        \chs_out_f[1][DATA][24] ) );
  HS65_LS_AOI222X2 U184 ( .A(n71), .B(\chs_in_f[2][DATA][24] ), .C(n35), .D(
        \chs_in_f[0][DATA][24] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][24] ), .Z(n387) );
  HS65_LS_OAI212X5 U185 ( .A(n275), .B(n25), .C(n310), .D(n10), .E(n388), .Z(
        \chs_out_f[1][DATA][25] ) );
  HS65_LS_AOI222X2 U186 ( .A(n71), .B(\chs_in_f[2][DATA][25] ), .C(n35), .D(
        \chs_in_f[0][DATA][25] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][25] ), .Z(n388) );
  HS65_LS_OAI212X5 U187 ( .A(n274), .B(n25), .C(n309), .D(n10), .E(n389), .Z(
        \chs_out_f[1][DATA][26] ) );
  HS65_LS_AOI222X2 U188 ( .A(n71), .B(\chs_in_f[2][DATA][26] ), .C(n35), .D(
        \chs_in_f[0][DATA][26] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][26] ), .Z(n389) );
  HS65_LS_OAI212X5 U189 ( .A(n273), .B(n25), .C(n308), .D(n10), .E(n390), .Z(
        \chs_out_f[1][DATA][27] ) );
  HS65_LS_AOI222X2 U190 ( .A(n71), .B(\chs_in_f[2][DATA][27] ), .C(n35), .D(
        \chs_in_f[0][DATA][27] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][27] ), .Z(n390) );
  HS65_LS_OAI212X5 U191 ( .A(n272), .B(n25), .C(n307), .D(n10), .E(n391), .Z(
        \chs_out_f[1][DATA][28] ) );
  HS65_LS_AOI222X2 U192 ( .A(n71), .B(\chs_in_f[2][DATA][28] ), .C(n35), .D(
        \chs_in_f[0][DATA][28] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][28] ), .Z(n391) );
  HS65_LS_OAI212X5 U193 ( .A(n271), .B(n25), .C(n306), .D(n10), .E(n392), .Z(
        \chs_out_f[1][DATA][29] ) );
  HS65_LS_AOI222X2 U194 ( .A(n71), .B(\chs_in_f[2][DATA][29] ), .C(n35), .D(
        \chs_in_f[0][DATA][29] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][29] ), .Z(n392) );
  HS65_LS_OAI212X5 U195 ( .A(n270), .B(n25), .C(n305), .D(n10), .E(n394), .Z(
        \chs_out_f[1][DATA][30] ) );
  HS65_LS_AOI222X2 U196 ( .A(n71), .B(\chs_in_f[2][DATA][30] ), .C(n35), .D(
        \chs_in_f[0][DATA][30] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][30] ), .Z(n394) );
  HS65_LS_IVX9 U197 ( .A(\chs_in_f[3][DATA][9] ), .Z(n291) );
  HS65_LS_IVX9 U198 ( .A(\chs_in_f[3][DATA][34] ), .Z(n266) );
  HS65_LS_IVX9 U199 ( .A(\chs_in_f[3][DATA][0] ), .Z(n300) );
  HS65_LS_IVX9 U200 ( .A(\chs_in_f[3][DATA][1] ), .Z(n299) );
  HS65_LS_IVX9 U201 ( .A(\chs_in_f[3][DATA][2] ), .Z(n298) );
  HS65_LS_IVX9 U202 ( .A(\chs_in_f[3][DATA][3] ), .Z(n297) );
  HS65_LS_IVX9 U203 ( .A(\chs_in_f[3][DATA][4] ), .Z(n296) );
  HS65_LS_IVX9 U204 ( .A(\chs_in_f[3][DATA][5] ), .Z(n295) );
  HS65_LS_IVX9 U205 ( .A(\chs_in_f[3][DATA][6] ), .Z(n294) );
  HS65_LS_IVX9 U206 ( .A(\chs_in_f[3][DATA][7] ), .Z(n293) );
  HS65_LS_IVX9 U207 ( .A(\chs_in_f[3][DATA][8] ), .Z(n292) );
  HS65_LS_IVX9 U208 ( .A(\chs_in_f[3][DATA][10] ), .Z(n290) );
  HS65_LS_IVX9 U209 ( .A(\chs_in_f[3][DATA][11] ), .Z(n289) );
  HS65_LS_IVX9 U210 ( .A(\chs_in_f[3][DATA][12] ), .Z(n288) );
  HS65_LS_IVX9 U211 ( .A(\chs_in_f[3][DATA][13] ), .Z(n287) );
  HS65_LS_IVX9 U212 ( .A(\chs_in_f[3][DATA][14] ), .Z(n286) );
  HS65_LS_IVX9 U213 ( .A(\chs_in_f[3][DATA][15] ), .Z(n285) );
  HS65_LS_IVX9 U214 ( .A(\chs_in_f[3][DATA][16] ), .Z(n284) );
  HS65_LS_IVX9 U215 ( .A(\chs_in_f[3][DATA][17] ), .Z(n283) );
  HS65_LS_IVX9 U216 ( .A(\chs_in_f[3][DATA][18] ), .Z(n282) );
  HS65_LS_IVX9 U217 ( .A(\chs_in_f[3][DATA][19] ), .Z(n281) );
  HS65_LS_IVX9 U218 ( .A(\chs_in_f[3][DATA][20] ), .Z(n280) );
  HS65_LS_IVX9 U219 ( .A(\chs_in_f[3][DATA][21] ), .Z(n279) );
  HS65_LS_IVX9 U220 ( .A(\chs_in_f[3][DATA][22] ), .Z(n278) );
  HS65_LS_IVX9 U221 ( .A(\chs_in_f[3][DATA][23] ), .Z(n277) );
  HS65_LS_IVX9 U222 ( .A(\chs_in_f[3][DATA][24] ), .Z(n276) );
  HS65_LS_IVX9 U223 ( .A(\chs_in_f[3][DATA][25] ), .Z(n275) );
  HS65_LS_IVX9 U224 ( .A(\chs_in_f[3][DATA][26] ), .Z(n274) );
  HS65_LS_IVX9 U225 ( .A(\chs_in_f[3][DATA][27] ), .Z(n273) );
  HS65_LS_IVX9 U226 ( .A(\chs_in_f[3][DATA][28] ), .Z(n272) );
  HS65_LS_IVX9 U227 ( .A(\chs_in_f[3][DATA][29] ), .Z(n271) );
  HS65_LS_IVX9 U228 ( .A(\chs_in_f[3][DATA][30] ), .Z(n270) );
  HS65_LS_IVX9 U229 ( .A(\chs_in_f[3][DATA][31] ), .Z(n269) );
  HS65_LS_IVX9 U230 ( .A(\chs_in_f[3][DATA][32] ), .Z(n268) );
  HS65_LS_IVX9 U231 ( .A(\chs_in_f[3][DATA][33] ), .Z(n267) );
  HS65_LS_IVX9 U232 ( .A(\chs_in_f[4][DATA][9] ), .Z(n326) );
  HS65_LS_IVX9 U233 ( .A(\chs_in_f[4][DATA][34] ), .Z(n301) );
  HS65_LS_IVX9 U234 ( .A(\chs_in_f[4][DATA][0] ), .Z(n335) );
  HS65_LS_IVX9 U235 ( .A(\chs_in_f[4][DATA][1] ), .Z(n334) );
  HS65_LS_IVX9 U236 ( .A(\chs_in_f[4][DATA][2] ), .Z(n333) );
  HS65_LS_IVX9 U237 ( .A(\chs_in_f[4][DATA][3] ), .Z(n332) );
  HS65_LS_IVX9 U238 ( .A(\chs_in_f[4][DATA][4] ), .Z(n331) );
  HS65_LS_IVX9 U239 ( .A(\chs_in_f[4][DATA][5] ), .Z(n330) );
  HS65_LS_IVX9 U240 ( .A(\chs_in_f[4][DATA][6] ), .Z(n329) );
  HS65_LS_IVX9 U241 ( .A(\chs_in_f[4][DATA][7] ), .Z(n328) );
  HS65_LS_IVX9 U242 ( .A(\chs_in_f[4][DATA][8] ), .Z(n327) );
  HS65_LS_IVX9 U243 ( .A(\chs_in_f[4][DATA][10] ), .Z(n325) );
  HS65_LS_IVX9 U244 ( .A(\chs_in_f[4][DATA][11] ), .Z(n324) );
  HS65_LS_IVX9 U245 ( .A(\chs_in_f[4][DATA][12] ), .Z(n323) );
  HS65_LS_IVX9 U246 ( .A(\chs_in_f[4][DATA][13] ), .Z(n322) );
  HS65_LS_IVX9 U247 ( .A(\chs_in_f[4][DATA][14] ), .Z(n321) );
  HS65_LS_IVX9 U248 ( .A(\chs_in_f[4][DATA][15] ), .Z(n320) );
  HS65_LS_IVX9 U249 ( .A(\chs_in_f[4][DATA][16] ), .Z(n319) );
  HS65_LS_IVX9 U250 ( .A(\chs_in_f[4][DATA][17] ), .Z(n318) );
  HS65_LS_IVX9 U251 ( .A(\chs_in_f[4][DATA][18] ), .Z(n317) );
  HS65_LS_IVX9 U252 ( .A(\chs_in_f[4][DATA][19] ), .Z(n316) );
  HS65_LS_IVX9 U253 ( .A(\chs_in_f[4][DATA][20] ), .Z(n315) );
  HS65_LS_IVX9 U254 ( .A(\chs_in_f[4][DATA][21] ), .Z(n314) );
  HS65_LS_IVX9 U255 ( .A(\chs_in_f[4][DATA][22] ), .Z(n313) );
  HS65_LS_IVX9 U256 ( .A(\chs_in_f[4][DATA][23] ), .Z(n312) );
  HS65_LS_IVX9 U257 ( .A(\chs_in_f[4][DATA][24] ), .Z(n311) );
  HS65_LS_IVX9 U258 ( .A(\chs_in_f[4][DATA][25] ), .Z(n310) );
  HS65_LS_IVX9 U259 ( .A(\chs_in_f[4][DATA][26] ), .Z(n309) );
  HS65_LS_IVX9 U260 ( .A(\chs_in_f[4][DATA][27] ), .Z(n308) );
  HS65_LS_IVX9 U261 ( .A(\chs_in_f[4][DATA][28] ), .Z(n307) );
  HS65_LS_IVX9 U262 ( .A(\chs_in_f[4][DATA][29] ), .Z(n306) );
  HS65_LS_IVX9 U263 ( .A(\chs_in_f[4][DATA][30] ), .Z(n305) );
  HS65_LS_IVX9 U264 ( .A(\chs_in_f[4][DATA][31] ), .Z(n304) );
  HS65_LS_IVX9 U265 ( .A(\chs_in_f[4][DATA][32] ), .Z(n303) );
  HS65_LS_IVX9 U266 ( .A(\chs_in_f[4][DATA][33] ), .Z(n302) );
  HS65_LS_BFX18 U267 ( .A(\switch_sel[2][4] ), .Z(n77) );
  HS65_LS_BFX18 U268 ( .A(\switch_sel[2][3] ), .Z(n73) );
  HS65_LS_BFX18 U269 ( .A(\switch_sel[0][2] ), .Z(n37) );
  HS65_LS_BFX18 U270 ( .A(\switch_sel[2][1] ), .Z(n69) );
  HS65_LS_BFX18 U271 ( .A(\switch_sel[2][0] ), .Z(n65) );
  HS65_LS_AOI222X2 U272 ( .A(\chs_in_f[2][DATA][0] ), .B(n80), .C(
        \chs_in_f[0][DATA][0] ), .D(n46), .E(\chs_in_f[1][DATA][0] ), .F(n64), 
        .Z(n476) );
  HS65_LS_AOI222X2 U273 ( .A(\chs_in_f[2][DATA][1] ), .B(n79), .C(
        \chs_in_f[0][DATA][1] ), .D(n46), .E(\chs_in_f[1][DATA][1] ), .F(n63), 
        .Z(n487) );
  HS65_LS_AOI222X2 U274 ( .A(\chs_in_f[2][DATA][2] ), .B(n78), .C(
        \chs_in_f[0][DATA][2] ), .D(n47), .E(\chs_in_f[1][DATA][2] ), .F(n62), 
        .Z(n498) );
  HS65_LS_AOI222X2 U275 ( .A(\chs_in_f[2][DATA][3] ), .B(n78), .C(
        \chs_in_f[0][DATA][3] ), .D(n48), .E(\chs_in_f[1][DATA][3] ), .F(n62), 
        .Z(n504) );
  HS65_LS_AOI222X2 U276 ( .A(\chs_in_f[2][DATA][4] ), .B(n78), .C(
        \chs_in_f[0][DATA][4] ), .D(n48), .E(\chs_in_f[1][DATA][4] ), .F(n62), 
        .Z(n505) );
  HS65_LS_OAI212X5 U277 ( .A(n20), .B(n295), .C(n17), .D(n330), .E(n506), .Z(
        \chs_out_f[4][DATA][5] ) );
  HS65_LS_AOI222X2 U278 ( .A(\chs_in_f[2][DATA][5] ), .B(n78), .C(
        \chs_in_f[0][DATA][5] ), .D(n48), .E(\chs_in_f[1][DATA][5] ), .F(n62), 
        .Z(n506) );
  HS65_LS_OAI212X5 U279 ( .A(n20), .B(n294), .C(n17), .D(n329), .E(n507), .Z(
        \chs_out_f[4][DATA][6] ) );
  HS65_LS_AOI222X2 U280 ( .A(\chs_in_f[2][DATA][6] ), .B(n78), .C(
        \chs_in_f[0][DATA][6] ), .D(n48), .E(\chs_in_f[1][DATA][6] ), .F(n62), 
        .Z(n507) );
  HS65_LS_OAI212X5 U281 ( .A(n20), .B(n293), .C(n17), .D(n328), .E(n508), .Z(
        \chs_out_f[4][DATA][7] ) );
  HS65_LS_AOI222X2 U282 ( .A(\chs_in_f[2][DATA][7] ), .B(n78), .C(
        \chs_in_f[0][DATA][7] ), .D(n48), .E(\chs_in_f[1][DATA][7] ), .F(n62), 
        .Z(n508) );
  HS65_LS_OAI212X5 U283 ( .A(n20), .B(n292), .C(n17), .D(n327), .E(n509), .Z(
        \chs_out_f[4][DATA][8] ) );
  HS65_LS_AOI222X2 U284 ( .A(\chs_in_f[2][DATA][8] ), .B(n78), .C(
        \chs_in_f[0][DATA][8] ), .D(n48), .E(\chs_in_f[1][DATA][8] ), .F(n62), 
        .Z(n509) );
  HS65_LS_AOI222X2 U285 ( .A(\chs_in_f[2][DATA][10] ), .B(n80), .C(
        \chs_in_f[0][DATA][10] ), .D(n46), .E(\chs_in_f[1][DATA][10] ), .F(n64), .Z(n477) );
  HS65_LS_AOI222X2 U286 ( .A(\chs_in_f[2][DATA][11] ), .B(n80), .C(
        \chs_in_f[0][DATA][11] ), .D(n46), .E(\chs_in_f[1][DATA][11] ), .F(n64), .Z(n478) );
  HS65_LS_AOI222X2 U287 ( .A(\chs_in_f[2][DATA][12] ), .B(n80), .C(
        \chs_in_f[0][DATA][12] ), .D(n46), .E(\chs_in_f[1][DATA][12] ), .F(n64), .Z(n479) );
  HS65_LS_AOI222X2 U288 ( .A(\chs_in_f[2][DATA][13] ), .B(n80), .C(
        \chs_in_f[0][DATA][13] ), .D(n46), .E(\chs_in_f[1][DATA][13] ), .F(n64), .Z(n480) );
  HS65_LS_OAI212X5 U289 ( .A(n18), .B(n286), .C(n15), .D(n321), .E(n481), .Z(
        \chs_out_f[4][DATA][14] ) );
  HS65_LS_AOI222X2 U290 ( .A(\chs_in_f[2][DATA][14] ), .B(n80), .C(
        \chs_in_f[0][DATA][14] ), .D(n46), .E(\chs_in_f[1][DATA][14] ), .F(n64), .Z(n481) );
  HS65_LS_OAI212X5 U291 ( .A(n18), .B(n285), .C(n15), .D(n320), .E(n482), .Z(
        \chs_out_f[4][DATA][15] ) );
  HS65_LS_AOI222X2 U292 ( .A(\chs_in_f[2][DATA][15] ), .B(n80), .C(
        \chs_in_f[0][DATA][15] ), .D(n46), .E(\chs_in_f[1][DATA][15] ), .F(n64), .Z(n482) );
  HS65_LS_OAI212X5 U293 ( .A(n18), .B(n284), .C(n15), .D(n319), .E(n483), .Z(
        \chs_out_f[4][DATA][16] ) );
  HS65_LS_AOI222X2 U294 ( .A(\chs_in_f[2][DATA][16] ), .B(n80), .C(
        \chs_in_f[0][DATA][16] ), .D(n46), .E(\chs_in_f[1][DATA][16] ), .F(n64), .Z(n483) );
  HS65_LS_OAI212X5 U295 ( .A(n18), .B(n283), .C(n15), .D(n318), .E(n484), .Z(
        \chs_out_f[4][DATA][17] ) );
  HS65_LS_AOI222X2 U296 ( .A(\chs_in_f[2][DATA][17] ), .B(n80), .C(
        \chs_in_f[0][DATA][17] ), .D(n46), .E(\chs_in_f[1][DATA][17] ), .F(n64), .Z(n484) );
  HS65_LS_OAI212X5 U297 ( .A(n18), .B(n282), .C(n15), .D(n317), .E(n485), .Z(
        \chs_out_f[4][DATA][18] ) );
  HS65_LS_AOI222X2 U298 ( .A(\chs_in_f[2][DATA][18] ), .B(n79), .C(
        \chs_in_f[0][DATA][18] ), .D(n46), .E(\chs_in_f[1][DATA][18] ), .F(n63), .Z(n485) );
  HS65_LS_OAI212X5 U299 ( .A(n18), .B(n281), .C(n15), .D(n316), .E(n486), .Z(
        \chs_out_f[4][DATA][19] ) );
  HS65_LS_AOI222X2 U300 ( .A(\chs_in_f[2][DATA][19] ), .B(n79), .C(
        \chs_in_f[0][DATA][19] ), .D(n46), .E(\chs_in_f[1][DATA][19] ), .F(n63), .Z(n486) );
  HS65_LS_OAI212X5 U301 ( .A(n19), .B(n280), .C(n15), .D(n315), .E(n488), .Z(
        \chs_out_f[4][DATA][20] ) );
  HS65_LS_AOI222X2 U302 ( .A(\chs_in_f[2][DATA][20] ), .B(n79), .C(
        \chs_in_f[0][DATA][20] ), .D(n47), .E(\chs_in_f[1][DATA][20] ), .F(n63), .Z(n488) );
  HS65_LS_OAI212X5 U303 ( .A(n19), .B(n279), .C(n16), .D(n314), .E(n489), .Z(
        \chs_out_f[4][DATA][21] ) );
  HS65_LS_AOI222X2 U304 ( .A(\chs_in_f[2][DATA][21] ), .B(n79), .C(
        \chs_in_f[0][DATA][21] ), .D(n47), .E(\chs_in_f[1][DATA][21] ), .F(n63), .Z(n489) );
  HS65_LS_OAI212X5 U305 ( .A(n19), .B(n278), .C(n16), .D(n313), .E(n490), .Z(
        \chs_out_f[4][DATA][22] ) );
  HS65_LS_AOI222X2 U306 ( .A(\chs_in_f[2][DATA][22] ), .B(n79), .C(
        \chs_in_f[0][DATA][22] ), .D(n47), .E(\chs_in_f[1][DATA][22] ), .F(n63), .Z(n490) );
  HS65_LS_OAI212X5 U307 ( .A(n19), .B(n277), .C(n16), .D(n312), .E(n491), .Z(
        \chs_out_f[4][DATA][23] ) );
  HS65_LS_AOI222X2 U308 ( .A(\chs_in_f[2][DATA][23] ), .B(n79), .C(
        \chs_in_f[0][DATA][23] ), .D(n47), .E(\chs_in_f[1][DATA][23] ), .F(n63), .Z(n491) );
  HS65_LS_OAI212X5 U309 ( .A(n19), .B(n276), .C(n16), .D(n311), .E(n492), .Z(
        \chs_out_f[4][DATA][24] ) );
  HS65_LS_AOI222X2 U310 ( .A(\chs_in_f[2][DATA][24] ), .B(n79), .C(
        \chs_in_f[0][DATA][24] ), .D(n47), .E(\chs_in_f[1][DATA][24] ), .F(n63), .Z(n492) );
  HS65_LS_OAI212X5 U311 ( .A(n19), .B(n275), .C(n16), .D(n310), .E(n493), .Z(
        \chs_out_f[4][DATA][25] ) );
  HS65_LS_AOI222X2 U312 ( .A(\chs_in_f[2][DATA][25] ), .B(n79), .C(
        \chs_in_f[0][DATA][25] ), .D(n47), .E(\chs_in_f[1][DATA][25] ), .F(n63), .Z(n493) );
  HS65_LS_OAI212X5 U313 ( .A(n19), .B(n274), .C(n16), .D(n309), .E(n494), .Z(
        \chs_out_f[4][DATA][26] ) );
  HS65_LS_AOI222X2 U314 ( .A(\chs_in_f[2][DATA][26] ), .B(n79), .C(
        \chs_in_f[0][DATA][26] ), .D(n47), .E(\chs_in_f[1][DATA][26] ), .F(n63), .Z(n494) );
  HS65_LS_OAI212X5 U315 ( .A(n19), .B(n273), .C(n16), .D(n308), .E(n495), .Z(
        \chs_out_f[4][DATA][27] ) );
  HS65_LS_AOI222X2 U316 ( .A(\chs_in_f[2][DATA][27] ), .B(n79), .C(
        \chs_in_f[0][DATA][27] ), .D(n47), .E(\chs_in_f[1][DATA][27] ), .F(n63), .Z(n495) );
  HS65_LS_OAI212X5 U317 ( .A(n19), .B(n272), .C(n16), .D(n307), .E(n496), .Z(
        \chs_out_f[4][DATA][28] ) );
  HS65_LS_AOI222X2 U318 ( .A(\chs_in_f[2][DATA][28] ), .B(n79), .C(
        \chs_in_f[0][DATA][28] ), .D(n47), .E(\chs_in_f[1][DATA][28] ), .F(n63), .Z(n496) );
  HS65_LS_OAI212X5 U319 ( .A(n19), .B(n271), .C(n16), .D(n306), .E(n497), .Z(
        \chs_out_f[4][DATA][29] ) );
  HS65_LS_AOI222X2 U320 ( .A(\chs_in_f[2][DATA][29] ), .B(n79), .C(
        \chs_in_f[0][DATA][29] ), .D(n47), .E(\chs_in_f[1][DATA][29] ), .F(n63), .Z(n497) );
  HS65_LS_OAI212X5 U321 ( .A(n19), .B(n270), .C(n16), .D(n305), .E(n499), .Z(
        \chs_out_f[4][DATA][30] ) );
  HS65_LS_AOI222X2 U322 ( .A(\chs_in_f[2][DATA][30] ), .B(n78), .C(
        \chs_in_f[0][DATA][30] ), .D(n47), .E(\chs_in_f[1][DATA][30] ), .F(n62), .Z(n499) );
  HS65_LS_OAI212X5 U323 ( .A(n20), .B(n269), .C(n16), .D(n304), .E(n500), .Z(
        \chs_out_f[4][DATA][31] ) );
  HS65_LS_AOI222X2 U324 ( .A(\chs_in_f[2][DATA][31] ), .B(n78), .C(
        \chs_in_f[0][DATA][31] ), .D(n48), .E(\chs_in_f[1][DATA][31] ), .F(n62), .Z(n500) );
  HS65_LS_OAI212X5 U325 ( .A(n20), .B(n268), .C(n16), .D(n303), .E(n501), .Z(
        \chs_out_f[4][DATA][32] ) );
  HS65_LS_AOI222X2 U326 ( .A(\chs_in_f[2][DATA][32] ), .B(n78), .C(
        \chs_in_f[0][DATA][32] ), .D(n48), .E(\chs_in_f[1][DATA][32] ), .F(n62), .Z(n501) );
  HS65_LS_OAI212X5 U327 ( .A(n20), .B(n267), .C(n17), .D(n302), .E(n502), .Z(
        \chs_out_f[4][DATA][33] ) );
  HS65_LS_AOI222X2 U328 ( .A(\chs_in_f[2][DATA][33] ), .B(n78), .C(
        \chs_in_f[0][DATA][33] ), .D(n48), .E(\chs_in_f[1][DATA][33] ), .F(n62), .Z(n502) );
  HS65_LS_OAI212X5 U329 ( .A(n291), .B(n23), .C(n326), .D(n8), .E(n440), .Z(
        \chs_out_f[2][DATA][9] ) );
  HS65_LS_AOI222X2 U330 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][9] ), 
        .C(n40), .D(\chs_in_f[0][DATA][9] ), .E(n56), .F(
        \chs_in_f[1][DATA][9] ), .Z(n440) );
  HS65_LS_OAI212X5 U331 ( .A(n291), .B(n26), .C(n326), .D(n11), .E(n405), .Z(
        \chs_out_f[1][DATA][9] ) );
  HS65_LS_AOI222X2 U332 ( .A(n72), .B(\chs_in_f[2][DATA][9] ), .C(n36), .D(
        \chs_in_f[0][DATA][9] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][9] ), .Z(n405) );
  HS65_LS_OAI212X5 U333 ( .A(n291), .B(n29), .C(n326), .D(n14), .E(n370), .Z(
        \chs_out_f[0][DATA][9] ) );
  HS65_LS_AOI222X2 U334 ( .A(n68), .B(\chs_in_f[2][DATA][9] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][9] ), .E(n52), .F(
        \chs_in_f[1][DATA][9] ), .Z(n370) );
  HS65_LS_OAI212X5 U335 ( .A(n269), .B(n22), .C(n304), .D(n8), .E(n430), .Z(
        \chs_out_f[2][DATA][31] ) );
  HS65_LS_AOI222X2 U336 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][31] ), 
        .C(n40), .D(\chs_in_f[0][DATA][31] ), .E(n56), .F(
        \chs_in_f[1][DATA][31] ), .Z(n430) );
  HS65_LS_OAI212X5 U337 ( .A(n268), .B(n22), .C(n303), .D(n8), .E(n431), .Z(
        \chs_out_f[2][DATA][32] ) );
  HS65_LS_AOI222X2 U338 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][32] ), 
        .C(n40), .D(\chs_in_f[0][DATA][32] ), .E(n56), .F(
        \chs_in_f[1][DATA][32] ), .Z(n431) );
  HS65_LS_OAI212X5 U339 ( .A(n269), .B(n25), .C(n304), .D(n11), .E(n395), .Z(
        \chs_out_f[1][DATA][31] ) );
  HS65_LS_AOI222X2 U340 ( .A(n72), .B(\chs_in_f[2][DATA][31] ), .C(n36), .D(
        \chs_in_f[0][DATA][31] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][31] ), .Z(n395) );
  HS65_LS_OAI212X5 U341 ( .A(n268), .B(n25), .C(n303), .D(n11), .E(n396), .Z(
        \chs_out_f[1][DATA][32] ) );
  HS65_LS_AOI222X2 U342 ( .A(n72), .B(\chs_in_f[2][DATA][32] ), .C(n36), .D(
        \chs_in_f[0][DATA][32] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][32] ), .Z(n396) );
  HS65_LS_OAI212X5 U343 ( .A(n300), .B(n27), .C(n335), .D(n12), .E(n336), .Z(
        \chs_out_f[0][DATA][0] ) );
  HS65_LS_AOI222X2 U344 ( .A(n66), .B(\chs_in_f[2][DATA][0] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][0] ), .E(n50), .F(
        \chs_in_f[1][DATA][0] ), .Z(n336) );
  HS65_LS_OAI212X5 U345 ( .A(n299), .B(n27), .C(n334), .D(n12), .E(n347), .Z(
        \chs_out_f[0][DATA][1] ) );
  HS65_LS_AOI222X2 U346 ( .A(n66), .B(\chs_in_f[2][DATA][1] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][1] ), .E(n50), .F(
        \chs_in_f[1][DATA][1] ), .Z(n347) );
  HS65_LS_OAI212X5 U347 ( .A(n298), .B(n28), .C(n333), .D(n13), .E(n358), .Z(
        \chs_out_f[0][DATA][2] ) );
  HS65_LS_AOI222X2 U348 ( .A(n67), .B(\chs_in_f[2][DATA][2] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][2] ), .E(n51), .F(
        \chs_in_f[1][DATA][2] ), .Z(n358) );
  HS65_LS_OAI212X5 U349 ( .A(n290), .B(n27), .C(n325), .D(n12), .E(n337), .Z(
        \chs_out_f[0][DATA][10] ) );
  HS65_LS_AOI222X2 U350 ( .A(n66), .B(\chs_in_f[2][DATA][10] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][10] ), .E(n50), .F(
        \chs_in_f[1][DATA][10] ), .Z(n337) );
  HS65_LS_OAI212X5 U351 ( .A(n289), .B(n27), .C(n324), .D(n12), .E(n338), .Z(
        \chs_out_f[0][DATA][11] ) );
  HS65_LS_AOI222X2 U352 ( .A(n66), .B(\chs_in_f[2][DATA][11] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][11] ), .E(n50), .F(
        \chs_in_f[1][DATA][11] ), .Z(n338) );
  HS65_LS_OAI212X5 U353 ( .A(n288), .B(n27), .C(n323), .D(n12), .E(n339), .Z(
        \chs_out_f[0][DATA][12] ) );
  HS65_LS_AOI222X2 U354 ( .A(n66), .B(\chs_in_f[2][DATA][12] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][12] ), .E(n50), .F(
        \chs_in_f[1][DATA][12] ), .Z(n339) );
  HS65_LS_OAI212X5 U355 ( .A(n287), .B(n27), .C(n322), .D(n12), .E(n340), .Z(
        \chs_out_f[0][DATA][13] ) );
  HS65_LS_AOI222X2 U356 ( .A(n66), .B(\chs_in_f[2][DATA][13] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][13] ), .E(n50), .F(
        \chs_in_f[1][DATA][13] ), .Z(n340) );
  HS65_LS_OAI212X5 U357 ( .A(n286), .B(n27), .C(n321), .D(n12), .E(n341), .Z(
        \chs_out_f[0][DATA][14] ) );
  HS65_LS_AOI222X2 U358 ( .A(n66), .B(\chs_in_f[2][DATA][14] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][14] ), .E(n50), .F(
        \chs_in_f[1][DATA][14] ), .Z(n341) );
  HS65_LS_OAI212X5 U359 ( .A(n285), .B(n27), .C(n320), .D(n12), .E(n342), .Z(
        \chs_out_f[0][DATA][15] ) );
  HS65_LS_AOI222X2 U360 ( .A(n66), .B(\chs_in_f[2][DATA][15] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][15] ), .E(n50), .F(
        \chs_in_f[1][DATA][15] ), .Z(n342) );
  HS65_LS_OAI212X5 U361 ( .A(n284), .B(n27), .C(n319), .D(n12), .E(n343), .Z(
        \chs_out_f[0][DATA][16] ) );
  HS65_LS_AOI222X2 U362 ( .A(n66), .B(\chs_in_f[2][DATA][16] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][16] ), .E(n50), .F(
        \chs_in_f[1][DATA][16] ), .Z(n343) );
  HS65_LS_OAI212X5 U363 ( .A(n283), .B(n27), .C(n318), .D(n12), .E(n344), .Z(
        \chs_out_f[0][DATA][17] ) );
  HS65_LS_AOI222X2 U364 ( .A(n66), .B(\chs_in_f[2][DATA][17] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][17] ), .E(n50), .F(
        \chs_in_f[1][DATA][17] ), .Z(n344) );
  HS65_LS_OAI212X5 U365 ( .A(n282), .B(n27), .C(n317), .D(n12), .E(n345), .Z(
        \chs_out_f[0][DATA][18] ) );
  HS65_LS_AOI222X2 U366 ( .A(n66), .B(\chs_in_f[2][DATA][18] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][18] ), .E(n50), .F(
        \chs_in_f[1][DATA][18] ), .Z(n345) );
  HS65_LS_OAI212X5 U367 ( .A(n281), .B(n27), .C(n316), .D(n12), .E(n346), .Z(
        \chs_out_f[0][DATA][19] ) );
  HS65_LS_AOI222X2 U368 ( .A(n66), .B(\chs_in_f[2][DATA][19] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][19] ), .E(n50), .F(
        \chs_in_f[1][DATA][19] ), .Z(n346) );
  HS65_LS_OAI212X5 U369 ( .A(n280), .B(n27), .C(n315), .D(n13), .E(n348), .Z(
        \chs_out_f[0][DATA][20] ) );
  HS65_LS_AOI222X2 U370 ( .A(n67), .B(\chs_in_f[2][DATA][20] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][20] ), .E(n51), .F(
        \chs_in_f[1][DATA][20] ), .Z(n348) );
  HS65_LS_OAI212X5 U371 ( .A(n279), .B(n28), .C(n314), .D(n13), .E(n349), .Z(
        \chs_out_f[0][DATA][21] ) );
  HS65_LS_AOI222X2 U372 ( .A(n67), .B(\chs_in_f[2][DATA][21] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][21] ), .E(n51), .F(
        \chs_in_f[1][DATA][21] ), .Z(n349) );
  HS65_LS_OAI212X5 U373 ( .A(n278), .B(n28), .C(n313), .D(n13), .E(n350), .Z(
        \chs_out_f[0][DATA][22] ) );
  HS65_LS_AOI222X2 U374 ( .A(n67), .B(\chs_in_f[2][DATA][22] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][22] ), .E(n51), .F(
        \chs_in_f[1][DATA][22] ), .Z(n350) );
  HS65_LS_OAI212X5 U375 ( .A(n277), .B(n28), .C(n312), .D(n13), .E(n351), .Z(
        \chs_out_f[0][DATA][23] ) );
  HS65_LS_AOI222X2 U376 ( .A(n67), .B(\chs_in_f[2][DATA][23] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][23] ), .E(n51), .F(
        \chs_in_f[1][DATA][23] ), .Z(n351) );
  HS65_LS_OAI212X5 U377 ( .A(n276), .B(n28), .C(n311), .D(n13), .E(n352), .Z(
        \chs_out_f[0][DATA][24] ) );
  HS65_LS_AOI222X2 U378 ( .A(n67), .B(\chs_in_f[2][DATA][24] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][24] ), .E(n51), .F(
        \chs_in_f[1][DATA][24] ), .Z(n352) );
  HS65_LS_OAI212X5 U379 ( .A(n275), .B(n28), .C(n310), .D(n13), .E(n353), .Z(
        \chs_out_f[0][DATA][25] ) );
  HS65_LS_AOI222X2 U380 ( .A(n67), .B(\chs_in_f[2][DATA][25] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][25] ), .E(n51), .F(
        \chs_in_f[1][DATA][25] ), .Z(n353) );
  HS65_LS_OAI212X5 U381 ( .A(n274), .B(n28), .C(n309), .D(n13), .E(n354), .Z(
        \chs_out_f[0][DATA][26] ) );
  HS65_LS_AOI222X2 U382 ( .A(n67), .B(\chs_in_f[2][DATA][26] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][26] ), .E(n51), .F(
        \chs_in_f[1][DATA][26] ), .Z(n354) );
  HS65_LS_OAI212X5 U383 ( .A(n273), .B(n28), .C(n308), .D(n13), .E(n355), .Z(
        \chs_out_f[0][DATA][27] ) );
  HS65_LS_AOI222X2 U384 ( .A(n67), .B(\chs_in_f[2][DATA][27] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][27] ), .E(n51), .F(
        \chs_in_f[1][DATA][27] ), .Z(n355) );
  HS65_LS_OAI212X5 U385 ( .A(n272), .B(n28), .C(n307), .D(n13), .E(n356), .Z(
        \chs_out_f[0][DATA][28] ) );
  HS65_LS_AOI222X2 U386 ( .A(n67), .B(\chs_in_f[2][DATA][28] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][28] ), .E(n51), .F(
        \chs_in_f[1][DATA][28] ), .Z(n356) );
  HS65_LS_OAI212X5 U387 ( .A(n271), .B(n28), .C(n306), .D(n13), .E(n357), .Z(
        \chs_out_f[0][DATA][29] ) );
  HS65_LS_AOI222X2 U388 ( .A(n67), .B(\chs_in_f[2][DATA][29] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][29] ), .E(n51), .F(
        \chs_in_f[1][DATA][29] ), .Z(n357) );
  HS65_LS_OAI212X5 U389 ( .A(n270), .B(n28), .C(n305), .D(n13), .E(n359), .Z(
        \chs_out_f[0][DATA][30] ) );
  HS65_LS_AOI222X2 U390 ( .A(n67), .B(\chs_in_f[2][DATA][30] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][30] ), .E(n51), .F(
        \chs_in_f[1][DATA][30] ), .Z(n359) );
  HS65_LS_OAI212X5 U391 ( .A(n269), .B(n28), .C(n304), .D(n14), .E(n360), .Z(
        \chs_out_f[0][DATA][31] ) );
  HS65_LS_AOI222X2 U392 ( .A(n68), .B(\chs_in_f[2][DATA][31] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][31] ), .E(n52), .F(
        \chs_in_f[1][DATA][31] ), .Z(n360) );
  HS65_LS_OAI212X5 U393 ( .A(n268), .B(n28), .C(n303), .D(n14), .E(n361), .Z(
        \chs_out_f[0][DATA][32] ) );
  HS65_LS_AOI222X2 U394 ( .A(n68), .B(\chs_in_f[2][DATA][32] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][32] ), .E(n52), .F(
        \chs_in_f[1][DATA][32] ), .Z(n361) );
  HS65_LS_OAI212X5 U395 ( .A(n297), .B(n23), .C(n332), .D(n8), .E(n434), .Z(
        \chs_out_f[2][DATA][3] ) );
  HS65_LS_AOI222X2 U396 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][3] ), 
        .C(n40), .D(\chs_in_f[0][DATA][3] ), .E(n56), .F(
        \chs_in_f[1][DATA][3] ), .Z(n434) );
  HS65_LS_OAI212X5 U397 ( .A(n296), .B(n23), .C(n331), .D(n8), .E(n435), .Z(
        \chs_out_f[2][DATA][4] ) );
  HS65_LS_AOI222X2 U398 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][4] ), 
        .C(n40), .D(\chs_in_f[0][DATA][4] ), .E(n56), .F(
        \chs_in_f[1][DATA][4] ), .Z(n435) );
  HS65_LS_OAI212X5 U399 ( .A(n295), .B(n23), .C(n330), .D(n8), .E(n436), .Z(
        \chs_out_f[2][DATA][5] ) );
  HS65_LS_AOI222X2 U400 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][5] ), 
        .C(n40), .D(\chs_in_f[0][DATA][5] ), .E(n56), .F(
        \chs_in_f[1][DATA][5] ), .Z(n436) );
  HS65_LS_OAI212X5 U401 ( .A(n294), .B(n23), .C(n329), .D(n8), .E(n437), .Z(
        \chs_out_f[2][DATA][6] ) );
  HS65_LS_AOI222X2 U402 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][6] ), 
        .C(n40), .D(\chs_in_f[0][DATA][6] ), .E(n56), .F(
        \chs_in_f[1][DATA][6] ), .Z(n437) );
  HS65_LS_OAI212X5 U403 ( .A(n293), .B(n23), .C(n328), .D(n8), .E(n438), .Z(
        \chs_out_f[2][DATA][7] ) );
  HS65_LS_AOI222X2 U404 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][7] ), 
        .C(n40), .D(\chs_in_f[0][DATA][7] ), .E(n56), .F(
        \chs_in_f[1][DATA][7] ), .Z(n438) );
  HS65_LS_OAI212X5 U405 ( .A(n292), .B(n23), .C(n327), .D(n8), .E(n439), .Z(
        \chs_out_f[2][DATA][8] ) );
  HS65_LS_AOI222X2 U406 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][8] ), 
        .C(n40), .D(\chs_in_f[0][DATA][8] ), .E(n56), .F(
        \chs_in_f[1][DATA][8] ), .Z(n439) );
  HS65_LS_OAI212X5 U407 ( .A(n267), .B(n23), .C(n302), .D(n8), .E(n432), .Z(
        \chs_out_f[2][DATA][33] ) );
  HS65_LS_AOI222X2 U408 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][33] ), 
        .C(n40), .D(\chs_in_f[0][DATA][33] ), .E(n56), .F(
        \chs_in_f[1][DATA][33] ), .Z(n432) );
  HS65_LS_OAI212X5 U409 ( .A(n297), .B(n26), .C(n332), .D(n11), .E(n399), .Z(
        \chs_out_f[1][DATA][3] ) );
  HS65_LS_AOI222X2 U410 ( .A(n72), .B(\chs_in_f[2][DATA][3] ), .C(n36), .D(
        \chs_in_f[0][DATA][3] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][3] ), .Z(n399) );
  HS65_LS_OAI212X5 U411 ( .A(n296), .B(n26), .C(n331), .D(n11), .E(n400), .Z(
        \chs_out_f[1][DATA][4] ) );
  HS65_LS_AOI222X2 U412 ( .A(n72), .B(\chs_in_f[2][DATA][4] ), .C(n36), .D(
        \chs_in_f[0][DATA][4] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][4] ), .Z(n400) );
  HS65_LS_OAI212X5 U413 ( .A(n295), .B(n26), .C(n330), .D(n11), .E(n401), .Z(
        \chs_out_f[1][DATA][5] ) );
  HS65_LS_AOI222X2 U414 ( .A(n72), .B(\chs_in_f[2][DATA][5] ), .C(n36), .D(
        \chs_in_f[0][DATA][5] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][5] ), .Z(n401) );
  HS65_LS_OAI212X5 U415 ( .A(n294), .B(n26), .C(n329), .D(n11), .E(n402), .Z(
        \chs_out_f[1][DATA][6] ) );
  HS65_LS_AOI222X2 U416 ( .A(n72), .B(\chs_in_f[2][DATA][6] ), .C(n36), .D(
        \chs_in_f[0][DATA][6] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][6] ), .Z(n402) );
  HS65_LS_OAI212X5 U417 ( .A(n293), .B(n26), .C(n328), .D(n11), .E(n403), .Z(
        \chs_out_f[1][DATA][7] ) );
  HS65_LS_AOI222X2 U418 ( .A(n72), .B(\chs_in_f[2][DATA][7] ), .C(n36), .D(
        \chs_in_f[0][DATA][7] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][7] ), .Z(n403) );
  HS65_LS_OAI212X5 U419 ( .A(n292), .B(n26), .C(n327), .D(n11), .E(n404), .Z(
        \chs_out_f[1][DATA][8] ) );
  HS65_LS_AOI222X2 U420 ( .A(n72), .B(\chs_in_f[2][DATA][8] ), .C(n36), .D(
        \chs_in_f[0][DATA][8] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][8] ), .Z(n404) );
  HS65_LS_OAI212X5 U421 ( .A(n267), .B(n26), .C(n302), .D(n11), .E(n397), .Z(
        \chs_out_f[1][DATA][33] ) );
  HS65_LS_AOI222X2 U422 ( .A(n72), .B(\chs_in_f[2][DATA][33] ), .C(n36), .D(
        \chs_in_f[0][DATA][33] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][33] ), .Z(n397) );
  HS65_LS_OAI212X5 U423 ( .A(n297), .B(n29), .C(n332), .D(n14), .E(n364), .Z(
        \chs_out_f[0][DATA][3] ) );
  HS65_LS_AOI222X2 U424 ( .A(n68), .B(\chs_in_f[2][DATA][3] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][3] ), .E(n52), .F(
        \chs_in_f[1][DATA][3] ), .Z(n364) );
  HS65_LS_OAI212X5 U425 ( .A(n296), .B(n29), .C(n331), .D(n14), .E(n365), .Z(
        \chs_out_f[0][DATA][4] ) );
  HS65_LS_AOI222X2 U426 ( .A(n68), .B(\chs_in_f[2][DATA][4] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][4] ), .E(n52), .F(
        \chs_in_f[1][DATA][4] ), .Z(n365) );
  HS65_LS_OAI212X5 U427 ( .A(n295), .B(n29), .C(n330), .D(n14), .E(n366), .Z(
        \chs_out_f[0][DATA][5] ) );
  HS65_LS_AOI222X2 U428 ( .A(n68), .B(\chs_in_f[2][DATA][5] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][5] ), .E(n52), .F(
        \chs_in_f[1][DATA][5] ), .Z(n366) );
  HS65_LS_OAI212X5 U429 ( .A(n294), .B(n29), .C(n329), .D(n14), .E(n367), .Z(
        \chs_out_f[0][DATA][6] ) );
  HS65_LS_AOI222X2 U430 ( .A(n68), .B(\chs_in_f[2][DATA][6] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][6] ), .E(n52), .F(
        \chs_in_f[1][DATA][6] ), .Z(n367) );
  HS65_LS_OAI212X5 U431 ( .A(n293), .B(n29), .C(n328), .D(n14), .E(n368), .Z(
        \chs_out_f[0][DATA][7] ) );
  HS65_LS_AOI222X2 U432 ( .A(n68), .B(\chs_in_f[2][DATA][7] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][7] ), .E(n52), .F(
        \chs_in_f[1][DATA][7] ), .Z(n368) );
  HS65_LS_OAI212X5 U433 ( .A(n292), .B(n29), .C(n327), .D(n14), .E(n369), .Z(
        \chs_out_f[0][DATA][8] ) );
  HS65_LS_AOI222X2 U434 ( .A(n68), .B(\chs_in_f[2][DATA][8] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][8] ), .E(n52), .F(
        \chs_in_f[1][DATA][8] ), .Z(n369) );
  HS65_LS_OAI212X5 U435 ( .A(n267), .B(n29), .C(n302), .D(n14), .E(n362), .Z(
        \chs_out_f[0][DATA][33] ) );
  HS65_LS_AOI222X2 U436 ( .A(n68), .B(\chs_in_f[2][DATA][33] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][33] ), .E(n52), .F(
        \chs_in_f[1][DATA][33] ), .Z(n362) );
  HS65_LS_OAI212X5 U437 ( .A(n291), .B(n32), .C(n326), .D(n5), .E(n475), .Z(
        \chs_out_f[3][DATA][9] ) );
  HS65_LS_AOI222X2 U438 ( .A(n76), .B(\chs_in_f[2][DATA][9] ), .C(n44), .D(
        \chs_in_f[0][DATA][9] ), .E(n60), .F(\chs_in_f[1][DATA][9] ), .Z(n475)
         );
  HS65_LS_OAI212X5 U439 ( .A(n300), .B(n30), .C(n335), .D(n3), .E(n441), .Z(
        \chs_out_f[3][DATA][0] ) );
  HS65_LS_AOI222X2 U440 ( .A(n74), .B(\chs_in_f[2][DATA][0] ), .C(n42), .D(
        \chs_in_f[0][DATA][0] ), .E(n58), .F(\chs_in_f[1][DATA][0] ), .Z(n441)
         );
  HS65_LS_OAI212X5 U441 ( .A(n299), .B(n30), .C(n334), .D(n3), .E(n452), .Z(
        \chs_out_f[3][DATA][1] ) );
  HS65_LS_AOI222X2 U442 ( .A(n74), .B(\chs_in_f[2][DATA][1] ), .C(n42), .D(
        \chs_in_f[0][DATA][1] ), .E(n58), .F(\chs_in_f[1][DATA][1] ), .Z(n452)
         );
  HS65_LS_OAI212X5 U443 ( .A(n298), .B(n31), .C(n333), .D(n4), .E(n463), .Z(
        \chs_out_f[3][DATA][2] ) );
  HS65_LS_AOI222X2 U444 ( .A(n75), .B(\chs_in_f[2][DATA][2] ), .C(n43), .D(
        \chs_in_f[0][DATA][2] ), .E(n59), .F(\chs_in_f[1][DATA][2] ), .Z(n463)
         );
  HS65_LS_OAI212X5 U445 ( .A(n297), .B(n32), .C(n332), .D(n5), .E(n469), .Z(
        \chs_out_f[3][DATA][3] ) );
  HS65_LS_AOI222X2 U446 ( .A(n76), .B(\chs_in_f[2][DATA][3] ), .C(n44), .D(
        \chs_in_f[0][DATA][3] ), .E(n60), .F(\chs_in_f[1][DATA][3] ), .Z(n469)
         );
  HS65_LS_OAI212X5 U447 ( .A(n296), .B(n32), .C(n331), .D(n5), .E(n470), .Z(
        \chs_out_f[3][DATA][4] ) );
  HS65_LS_AOI222X2 U448 ( .A(n76), .B(\chs_in_f[2][DATA][4] ), .C(n44), .D(
        \chs_in_f[0][DATA][4] ), .E(n60), .F(\chs_in_f[1][DATA][4] ), .Z(n470)
         );
  HS65_LS_OAI212X5 U449 ( .A(n295), .B(n32), .C(n330), .D(n5), .E(n471), .Z(
        \chs_out_f[3][DATA][5] ) );
  HS65_LS_AOI222X2 U450 ( .A(n76), .B(\chs_in_f[2][DATA][5] ), .C(n44), .D(
        \chs_in_f[0][DATA][5] ), .E(n60), .F(\chs_in_f[1][DATA][5] ), .Z(n471)
         );
  HS65_LS_OAI212X5 U451 ( .A(n294), .B(n32), .C(n329), .D(n5), .E(n472), .Z(
        \chs_out_f[3][DATA][6] ) );
  HS65_LS_AOI222X2 U452 ( .A(n76), .B(\chs_in_f[2][DATA][6] ), .C(n44), .D(
        \chs_in_f[0][DATA][6] ), .E(n60), .F(\chs_in_f[1][DATA][6] ), .Z(n472)
         );
  HS65_LS_OAI212X5 U453 ( .A(n293), .B(n32), .C(n328), .D(n5), .E(n473), .Z(
        \chs_out_f[3][DATA][7] ) );
  HS65_LS_AOI222X2 U454 ( .A(n76), .B(\chs_in_f[2][DATA][7] ), .C(n44), .D(
        \chs_in_f[0][DATA][7] ), .E(n60), .F(\chs_in_f[1][DATA][7] ), .Z(n473)
         );
  HS65_LS_OAI212X5 U455 ( .A(n292), .B(n32), .C(n327), .D(n5), .E(n474), .Z(
        \chs_out_f[3][DATA][8] ) );
  HS65_LS_AOI222X2 U456 ( .A(n76), .B(\chs_in_f[2][DATA][8] ), .C(n44), .D(
        \chs_in_f[0][DATA][8] ), .E(n60), .F(\chs_in_f[1][DATA][8] ), .Z(n474)
         );
  HS65_LS_OAI212X5 U457 ( .A(n290), .B(n30), .C(n325), .D(n3), .E(n442), .Z(
        \chs_out_f[3][DATA][10] ) );
  HS65_LS_AOI222X2 U458 ( .A(n74), .B(\chs_in_f[2][DATA][10] ), .C(n42), .D(
        \chs_in_f[0][DATA][10] ), .E(n58), .F(\chs_in_f[1][DATA][10] ), .Z(
        n442) );
  HS65_LS_OAI212X5 U459 ( .A(n289), .B(n30), .C(n324), .D(n3), .E(n443), .Z(
        \chs_out_f[3][DATA][11] ) );
  HS65_LS_AOI222X2 U460 ( .A(n74), .B(\chs_in_f[2][DATA][11] ), .C(n42), .D(
        \chs_in_f[0][DATA][11] ), .E(n58), .F(\chs_in_f[1][DATA][11] ), .Z(
        n443) );
  HS65_LS_OAI212X5 U461 ( .A(n288), .B(n30), .C(n323), .D(n3), .E(n444), .Z(
        \chs_out_f[3][DATA][12] ) );
  HS65_LS_AOI222X2 U462 ( .A(n74), .B(\chs_in_f[2][DATA][12] ), .C(n42), .D(
        \chs_in_f[0][DATA][12] ), .E(n58), .F(\chs_in_f[1][DATA][12] ), .Z(
        n444) );
  HS65_LS_OAI212X5 U463 ( .A(n287), .B(n30), .C(n322), .D(n3), .E(n445), .Z(
        \chs_out_f[3][DATA][13] ) );
  HS65_LS_AOI222X2 U464 ( .A(n74), .B(\chs_in_f[2][DATA][13] ), .C(n42), .D(
        \chs_in_f[0][DATA][13] ), .E(n58), .F(\chs_in_f[1][DATA][13] ), .Z(
        n445) );
  HS65_LS_OAI212X5 U465 ( .A(n286), .B(n30), .C(n321), .D(n3), .E(n446), .Z(
        \chs_out_f[3][DATA][14] ) );
  HS65_LS_AOI222X2 U466 ( .A(n74), .B(\chs_in_f[2][DATA][14] ), .C(n42), .D(
        \chs_in_f[0][DATA][14] ), .E(n58), .F(\chs_in_f[1][DATA][14] ), .Z(
        n446) );
  HS65_LS_OAI212X5 U467 ( .A(n285), .B(n30), .C(n320), .D(n3), .E(n447), .Z(
        \chs_out_f[3][DATA][15] ) );
  HS65_LS_AOI222X2 U468 ( .A(n74), .B(\chs_in_f[2][DATA][15] ), .C(n42), .D(
        \chs_in_f[0][DATA][15] ), .E(n58), .F(\chs_in_f[1][DATA][15] ), .Z(
        n447) );
  HS65_LS_OAI212X5 U469 ( .A(n284), .B(n30), .C(n319), .D(n3), .E(n448), .Z(
        \chs_out_f[3][DATA][16] ) );
  HS65_LS_AOI222X2 U470 ( .A(n74), .B(\chs_in_f[2][DATA][16] ), .C(n42), .D(
        \chs_in_f[0][DATA][16] ), .E(n58), .F(\chs_in_f[1][DATA][16] ), .Z(
        n448) );
  HS65_LS_OAI212X5 U471 ( .A(n283), .B(n30), .C(n318), .D(n3), .E(n449), .Z(
        \chs_out_f[3][DATA][17] ) );
  HS65_LS_AOI222X2 U472 ( .A(n74), .B(\chs_in_f[2][DATA][17] ), .C(n42), .D(
        \chs_in_f[0][DATA][17] ), .E(n58), .F(\chs_in_f[1][DATA][17] ), .Z(
        n449) );
  HS65_LS_OAI212X5 U473 ( .A(n282), .B(n30), .C(n317), .D(n3), .E(n450), .Z(
        \chs_out_f[3][DATA][18] ) );
  HS65_LS_AOI222X2 U474 ( .A(n74), .B(\chs_in_f[2][DATA][18] ), .C(n42), .D(
        \chs_in_f[0][DATA][18] ), .E(n58), .F(\chs_in_f[1][DATA][18] ), .Z(
        n450) );
  HS65_LS_OAI212X5 U475 ( .A(n281), .B(n30), .C(n316), .D(n3), .E(n451), .Z(
        \chs_out_f[3][DATA][19] ) );
  HS65_LS_AOI222X2 U476 ( .A(n74), .B(\chs_in_f[2][DATA][19] ), .C(n42), .D(
        \chs_in_f[0][DATA][19] ), .E(n58), .F(\chs_in_f[1][DATA][19] ), .Z(
        n451) );
  HS65_LS_OAI212X5 U477 ( .A(n280), .B(n30), .C(n315), .D(n4), .E(n453), .Z(
        \chs_out_f[3][DATA][20] ) );
  HS65_LS_AOI222X2 U478 ( .A(n75), .B(\chs_in_f[2][DATA][20] ), .C(n43), .D(
        \chs_in_f[0][DATA][20] ), .E(n59), .F(\chs_in_f[1][DATA][20] ), .Z(
        n453) );
  HS65_LS_OAI212X5 U479 ( .A(n279), .B(n31), .C(n314), .D(n4), .E(n454), .Z(
        \chs_out_f[3][DATA][21] ) );
  HS65_LS_AOI222X2 U480 ( .A(n75), .B(\chs_in_f[2][DATA][21] ), .C(n43), .D(
        \chs_in_f[0][DATA][21] ), .E(n59), .F(\chs_in_f[1][DATA][21] ), .Z(
        n454) );
  HS65_LS_OAI212X5 U481 ( .A(n278), .B(n31), .C(n313), .D(n4), .E(n455), .Z(
        \chs_out_f[3][DATA][22] ) );
  HS65_LS_AOI222X2 U482 ( .A(n75), .B(\chs_in_f[2][DATA][22] ), .C(n43), .D(
        \chs_in_f[0][DATA][22] ), .E(n59), .F(\chs_in_f[1][DATA][22] ), .Z(
        n455) );
  HS65_LS_OAI212X5 U483 ( .A(n277), .B(n31), .C(n312), .D(n4), .E(n456), .Z(
        \chs_out_f[3][DATA][23] ) );
  HS65_LS_AOI222X2 U484 ( .A(n75), .B(\chs_in_f[2][DATA][23] ), .C(n43), .D(
        \chs_in_f[0][DATA][23] ), .E(n59), .F(\chs_in_f[1][DATA][23] ), .Z(
        n456) );
  HS65_LS_OAI212X5 U485 ( .A(n276), .B(n31), .C(n311), .D(n4), .E(n457), .Z(
        \chs_out_f[3][DATA][24] ) );
  HS65_LS_AOI222X2 U486 ( .A(n75), .B(\chs_in_f[2][DATA][24] ), .C(n43), .D(
        \chs_in_f[0][DATA][24] ), .E(n59), .F(\chs_in_f[1][DATA][24] ), .Z(
        n457) );
  HS65_LS_OAI212X5 U487 ( .A(n275), .B(n31), .C(n310), .D(n4), .E(n458), .Z(
        \chs_out_f[3][DATA][25] ) );
  HS65_LS_AOI222X2 U488 ( .A(n75), .B(\chs_in_f[2][DATA][25] ), .C(n43), .D(
        \chs_in_f[0][DATA][25] ), .E(n59), .F(\chs_in_f[1][DATA][25] ), .Z(
        n458) );
  HS65_LS_OAI212X5 U489 ( .A(n274), .B(n31), .C(n309), .D(n4), .E(n459), .Z(
        \chs_out_f[3][DATA][26] ) );
  HS65_LS_AOI222X2 U490 ( .A(n75), .B(\chs_in_f[2][DATA][26] ), .C(n43), .D(
        \chs_in_f[0][DATA][26] ), .E(n59), .F(\chs_in_f[1][DATA][26] ), .Z(
        n459) );
  HS65_LS_OAI212X5 U491 ( .A(n273), .B(n31), .C(n308), .D(n4), .E(n460), .Z(
        \chs_out_f[3][DATA][27] ) );
  HS65_LS_AOI222X2 U492 ( .A(n75), .B(\chs_in_f[2][DATA][27] ), .C(n43), .D(
        \chs_in_f[0][DATA][27] ), .E(n59), .F(\chs_in_f[1][DATA][27] ), .Z(
        n460) );
  HS65_LS_OAI212X5 U493 ( .A(n272), .B(n31), .C(n307), .D(n4), .E(n461), .Z(
        \chs_out_f[3][DATA][28] ) );
  HS65_LS_AOI222X2 U494 ( .A(n75), .B(\chs_in_f[2][DATA][28] ), .C(n43), .D(
        \chs_in_f[0][DATA][28] ), .E(n59), .F(\chs_in_f[1][DATA][28] ), .Z(
        n461) );
  HS65_LS_OAI212X5 U495 ( .A(n271), .B(n31), .C(n306), .D(n4), .E(n462), .Z(
        \chs_out_f[3][DATA][29] ) );
  HS65_LS_AOI222X2 U496 ( .A(n75), .B(\chs_in_f[2][DATA][29] ), .C(n43), .D(
        \chs_in_f[0][DATA][29] ), .E(n59), .F(\chs_in_f[1][DATA][29] ), .Z(
        n462) );
  HS65_LS_OAI212X5 U497 ( .A(n270), .B(n31), .C(n305), .D(n4), .E(n464), .Z(
        \chs_out_f[3][DATA][30] ) );
  HS65_LS_AOI222X2 U498 ( .A(n75), .B(\chs_in_f[2][DATA][30] ), .C(n43), .D(
        \chs_in_f[0][DATA][30] ), .E(n59), .F(\chs_in_f[1][DATA][30] ), .Z(
        n464) );
  HS65_LS_OAI212X5 U499 ( .A(n269), .B(n31), .C(n304), .D(n5), .E(n465), .Z(
        \chs_out_f[3][DATA][31] ) );
  HS65_LS_AOI222X2 U500 ( .A(n76), .B(\chs_in_f[2][DATA][31] ), .C(n44), .D(
        \chs_in_f[0][DATA][31] ), .E(n60), .F(\chs_in_f[1][DATA][31] ), .Z(
        n465) );
  HS65_LS_OAI212X5 U501 ( .A(n268), .B(n31), .C(n303), .D(n5), .E(n466), .Z(
        \chs_out_f[3][DATA][32] ) );
  HS65_LS_AOI222X2 U502 ( .A(n76), .B(\chs_in_f[2][DATA][32] ), .C(n44), .D(
        \chs_in_f[0][DATA][32] ), .E(n60), .F(\chs_in_f[1][DATA][32] ), .Z(
        n466) );
  HS65_LS_OAI212X5 U503 ( .A(n267), .B(n32), .C(n302), .D(n5), .E(n467), .Z(
        \chs_out_f[3][DATA][33] ) );
  HS65_LS_AOI222X2 U504 ( .A(n76), .B(\chs_in_f[2][DATA][33] ), .C(n44), .D(
        \chs_in_f[0][DATA][33] ), .E(n60), .F(\chs_in_f[1][DATA][33] ), .Z(
        n467) );
  HS65_LS_OAI212X5 U505 ( .A(n266), .B(n32), .C(n301), .D(n5), .E(n468), .Z(
        \chs_out_f[3][DATA][34] ) );
  HS65_LS_OAI212X5 U506 ( .A(n20), .B(n266), .C(n17), .D(n301), .E(n503), .Z(
        \chs_out_f[4][DATA][34] ) );
  HS65_LS_OAI212X5 U507 ( .A(n266), .B(n23), .C(n301), .D(n8), .E(n433), .Z(
        \chs_out_f[2][DATA][34] ) );
  HS65_LS_OAI212X5 U508 ( .A(n266), .B(n26), .C(n301), .D(n11), .E(n398), .Z(
        \chs_out_f[1][DATA][34] ) );
  HS65_LS_OAI212X5 U509 ( .A(n266), .B(n29), .C(n301), .D(n14), .E(n363), .Z(
        \chs_out_f[0][DATA][34] ) );
  HS65_LS_IVX9 U510 ( .A(\switch_sel[4][4] ), .Z(n260) );
  HS65_LS_IVX9 U511 ( .A(\switch_sel[3][3] ), .Z(n265) );
endmodule


module latch_controller_0_10 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_0_000000000_10 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, n3, n5, n6, n7, n8, n9, n10;
  assign N0 = preset;

  latch_controller_0_10 controller ( .preset(n6), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLQX9 type_out_reg ( .D(N4), .GN(n8), .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U8 ( .A(\left_in[DATA][34] ), .B(n3), .Z(n9) );
  HS65_LS_AND2X4 U7 ( .A(1'b0), .B(n7), .Z(n10) );
  HS65_LS_OR2X9 U9 ( .A(n10), .B(n9), .Z(N4) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(N39), .Q(\right_out[DATA][33] )
         );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(N38), .Q(\right_out[DATA][32] )
         );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(N37), .Q(\right_out[DATA][31] )
         );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(N36), .Q(\right_out[DATA][30] )
         );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(N35), .Q(\right_out[DATA][29] )
         );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(N34), .Q(\right_out[DATA][28] )
         );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(N33), .Q(\right_out[DATA][27] )
         );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(N32), .Q(\right_out[DATA][26] )
         );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(N31), .Q(\right_out[DATA][25] )
         );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(N30), .Q(\right_out[DATA][24] )
         );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(N29), .Q(\right_out[DATA][23] )
         );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(N28), .Q(\right_out[DATA][22] )
         );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(N27), .Q(\right_out[DATA][21] )
         );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(N26), .Q(\right_out[DATA][20] )
         );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(N25), .Q(\right_out[DATA][19] )
         );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(N24), .Q(\right_out[DATA][18] )
         );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(N23), .Q(\right_out[DATA][17] )
         );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(N22), .Q(\right_out[DATA][16] )
         );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(N21), .Q(\right_out[DATA][15] )
         );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(N20), .Q(\right_out[DATA][14] )
         );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(N19), .Q(\right_out[DATA][13] )
         );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(N18), .Q(\right_out[DATA][12] )
         );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(N17), .Q(\right_out[DATA][11] )
         );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(N16), .Q(\right_out[DATA][10] )
         );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(N15), .Q(\right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(N14), .Q(\right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(N13), .Q(\right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(N12), .Q(\right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(N11), .Q(\right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(N10), .Q(\right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(N9), .Q(\right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(N8), .Q(\right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(N7), .Q(\right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(N6), .Q(\right_out[DATA][0] ) );
  HS65_LS_BFX9 U3 ( .A(N0), .Z(n6) );
  HS65_LS_IVX9 U4 ( .A(n6), .Z(n3) );
  HS65_LS_IVX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_NOR2X6 U6 ( .A(lt_enable), .B(n7), .Z(n8) );
  HS65_LS_AND2X4 U10 ( .A(\left_in[DATA][9] ), .B(n3), .Z(N15) );
  HS65_LS_AND2X4 U11 ( .A(\left_in[DATA][0] ), .B(n3), .Z(N6) );
  HS65_LS_AND2X4 U12 ( .A(\left_in[DATA][1] ), .B(n5), .Z(N7) );
  HS65_LS_AND2X4 U13 ( .A(\left_in[DATA][2] ), .B(n3), .Z(N8) );
  HS65_LS_AND2X4 U14 ( .A(\left_in[DATA][3] ), .B(n5), .Z(N9) );
  HS65_LS_AND2X4 U15 ( .A(\left_in[DATA][4] ), .B(n3), .Z(N10) );
  HS65_LS_AND2X4 U16 ( .A(\left_in[DATA][5] ), .B(n3), .Z(N11) );
  HS65_LS_AND2X4 U17 ( .A(\left_in[DATA][6] ), .B(n3), .Z(N12) );
  HS65_LS_AND2X4 U18 ( .A(\left_in[DATA][7] ), .B(n3), .Z(N13) );
  HS65_LS_AND2X4 U19 ( .A(\left_in[DATA][8] ), .B(n3), .Z(N14) );
  HS65_LS_AND2X4 U20 ( .A(\left_in[DATA][10] ), .B(n3), .Z(N16) );
  HS65_LS_AND2X4 U21 ( .A(\left_in[DATA][11] ), .B(n3), .Z(N17) );
  HS65_LS_AND2X4 U22 ( .A(\left_in[DATA][12] ), .B(n3), .Z(N18) );
  HS65_LS_AND2X4 U23 ( .A(\left_in[DATA][13] ), .B(n3), .Z(N19) );
  HS65_LS_AND2X4 U24 ( .A(\left_in[DATA][14] ), .B(n3), .Z(N20) );
  HS65_LS_AND2X4 U25 ( .A(\left_in[DATA][15] ), .B(n3), .Z(N21) );
  HS65_LS_AND2X4 U26 ( .A(\left_in[DATA][16] ), .B(n3), .Z(N22) );
  HS65_LS_AND2X4 U27 ( .A(\left_in[DATA][17] ), .B(n5), .Z(N23) );
  HS65_LS_AND2X4 U28 ( .A(\left_in[DATA][18] ), .B(n5), .Z(N24) );
  HS65_LS_AND2X4 U29 ( .A(\left_in[DATA][19] ), .B(n5), .Z(N25) );
  HS65_LS_AND2X4 U30 ( .A(\left_in[DATA][20] ), .B(n5), .Z(N26) );
  HS65_LS_AND2X4 U31 ( .A(\left_in[DATA][21] ), .B(n5), .Z(N27) );
  HS65_LS_AND2X4 U32 ( .A(\left_in[DATA][22] ), .B(n5), .Z(N28) );
  HS65_LS_AND2X4 U33 ( .A(\left_in[DATA][23] ), .B(n5), .Z(N29) );
  HS65_LS_AND2X4 U34 ( .A(\left_in[DATA][24] ), .B(n5), .Z(N30) );
  HS65_LS_AND2X4 U35 ( .A(\left_in[DATA][25] ), .B(n5), .Z(N31) );
  HS65_LS_AND2X4 U36 ( .A(\left_in[DATA][26] ), .B(n5), .Z(N32) );
  HS65_LS_AND2X4 U37 ( .A(\left_in[DATA][27] ), .B(n5), .Z(N33) );
  HS65_LS_AND2X4 U38 ( .A(\left_in[DATA][28] ), .B(n5), .Z(N34) );
  HS65_LS_AND2X4 U39 ( .A(\left_in[DATA][29] ), .B(n5), .Z(N35) );
  HS65_LS_AND2X4 U40 ( .A(\left_in[DATA][30] ), .B(n3), .Z(N36) );
  HS65_LS_AND2X4 U41 ( .A(\left_in[DATA][31] ), .B(n5), .Z(N37) );
  HS65_LS_AND2X4 U42 ( .A(\left_in[DATA][32] ), .B(n3), .Z(N38) );
  HS65_LS_AND2X4 U43 ( .A(\left_in[DATA][33] ), .B(n5), .Z(N39) );
  HS65_LS_BFX9 U44 ( .A(N0), .Z(n7) );
  HS65_LS_NAND2X7 U45 ( .A(\right_out[DATA][34] ), .B(n8), .Z(N5) );
endmodule


module latch_controller_0_9 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_0_000000000_9 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, n3, n5, n6, n7, n8, n9, n10;
  assign N0 = preset;

  latch_controller_0_9 controller ( .preset(n6), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLQX9 type_out_reg ( .D(N4), .GN(n8), .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(1'b0), .B(n7), .Z(n10) );
  HS65_LS_OR2X9 U9 ( .A(n10), .B(n9), .Z(N4) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(N39), .Q(\right_out[DATA][33] )
         );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(N38), .Q(\right_out[DATA][32] )
         );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(N37), .Q(\right_out[DATA][31] )
         );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(N36), .Q(\right_out[DATA][30] )
         );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(N35), .Q(\right_out[DATA][29] )
         );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(N34), .Q(\right_out[DATA][28] )
         );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(N33), .Q(\right_out[DATA][27] )
         );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(N32), .Q(\right_out[DATA][26] )
         );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(N31), .Q(\right_out[DATA][25] )
         );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(N30), .Q(\right_out[DATA][24] )
         );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(N29), .Q(\right_out[DATA][23] )
         );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(N28), .Q(\right_out[DATA][22] )
         );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(N27), .Q(\right_out[DATA][21] )
         );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(N26), .Q(\right_out[DATA][20] )
         );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(N25), .Q(\right_out[DATA][19] )
         );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(N24), .Q(\right_out[DATA][18] )
         );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(N23), .Q(\right_out[DATA][17] )
         );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(N22), .Q(\right_out[DATA][16] )
         );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(N21), .Q(\right_out[DATA][15] )
         );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(N20), .Q(\right_out[DATA][14] )
         );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(N19), .Q(\right_out[DATA][13] )
         );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(N18), .Q(\right_out[DATA][12] )
         );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(N17), .Q(\right_out[DATA][11] )
         );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(N16), .Q(\right_out[DATA][10] )
         );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(N15), .Q(\right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(N14), .Q(\right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(N13), .Q(\right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(N12), .Q(\right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(N11), .Q(\right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(N10), .Q(\right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(N9), .Q(\right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(N8), .Q(\right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(N7), .Q(\right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(N6), .Q(\right_out[DATA][0] ) );
  HS65_LS_AND2X4 U8 ( .A(\left_in[DATA][34] ), .B(n3), .Z(n9) );
  HS65_LS_AND2X4 U3 ( .A(\left_in[DATA][0] ), .B(n3), .Z(N6) );
  HS65_LS_AND2X4 U4 ( .A(\left_in[DATA][1] ), .B(n5), .Z(N7) );
  HS65_LS_AND2X4 U5 ( .A(\left_in[DATA][2] ), .B(n3), .Z(N8) );
  HS65_LS_AND2X4 U6 ( .A(\left_in[DATA][10] ), .B(n3), .Z(N16) );
  HS65_LS_AND2X4 U10 ( .A(\left_in[DATA][11] ), .B(n3), .Z(N17) );
  HS65_LS_AND2X4 U11 ( .A(\left_in[DATA][12] ), .B(n3), .Z(N18) );
  HS65_LS_AND2X4 U12 ( .A(\left_in[DATA][13] ), .B(n3), .Z(N19) );
  HS65_LS_AND2X4 U13 ( .A(\left_in[DATA][14] ), .B(n3), .Z(N20) );
  HS65_LS_AND2X4 U14 ( .A(\left_in[DATA][15] ), .B(n3), .Z(N21) );
  HS65_LS_AND2X4 U15 ( .A(\left_in[DATA][3] ), .B(n5), .Z(N9) );
  HS65_LS_AND2X4 U16 ( .A(\left_in[DATA][4] ), .B(n3), .Z(N10) );
  HS65_LS_AND2X4 U17 ( .A(\left_in[DATA][5] ), .B(n3), .Z(N11) );
  HS65_LS_AND2X4 U18 ( .A(\left_in[DATA][6] ), .B(n3), .Z(N12) );
  HS65_LS_AND2X4 U19 ( .A(\left_in[DATA][7] ), .B(n3), .Z(N13) );
  HS65_LS_AND2X4 U20 ( .A(\left_in[DATA][8] ), .B(n3), .Z(N14) );
  HS65_LS_AND2X4 U21 ( .A(\left_in[DATA][9] ), .B(n3), .Z(N15) );
  HS65_LS_BFX9 U22 ( .A(N0), .Z(n6) );
  HS65_LS_IVX9 U23 ( .A(n6), .Z(n3) );
  HS65_LS_IVX9 U24 ( .A(n6), .Z(n5) );
  HS65_LS_NOR2X6 U25 ( .A(lt_enable), .B(n7), .Z(n8) );
  HS65_LS_AND2X4 U26 ( .A(\left_in[DATA][16] ), .B(n3), .Z(N22) );
  HS65_LS_AND2X4 U27 ( .A(\left_in[DATA][17] ), .B(n5), .Z(N23) );
  HS65_LS_AND2X4 U28 ( .A(\left_in[DATA][18] ), .B(n5), .Z(N24) );
  HS65_LS_AND2X4 U29 ( .A(\left_in[DATA][19] ), .B(n5), .Z(N25) );
  HS65_LS_AND2X4 U30 ( .A(\left_in[DATA][20] ), .B(n5), .Z(N26) );
  HS65_LS_AND2X4 U31 ( .A(\left_in[DATA][21] ), .B(n5), .Z(N27) );
  HS65_LS_AND2X4 U32 ( .A(\left_in[DATA][22] ), .B(n5), .Z(N28) );
  HS65_LS_AND2X4 U33 ( .A(\left_in[DATA][23] ), .B(n5), .Z(N29) );
  HS65_LS_AND2X4 U34 ( .A(\left_in[DATA][24] ), .B(n5), .Z(N30) );
  HS65_LS_AND2X4 U35 ( .A(\left_in[DATA][25] ), .B(n5), .Z(N31) );
  HS65_LS_AND2X4 U36 ( .A(\left_in[DATA][26] ), .B(n5), .Z(N32) );
  HS65_LS_AND2X4 U37 ( .A(\left_in[DATA][27] ), .B(n5), .Z(N33) );
  HS65_LS_AND2X4 U38 ( .A(\left_in[DATA][28] ), .B(n5), .Z(N34) );
  HS65_LS_AND2X4 U39 ( .A(\left_in[DATA][29] ), .B(n5), .Z(N35) );
  HS65_LS_AND2X4 U40 ( .A(\left_in[DATA][30] ), .B(n5), .Z(N36) );
  HS65_LS_AND2X4 U41 ( .A(\left_in[DATA][31] ), .B(n3), .Z(N37) );
  HS65_LS_AND2X4 U42 ( .A(\left_in[DATA][32] ), .B(n5), .Z(N38) );
  HS65_LS_AND2X4 U43 ( .A(\left_in[DATA][33] ), .B(n3), .Z(N39) );
  HS65_LS_BFX9 U44 ( .A(N0), .Z(n7) );
  HS65_LS_NAND2X7 U45 ( .A(\right_out[DATA][34] ), .B(n8), .Z(N5) );
endmodule


module latch_controller_0_8 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_0_000000000_8 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, n3, n5, n6, n7, n8, n9, n10;
  assign N0 = preset;

  latch_controller_0_8 controller ( .preset(n6), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLQX9 type_out_reg ( .D(N4), .GN(n8), .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U8 ( .A(\left_in[DATA][34] ), .B(n3), .Z(n9) );
  HS65_LS_AND2X4 U7 ( .A(1'b0), .B(n7), .Z(n10) );
  HS65_LS_OR2X9 U9 ( .A(n10), .B(n9), .Z(N4) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(N39), .Q(\right_out[DATA][33] )
         );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(N38), .Q(\right_out[DATA][32] )
         );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(N37), .Q(\right_out[DATA][31] )
         );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(N36), .Q(\right_out[DATA][30] )
         );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(N35), .Q(\right_out[DATA][29] )
         );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(N34), .Q(\right_out[DATA][28] )
         );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(N33), .Q(\right_out[DATA][27] )
         );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(N32), .Q(\right_out[DATA][26] )
         );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(N31), .Q(\right_out[DATA][25] )
         );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(N30), .Q(\right_out[DATA][24] )
         );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(N29), .Q(\right_out[DATA][23] )
         );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(N28), .Q(\right_out[DATA][22] )
         );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(N27), .Q(\right_out[DATA][21] )
         );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(N26), .Q(\right_out[DATA][20] )
         );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(N25), .Q(\right_out[DATA][19] )
         );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(N24), .Q(\right_out[DATA][18] )
         );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(N23), .Q(\right_out[DATA][17] )
         );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(N22), .Q(\right_out[DATA][16] )
         );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(N21), .Q(\right_out[DATA][15] )
         );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(N20), .Q(\right_out[DATA][14] )
         );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(N19), .Q(\right_out[DATA][13] )
         );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(N18), .Q(\right_out[DATA][12] )
         );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(N17), .Q(\right_out[DATA][11] )
         );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(N16), .Q(\right_out[DATA][10] )
         );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(N15), .Q(\right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(N14), .Q(\right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(N13), .Q(\right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(N12), .Q(\right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(N11), .Q(\right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(N10), .Q(\right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(N9), .Q(\right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(N8), .Q(\right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(N7), .Q(\right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(N6), .Q(\right_out[DATA][0] ) );
  HS65_LS_AND2X4 U3 ( .A(\left_in[DATA][4] ), .B(n3), .Z(N10) );
  HS65_LS_AND2X4 U4 ( .A(\left_in[DATA][5] ), .B(n3), .Z(N11) );
  HS65_LS_AND2X4 U5 ( .A(\left_in[DATA][6] ), .B(n3), .Z(N12) );
  HS65_LS_AND2X4 U6 ( .A(\left_in[DATA][7] ), .B(n3), .Z(N13) );
  HS65_LS_AND2X4 U10 ( .A(\left_in[DATA][8] ), .B(n3), .Z(N14) );
  HS65_LS_AND2X4 U11 ( .A(\left_in[DATA][9] ), .B(n3), .Z(N15) );
  HS65_LS_AND2X4 U12 ( .A(\left_in[DATA][10] ), .B(n3), .Z(N16) );
  HS65_LS_AND2X4 U13 ( .A(\left_in[DATA][11] ), .B(n3), .Z(N17) );
  HS65_LS_AND2X4 U14 ( .A(\left_in[DATA][12] ), .B(n3), .Z(N18) );
  HS65_LS_AND2X4 U15 ( .A(\left_in[DATA][13] ), .B(n3), .Z(N19) );
  HS65_LS_AND2X4 U16 ( .A(\left_in[DATA][14] ), .B(n3), .Z(N20) );
  HS65_LS_AND2X4 U17 ( .A(\left_in[DATA][15] ), .B(n3), .Z(N21) );
  HS65_LS_AND2X4 U18 ( .A(\left_in[DATA][0] ), .B(n3), .Z(N6) );
  HS65_LS_AND2X4 U19 ( .A(\left_in[DATA][1] ), .B(n5), .Z(N7) );
  HS65_LS_AND2X4 U20 ( .A(\left_in[DATA][2] ), .B(n3), .Z(N8) );
  HS65_LS_AND2X4 U21 ( .A(\left_in[DATA][3] ), .B(n5), .Z(N9) );
  HS65_LS_BFX9 U22 ( .A(N0), .Z(n6) );
  HS65_LS_IVX9 U23 ( .A(n6), .Z(n3) );
  HS65_LS_IVX9 U24 ( .A(n6), .Z(n5) );
  HS65_LS_NOR2X6 U25 ( .A(lt_enable), .B(n7), .Z(n8) );
  HS65_LS_AND2X4 U26 ( .A(\left_in[DATA][16] ), .B(n3), .Z(N22) );
  HS65_LS_AND2X4 U27 ( .A(\left_in[DATA][17] ), .B(n5), .Z(N23) );
  HS65_LS_AND2X4 U28 ( .A(\left_in[DATA][18] ), .B(n5), .Z(N24) );
  HS65_LS_AND2X4 U29 ( .A(\left_in[DATA][19] ), .B(n5), .Z(N25) );
  HS65_LS_AND2X4 U30 ( .A(\left_in[DATA][20] ), .B(n5), .Z(N26) );
  HS65_LS_AND2X4 U31 ( .A(\left_in[DATA][21] ), .B(n5), .Z(N27) );
  HS65_LS_AND2X4 U32 ( .A(\left_in[DATA][22] ), .B(n5), .Z(N28) );
  HS65_LS_AND2X4 U33 ( .A(\left_in[DATA][23] ), .B(n5), .Z(N29) );
  HS65_LS_AND2X4 U34 ( .A(\left_in[DATA][24] ), .B(n5), .Z(N30) );
  HS65_LS_AND2X4 U35 ( .A(\left_in[DATA][25] ), .B(n5), .Z(N31) );
  HS65_LS_AND2X4 U36 ( .A(\left_in[DATA][26] ), .B(n5), .Z(N32) );
  HS65_LS_AND2X4 U37 ( .A(\left_in[DATA][27] ), .B(n5), .Z(N33) );
  HS65_LS_AND2X4 U38 ( .A(\left_in[DATA][28] ), .B(n5), .Z(N34) );
  HS65_LS_AND2X4 U39 ( .A(\left_in[DATA][29] ), .B(n5), .Z(N35) );
  HS65_LS_AND2X4 U40 ( .A(\left_in[DATA][30] ), .B(n3), .Z(N36) );
  HS65_LS_AND2X4 U41 ( .A(\left_in[DATA][31] ), .B(n5), .Z(N37) );
  HS65_LS_AND2X4 U42 ( .A(\left_in[DATA][32] ), .B(n3), .Z(N38) );
  HS65_LS_AND2X4 U43 ( .A(\left_in[DATA][33] ), .B(n5), .Z(N39) );
  HS65_LS_BFX9 U44 ( .A(N0), .Z(n7) );
  HS65_LS_NAND2X7 U45 ( .A(\right_out[DATA][34] ), .B(n8), .Z(N5) );
endmodule


module latch_controller_0_7 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_0_000000000_7 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, n3, n5, n6, n7, n8, n9, n10;
  assign N0 = preset;

  latch_controller_0_7 controller ( .preset(n6), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLQX9 type_out_reg ( .D(N4), .GN(n8), .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U8 ( .A(\left_in[DATA][34] ), .B(n3), .Z(n9) );
  HS65_LS_AND2X4 U7 ( .A(1'b0), .B(n7), .Z(n10) );
  HS65_LS_OR2X9 U9 ( .A(n10), .B(n9), .Z(N4) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(N39), .Q(\right_out[DATA][33] )
         );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(N38), .Q(\right_out[DATA][32] )
         );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(N37), .Q(\right_out[DATA][31] )
         );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(N36), .Q(\right_out[DATA][30] )
         );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(N35), .Q(\right_out[DATA][29] )
         );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(N34), .Q(\right_out[DATA][28] )
         );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(N33), .Q(\right_out[DATA][27] )
         );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(N32), .Q(\right_out[DATA][26] )
         );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(N31), .Q(\right_out[DATA][25] )
         );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(N30), .Q(\right_out[DATA][24] )
         );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(N29), .Q(\right_out[DATA][23] )
         );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(N28), .Q(\right_out[DATA][22] )
         );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(N27), .Q(\right_out[DATA][21] )
         );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(N26), .Q(\right_out[DATA][20] )
         );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(N25), .Q(\right_out[DATA][19] )
         );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(N24), .Q(\right_out[DATA][18] )
         );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(N23), .Q(\right_out[DATA][17] )
         );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(N22), .Q(\right_out[DATA][16] )
         );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(N21), .Q(\right_out[DATA][15] )
         );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(N20), .Q(\right_out[DATA][14] )
         );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(N19), .Q(\right_out[DATA][13] )
         );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(N18), .Q(\right_out[DATA][12] )
         );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(N17), .Q(\right_out[DATA][11] )
         );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(N16), .Q(\right_out[DATA][10] )
         );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(N15), .Q(\right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(N14), .Q(\right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(N13), .Q(\right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(N12), .Q(\right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(N11), .Q(\right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(N10), .Q(\right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(N9), .Q(\right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(N8), .Q(\right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(N7), .Q(\right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(N6), .Q(\right_out[DATA][0] ) );
  HS65_LS_AND2X4 U3 ( .A(\left_in[DATA][4] ), .B(n3), .Z(N10) );
  HS65_LS_AND2X4 U4 ( .A(\left_in[DATA][5] ), .B(n3), .Z(N11) );
  HS65_LS_AND2X4 U5 ( .A(\left_in[DATA][6] ), .B(n3), .Z(N12) );
  HS65_LS_AND2X4 U6 ( .A(\left_in[DATA][7] ), .B(n3), .Z(N13) );
  HS65_LS_AND2X4 U10 ( .A(\left_in[DATA][8] ), .B(n3), .Z(N14) );
  HS65_LS_AND2X4 U11 ( .A(\left_in[DATA][9] ), .B(n3), .Z(N15) );
  HS65_LS_AND2X4 U12 ( .A(\left_in[DATA][10] ), .B(n3), .Z(N16) );
  HS65_LS_AND2X4 U13 ( .A(\left_in[DATA][11] ), .B(n3), .Z(N17) );
  HS65_LS_AND2X4 U14 ( .A(\left_in[DATA][12] ), .B(n3), .Z(N18) );
  HS65_LS_AND2X4 U15 ( .A(\left_in[DATA][13] ), .B(n3), .Z(N19) );
  HS65_LS_AND2X4 U16 ( .A(\left_in[DATA][14] ), .B(n3), .Z(N20) );
  HS65_LS_AND2X4 U17 ( .A(\left_in[DATA][15] ), .B(n3), .Z(N21) );
  HS65_LS_AND2X4 U18 ( .A(\left_in[DATA][0] ), .B(n3), .Z(N6) );
  HS65_LS_AND2X4 U19 ( .A(\left_in[DATA][1] ), .B(n5), .Z(N7) );
  HS65_LS_AND2X4 U20 ( .A(\left_in[DATA][2] ), .B(n3), .Z(N8) );
  HS65_LS_AND2X4 U21 ( .A(\left_in[DATA][3] ), .B(n5), .Z(N9) );
  HS65_LS_BFX9 U22 ( .A(N0), .Z(n6) );
  HS65_LS_IVX9 U23 ( .A(n6), .Z(n3) );
  HS65_LS_IVX9 U24 ( .A(n6), .Z(n5) );
  HS65_LS_NOR2X6 U25 ( .A(lt_enable), .B(n7), .Z(n8) );
  HS65_LS_AND2X4 U26 ( .A(\left_in[DATA][16] ), .B(n3), .Z(N22) );
  HS65_LS_AND2X4 U27 ( .A(\left_in[DATA][17] ), .B(n5), .Z(N23) );
  HS65_LS_AND2X4 U28 ( .A(\left_in[DATA][18] ), .B(n5), .Z(N24) );
  HS65_LS_AND2X4 U29 ( .A(\left_in[DATA][19] ), .B(n5), .Z(N25) );
  HS65_LS_AND2X4 U30 ( .A(\left_in[DATA][20] ), .B(n5), .Z(N26) );
  HS65_LS_AND2X4 U31 ( .A(\left_in[DATA][21] ), .B(n5), .Z(N27) );
  HS65_LS_AND2X4 U32 ( .A(\left_in[DATA][22] ), .B(n5), .Z(N28) );
  HS65_LS_AND2X4 U33 ( .A(\left_in[DATA][23] ), .B(n5), .Z(N29) );
  HS65_LS_AND2X4 U34 ( .A(\left_in[DATA][24] ), .B(n5), .Z(N30) );
  HS65_LS_AND2X4 U35 ( .A(\left_in[DATA][25] ), .B(n5), .Z(N31) );
  HS65_LS_AND2X4 U36 ( .A(\left_in[DATA][26] ), .B(n5), .Z(N32) );
  HS65_LS_AND2X4 U37 ( .A(\left_in[DATA][27] ), .B(n5), .Z(N33) );
  HS65_LS_AND2X4 U38 ( .A(\left_in[DATA][28] ), .B(n5), .Z(N34) );
  HS65_LS_AND2X4 U39 ( .A(\left_in[DATA][29] ), .B(n5), .Z(N35) );
  HS65_LS_AND2X4 U40 ( .A(\left_in[DATA][30] ), .B(n3), .Z(N36) );
  HS65_LS_AND2X4 U41 ( .A(\left_in[DATA][31] ), .B(n5), .Z(N37) );
  HS65_LS_AND2X4 U42 ( .A(\left_in[DATA][32] ), .B(n3), .Z(N38) );
  HS65_LS_AND2X4 U43 ( .A(\left_in[DATA][33] ), .B(n5), .Z(N39) );
  HS65_LS_BFX9 U44 ( .A(N0), .Z(n7) );
  HS65_LS_NAND2X7 U45 ( .A(\right_out[DATA][34] ), .B(n8), .Z(N5) );
endmodule


module latch_controller_0_6 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_0_000000000_6 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, n3, n5, n6, n7, n8, n9, n10;
  assign N0 = preset;

  latch_controller_0_6 controller ( .preset(n6), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLQX9 type_out_reg ( .D(N4), .GN(n8), .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U8 ( .A(\left_in[DATA][34] ), .B(n3), .Z(n9) );
  HS65_LS_AND2X4 U7 ( .A(1'b0), .B(n7), .Z(n10) );
  HS65_LS_OR2X9 U9 ( .A(n10), .B(n9), .Z(N4) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(N39), .Q(\right_out[DATA][33] )
         );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(N38), .Q(\right_out[DATA][32] )
         );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(N37), .Q(\right_out[DATA][31] )
         );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(N36), .Q(\right_out[DATA][30] )
         );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(N35), .Q(\right_out[DATA][29] )
         );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(N34), .Q(\right_out[DATA][28] )
         );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(N33), .Q(\right_out[DATA][27] )
         );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(N32), .Q(\right_out[DATA][26] )
         );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(N31), .Q(\right_out[DATA][25] )
         );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(N30), .Q(\right_out[DATA][24] )
         );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(N29), .Q(\right_out[DATA][23] )
         );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(N28), .Q(\right_out[DATA][22] )
         );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(N27), .Q(\right_out[DATA][21] )
         );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(N26), .Q(\right_out[DATA][20] )
         );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(N25), .Q(\right_out[DATA][19] )
         );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(N24), .Q(\right_out[DATA][18] )
         );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(N23), .Q(\right_out[DATA][17] )
         );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(N22), .Q(\right_out[DATA][16] )
         );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(N21), .Q(\right_out[DATA][15] )
         );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(N20), .Q(\right_out[DATA][14] )
         );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(N19), .Q(\right_out[DATA][13] )
         );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(N18), .Q(\right_out[DATA][12] )
         );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(N17), .Q(\right_out[DATA][11] )
         );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(N16), .Q(\right_out[DATA][10] )
         );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(N15), .Q(\right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(N14), .Q(\right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(N13), .Q(\right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(N12), .Q(\right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(N11), .Q(\right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(N10), .Q(\right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(N9), .Q(\right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(N8), .Q(\right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(N7), .Q(\right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(N6), .Q(\right_out[DATA][0] ) );
  HS65_LS_AND2X4 U3 ( .A(\left_in[DATA][5] ), .B(n3), .Z(N11) );
  HS65_LS_AND2X4 U4 ( .A(\left_in[DATA][6] ), .B(n3), .Z(N12) );
  HS65_LS_AND2X4 U5 ( .A(\left_in[DATA][7] ), .B(n3), .Z(N13) );
  HS65_LS_AND2X4 U6 ( .A(\left_in[DATA][8] ), .B(n3), .Z(N14) );
  HS65_LS_AND2X4 U10 ( .A(\left_in[DATA][14] ), .B(n3), .Z(N20) );
  HS65_LS_AND2X4 U11 ( .A(\left_in[DATA][15] ), .B(n3), .Z(N21) );
  HS65_LS_BFX9 U12 ( .A(N0), .Z(n6) );
  HS65_LS_IVX9 U13 ( .A(n6), .Z(n3) );
  HS65_LS_IVX9 U14 ( .A(n6), .Z(n5) );
  HS65_LS_NOR2X6 U15 ( .A(lt_enable), .B(n7), .Z(n8) );
  HS65_LS_AND2X4 U16 ( .A(\left_in[DATA][9] ), .B(n3), .Z(N15) );
  HS65_LS_AND2X4 U17 ( .A(\left_in[DATA][0] ), .B(n3), .Z(N6) );
  HS65_LS_AND2X4 U18 ( .A(\left_in[DATA][1] ), .B(n5), .Z(N7) );
  HS65_LS_AND2X4 U19 ( .A(\left_in[DATA][2] ), .B(n3), .Z(N8) );
  HS65_LS_AND2X4 U20 ( .A(\left_in[DATA][10] ), .B(n3), .Z(N16) );
  HS65_LS_AND2X4 U21 ( .A(\left_in[DATA][11] ), .B(n3), .Z(N17) );
  HS65_LS_AND2X4 U22 ( .A(\left_in[DATA][12] ), .B(n3), .Z(N18) );
  HS65_LS_AND2X4 U23 ( .A(\left_in[DATA][13] ), .B(n3), .Z(N19) );
  HS65_LS_AND2X4 U24 ( .A(\left_in[DATA][16] ), .B(n3), .Z(N22) );
  HS65_LS_AND2X4 U25 ( .A(\left_in[DATA][17] ), .B(n5), .Z(N23) );
  HS65_LS_AND2X4 U26 ( .A(\left_in[DATA][18] ), .B(n5), .Z(N24) );
  HS65_LS_AND2X4 U27 ( .A(\left_in[DATA][19] ), .B(n5), .Z(N25) );
  HS65_LS_AND2X4 U28 ( .A(\left_in[DATA][20] ), .B(n5), .Z(N26) );
  HS65_LS_AND2X4 U29 ( .A(\left_in[DATA][21] ), .B(n5), .Z(N27) );
  HS65_LS_AND2X4 U30 ( .A(\left_in[DATA][22] ), .B(n5), .Z(N28) );
  HS65_LS_AND2X4 U31 ( .A(\left_in[DATA][23] ), .B(n5), .Z(N29) );
  HS65_LS_AND2X4 U32 ( .A(\left_in[DATA][24] ), .B(n5), .Z(N30) );
  HS65_LS_AND2X4 U33 ( .A(\left_in[DATA][25] ), .B(n5), .Z(N31) );
  HS65_LS_AND2X4 U34 ( .A(\left_in[DATA][26] ), .B(n5), .Z(N32) );
  HS65_LS_AND2X4 U35 ( .A(\left_in[DATA][27] ), .B(n5), .Z(N33) );
  HS65_LS_AND2X4 U36 ( .A(\left_in[DATA][28] ), .B(n5), .Z(N34) );
  HS65_LS_AND2X4 U37 ( .A(\left_in[DATA][29] ), .B(n5), .Z(N35) );
  HS65_LS_AND2X4 U38 ( .A(\left_in[DATA][30] ), .B(n5), .Z(N36) );
  HS65_LS_AND2X4 U39 ( .A(\left_in[DATA][31] ), .B(n3), .Z(N37) );
  HS65_LS_AND2X4 U40 ( .A(\left_in[DATA][32] ), .B(n5), .Z(N38) );
  HS65_LS_AND2X4 U41 ( .A(\left_in[DATA][3] ), .B(n3), .Z(N9) );
  HS65_LS_AND2X4 U42 ( .A(\left_in[DATA][4] ), .B(n3), .Z(N10) );
  HS65_LS_AND2X4 U43 ( .A(\left_in[DATA][33] ), .B(n5), .Z(N39) );
  HS65_LS_BFX9 U44 ( .A(N0), .Z(n7) );
  HS65_LS_NAND2X7 U45 ( .A(\right_out[DATA][34] ), .B(n8), .Z(N5) );
endmodule


module crossbar_stage_2 ( preset, .switch_sel({\switch_sel[4][4] , 
        \switch_sel[4][3] , \switch_sel[4][2] , \switch_sel[4][1] , 
        \switch_sel[4][0] , \switch_sel[3][4] , \switch_sel[3][3] , 
        \switch_sel[3][2] , \switch_sel[3][1] , \switch_sel[3][0] , 
        \switch_sel[2][4] , \switch_sel[2][3] , \switch_sel[2][2] , 
        \switch_sel[2][1] , \switch_sel[2][0] , \switch_sel[1][4] , 
        \switch_sel[1][3] , \switch_sel[1][2] , \switch_sel[1][1] , 
        \switch_sel[1][0] , \switch_sel[0][4] , \switch_sel[0][3] , 
        \switch_sel[0][2] , \switch_sel[0][1] , \switch_sel[0][0] }), 
    .chs_in_f({\chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] , 
        \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] , 
        \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] , 
        \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] , 
        \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] , 
        \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] , 
        \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] , 
        \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] , 
        \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] , 
        \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] , 
        \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] , 
        \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] , 
        \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] , 
        \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] , \chs_in_f[4][DATA][7] , 
        \chs_in_f[4][DATA][6] , \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] , 
        \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] , \chs_in_f[4][DATA][1] , 
        \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] , \chs_in_f[3][DATA][34] , 
        \chs_in_f[3][DATA][33] , \chs_in_f[3][DATA][32] , 
        \chs_in_f[3][DATA][31] , \chs_in_f[3][DATA][30] , 
        \chs_in_f[3][DATA][29] , \chs_in_f[3][DATA][28] , 
        \chs_in_f[3][DATA][27] , \chs_in_f[3][DATA][26] , 
        \chs_in_f[3][DATA][25] , \chs_in_f[3][DATA][24] , 
        \chs_in_f[3][DATA][23] , \chs_in_f[3][DATA][22] , 
        \chs_in_f[3][DATA][21] , \chs_in_f[3][DATA][20] , 
        \chs_in_f[3][DATA][19] , \chs_in_f[3][DATA][18] , 
        \chs_in_f[3][DATA][17] , \chs_in_f[3][DATA][16] , 
        \chs_in_f[3][DATA][15] , \chs_in_f[3][DATA][14] , 
        \chs_in_f[3][DATA][13] , \chs_in_f[3][DATA][12] , 
        \chs_in_f[3][DATA][11] , \chs_in_f[3][DATA][10] , 
        \chs_in_f[3][DATA][9] , \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] , 
        \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] , \chs_in_f[3][DATA][4] , 
        \chs_in_f[3][DATA][3] , \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] , 
        \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] , 
        \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] , 
        \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] , 
        \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] , 
        \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] , 
        \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] , 
        \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] , 
        \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] , 
        \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] , 
        \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] , 
        \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] , 
        \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] , 
        \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] , 
        \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] , \chs_in_f[2][DATA][7] , 
        \chs_in_f[2][DATA][6] , \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] , 
        \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] , \chs_in_f[2][DATA][1] , 
        \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] , \chs_in_f[1][DATA][34] , 
        \chs_in_f[1][DATA][33] , \chs_in_f[1][DATA][32] , 
        \chs_in_f[1][DATA][31] , \chs_in_f[1][DATA][30] , 
        \chs_in_f[1][DATA][29] , \chs_in_f[1][DATA][28] , 
        \chs_in_f[1][DATA][27] , \chs_in_f[1][DATA][26] , 
        \chs_in_f[1][DATA][25] , \chs_in_f[1][DATA][24] , 
        \chs_in_f[1][DATA][23] , \chs_in_f[1][DATA][22] , 
        \chs_in_f[1][DATA][21] , \chs_in_f[1][DATA][20] , 
        \chs_in_f[1][DATA][19] , \chs_in_f[1][DATA][18] , 
        \chs_in_f[1][DATA][17] , \chs_in_f[1][DATA][16] , 
        \chs_in_f[1][DATA][15] , \chs_in_f[1][DATA][14] , 
        \chs_in_f[1][DATA][13] , \chs_in_f[1][DATA][12] , 
        \chs_in_f[1][DATA][11] , \chs_in_f[1][DATA][10] , 
        \chs_in_f[1][DATA][9] , \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] , 
        \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] , \chs_in_f[1][DATA][4] , 
        \chs_in_f[1][DATA][3] , \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] , 
        \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] , 
        \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] , 
        \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] , 
        \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] , 
        \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] , 
        \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] , 
        \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] , 
        \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] , 
        \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] , 
        \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] , 
        \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] , 
        \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] , 
        \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] , 
        \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] , \chs_in_f[0][DATA][7] , 
        \chs_in_f[0][DATA][6] , \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] , 
        \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] , \chs_in_f[0][DATA][1] , 
        \chs_in_f[0][DATA][0] }), .chs_in_b({\chs_in_b[4][ACK] , 
        \chs_in_b[3][ACK] , \chs_in_b[2][ACK] , \chs_in_b[1][ACK] , 
        \chs_in_b[0][ACK] }), .latches_out_f({\latches_out_f[4][REQ] , 
        \latches_out_f[4][DATA][34] , \latches_out_f[4][DATA][33] , 
        \latches_out_f[4][DATA][32] , \latches_out_f[4][DATA][31] , 
        \latches_out_f[4][DATA][30] , \latches_out_f[4][DATA][29] , 
        \latches_out_f[4][DATA][28] , \latches_out_f[4][DATA][27] , 
        \latches_out_f[4][DATA][26] , \latches_out_f[4][DATA][25] , 
        \latches_out_f[4][DATA][24] , \latches_out_f[4][DATA][23] , 
        \latches_out_f[4][DATA][22] , \latches_out_f[4][DATA][21] , 
        \latches_out_f[4][DATA][20] , \latches_out_f[4][DATA][19] , 
        \latches_out_f[4][DATA][18] , \latches_out_f[4][DATA][17] , 
        \latches_out_f[4][DATA][16] , \latches_out_f[4][DATA][15] , 
        \latches_out_f[4][DATA][14] , \latches_out_f[4][DATA][13] , 
        \latches_out_f[4][DATA][12] , \latches_out_f[4][DATA][11] , 
        \latches_out_f[4][DATA][10] , \latches_out_f[4][DATA][9] , 
        \latches_out_f[4][DATA][8] , \latches_out_f[4][DATA][7] , 
        \latches_out_f[4][DATA][6] , \latches_out_f[4][DATA][5] , 
        \latches_out_f[4][DATA][4] , \latches_out_f[4][DATA][3] , 
        \latches_out_f[4][DATA][2] , \latches_out_f[4][DATA][1] , 
        \latches_out_f[4][DATA][0] , \latches_out_f[3][REQ] , 
        \latches_out_f[3][DATA][34] , \latches_out_f[3][DATA][33] , 
        \latches_out_f[3][DATA][32] , \latches_out_f[3][DATA][31] , 
        \latches_out_f[3][DATA][30] , \latches_out_f[3][DATA][29] , 
        \latches_out_f[3][DATA][28] , \latches_out_f[3][DATA][27] , 
        \latches_out_f[3][DATA][26] , \latches_out_f[3][DATA][25] , 
        \latches_out_f[3][DATA][24] , \latches_out_f[3][DATA][23] , 
        \latches_out_f[3][DATA][22] , \latches_out_f[3][DATA][21] , 
        \latches_out_f[3][DATA][20] , \latches_out_f[3][DATA][19] , 
        \latches_out_f[3][DATA][18] , \latches_out_f[3][DATA][17] , 
        \latches_out_f[3][DATA][16] , \latches_out_f[3][DATA][15] , 
        \latches_out_f[3][DATA][14] , \latches_out_f[3][DATA][13] , 
        \latches_out_f[3][DATA][12] , \latches_out_f[3][DATA][11] , 
        \latches_out_f[3][DATA][10] , \latches_out_f[3][DATA][9] , 
        \latches_out_f[3][DATA][8] , \latches_out_f[3][DATA][7] , 
        \latches_out_f[3][DATA][6] , \latches_out_f[3][DATA][5] , 
        \latches_out_f[3][DATA][4] , \latches_out_f[3][DATA][3] , 
        \latches_out_f[3][DATA][2] , \latches_out_f[3][DATA][1] , 
        \latches_out_f[3][DATA][0] , \latches_out_f[2][REQ] , 
        \latches_out_f[2][DATA][34] , \latches_out_f[2][DATA][33] , 
        \latches_out_f[2][DATA][32] , \latches_out_f[2][DATA][31] , 
        \latches_out_f[2][DATA][30] , \latches_out_f[2][DATA][29] , 
        \latches_out_f[2][DATA][28] , \latches_out_f[2][DATA][27] , 
        \latches_out_f[2][DATA][26] , \latches_out_f[2][DATA][25] , 
        \latches_out_f[2][DATA][24] , \latches_out_f[2][DATA][23] , 
        \latches_out_f[2][DATA][22] , \latches_out_f[2][DATA][21] , 
        \latches_out_f[2][DATA][20] , \latches_out_f[2][DATA][19] , 
        \latches_out_f[2][DATA][18] , \latches_out_f[2][DATA][17] , 
        \latches_out_f[2][DATA][16] , \latches_out_f[2][DATA][15] , 
        \latches_out_f[2][DATA][14] , \latches_out_f[2][DATA][13] , 
        \latches_out_f[2][DATA][12] , \latches_out_f[2][DATA][11] , 
        \latches_out_f[2][DATA][10] , \latches_out_f[2][DATA][9] , 
        \latches_out_f[2][DATA][8] , \latches_out_f[2][DATA][7] , 
        \latches_out_f[2][DATA][6] , \latches_out_f[2][DATA][5] , 
        \latches_out_f[2][DATA][4] , \latches_out_f[2][DATA][3] , 
        \latches_out_f[2][DATA][2] , \latches_out_f[2][DATA][1] , 
        \latches_out_f[2][DATA][0] , \latches_out_f[1][REQ] , 
        \latches_out_f[1][DATA][34] , \latches_out_f[1][DATA][33] , 
        \latches_out_f[1][DATA][32] , \latches_out_f[1][DATA][31] , 
        \latches_out_f[1][DATA][30] , \latches_out_f[1][DATA][29] , 
        \latches_out_f[1][DATA][28] , \latches_out_f[1][DATA][27] , 
        \latches_out_f[1][DATA][26] , \latches_out_f[1][DATA][25] , 
        \latches_out_f[1][DATA][24] , \latches_out_f[1][DATA][23] , 
        \latches_out_f[1][DATA][22] , \latches_out_f[1][DATA][21] , 
        \latches_out_f[1][DATA][20] , \latches_out_f[1][DATA][19] , 
        \latches_out_f[1][DATA][18] , \latches_out_f[1][DATA][17] , 
        \latches_out_f[1][DATA][16] , \latches_out_f[1][DATA][15] , 
        \latches_out_f[1][DATA][14] , \latches_out_f[1][DATA][13] , 
        \latches_out_f[1][DATA][12] , \latches_out_f[1][DATA][11] , 
        \latches_out_f[1][DATA][10] , \latches_out_f[1][DATA][9] , 
        \latches_out_f[1][DATA][8] , \latches_out_f[1][DATA][7] , 
        \latches_out_f[1][DATA][6] , \latches_out_f[1][DATA][5] , 
        \latches_out_f[1][DATA][4] , \latches_out_f[1][DATA][3] , 
        \latches_out_f[1][DATA][2] , \latches_out_f[1][DATA][1] , 
        \latches_out_f[1][DATA][0] , \latches_out_f[0][REQ] , 
        \latches_out_f[0][DATA][34] , \latches_out_f[0][DATA][33] , 
        \latches_out_f[0][DATA][32] , \latches_out_f[0][DATA][31] , 
        \latches_out_f[0][DATA][30] , \latches_out_f[0][DATA][29] , 
        \latches_out_f[0][DATA][28] , \latches_out_f[0][DATA][27] , 
        \latches_out_f[0][DATA][26] , \latches_out_f[0][DATA][25] , 
        \latches_out_f[0][DATA][24] , \latches_out_f[0][DATA][23] , 
        \latches_out_f[0][DATA][22] , \latches_out_f[0][DATA][21] , 
        \latches_out_f[0][DATA][20] , \latches_out_f[0][DATA][19] , 
        \latches_out_f[0][DATA][18] , \latches_out_f[0][DATA][17] , 
        \latches_out_f[0][DATA][16] , \latches_out_f[0][DATA][15] , 
        \latches_out_f[0][DATA][14] , \latches_out_f[0][DATA][13] , 
        \latches_out_f[0][DATA][12] , \latches_out_f[0][DATA][11] , 
        \latches_out_f[0][DATA][10] , \latches_out_f[0][DATA][9] , 
        \latches_out_f[0][DATA][8] , \latches_out_f[0][DATA][7] , 
        \latches_out_f[0][DATA][6] , \latches_out_f[0][DATA][5] , 
        \latches_out_f[0][DATA][4] , \latches_out_f[0][DATA][3] , 
        \latches_out_f[0][DATA][2] , \latches_out_f[0][DATA][1] , 
        \latches_out_f[0][DATA][0] }), .latches_out_b({\latches_out_b[4][ACK] , 
        \latches_out_b[3][ACK] , \latches_out_b[2][ACK] , 
        \latches_out_b[1][ACK] , \latches_out_b[0][ACK] }) );
  input preset, \switch_sel[4][4] , \switch_sel[4][3] , \switch_sel[4][2] ,
         \switch_sel[4][1] , \switch_sel[4][0] , \switch_sel[3][4] ,
         \switch_sel[3][3] , \switch_sel[3][2] , \switch_sel[3][1] ,
         \switch_sel[3][0] , \switch_sel[2][4] , \switch_sel[2][3] ,
         \switch_sel[2][2] , \switch_sel[2][1] , \switch_sel[2][0] ,
         \switch_sel[1][4] , \switch_sel[1][3] , \switch_sel[1][2] ,
         \switch_sel[1][1] , \switch_sel[1][0] , \switch_sel[0][4] ,
         \switch_sel[0][3] , \switch_sel[0][2] , \switch_sel[0][1] ,
         \switch_sel[0][0] , \chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] ,
         \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] ,
         \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] ,
         \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] ,
         \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] ,
         \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] ,
         \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] ,
         \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] ,
         \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] ,
         \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] ,
         \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] ,
         \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] ,
         \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] ,
         \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] ,
         \chs_in_f[4][DATA][7] , \chs_in_f[4][DATA][6] ,
         \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] ,
         \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] ,
         \chs_in_f[4][DATA][1] , \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] ,
         \chs_in_f[3][DATA][34] , \chs_in_f[3][DATA][33] ,
         \chs_in_f[3][DATA][32] , \chs_in_f[3][DATA][31] ,
         \chs_in_f[3][DATA][30] , \chs_in_f[3][DATA][29] ,
         \chs_in_f[3][DATA][28] , \chs_in_f[3][DATA][27] ,
         \chs_in_f[3][DATA][26] , \chs_in_f[3][DATA][25] ,
         \chs_in_f[3][DATA][24] , \chs_in_f[3][DATA][23] ,
         \chs_in_f[3][DATA][22] , \chs_in_f[3][DATA][21] ,
         \chs_in_f[3][DATA][20] , \chs_in_f[3][DATA][19] ,
         \chs_in_f[3][DATA][18] , \chs_in_f[3][DATA][17] ,
         \chs_in_f[3][DATA][16] , \chs_in_f[3][DATA][15] ,
         \chs_in_f[3][DATA][14] , \chs_in_f[3][DATA][13] ,
         \chs_in_f[3][DATA][12] , \chs_in_f[3][DATA][11] ,
         \chs_in_f[3][DATA][10] , \chs_in_f[3][DATA][9] ,
         \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] ,
         \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] ,
         \chs_in_f[3][DATA][4] , \chs_in_f[3][DATA][3] ,
         \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] ,
         \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] ,
         \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] ,
         \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] ,
         \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] ,
         \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] ,
         \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] ,
         \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] ,
         \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] ,
         \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] ,
         \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] ,
         \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] ,
         \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] ,
         \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] ,
         \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] ,
         \chs_in_f[2][DATA][7] , \chs_in_f[2][DATA][6] ,
         \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] ,
         \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] ,
         \chs_in_f[2][DATA][1] , \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] ,
         \chs_in_f[1][DATA][34] , \chs_in_f[1][DATA][33] ,
         \chs_in_f[1][DATA][32] , \chs_in_f[1][DATA][31] ,
         \chs_in_f[1][DATA][30] , \chs_in_f[1][DATA][29] ,
         \chs_in_f[1][DATA][28] , \chs_in_f[1][DATA][27] ,
         \chs_in_f[1][DATA][26] , \chs_in_f[1][DATA][25] ,
         \chs_in_f[1][DATA][24] , \chs_in_f[1][DATA][23] ,
         \chs_in_f[1][DATA][22] , \chs_in_f[1][DATA][21] ,
         \chs_in_f[1][DATA][20] , \chs_in_f[1][DATA][19] ,
         \chs_in_f[1][DATA][18] , \chs_in_f[1][DATA][17] ,
         \chs_in_f[1][DATA][16] , \chs_in_f[1][DATA][15] ,
         \chs_in_f[1][DATA][14] , \chs_in_f[1][DATA][13] ,
         \chs_in_f[1][DATA][12] , \chs_in_f[1][DATA][11] ,
         \chs_in_f[1][DATA][10] , \chs_in_f[1][DATA][9] ,
         \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] ,
         \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] ,
         \chs_in_f[1][DATA][4] , \chs_in_f[1][DATA][3] ,
         \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] ,
         \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] ,
         \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] ,
         \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] ,
         \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] ,
         \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] ,
         \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] ,
         \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] ,
         \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] ,
         \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] ,
         \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] ,
         \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] ,
         \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] ,
         \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] ,
         \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] ,
         \chs_in_f[0][DATA][7] , \chs_in_f[0][DATA][6] ,
         \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] ,
         \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] ,
         \chs_in_f[0][DATA][1] , \chs_in_f[0][DATA][0] ,
         \latches_out_b[4][ACK] , \latches_out_b[3][ACK] ,
         \latches_out_b[2][ACK] , \latches_out_b[1][ACK] ,
         \latches_out_b[0][ACK] ;
  output \chs_in_b[4][ACK] , \chs_in_b[3][ACK] , \chs_in_b[2][ACK] ,
         \chs_in_b[1][ACK] , \chs_in_b[0][ACK] , \latches_out_f[4][REQ] ,
         \latches_out_f[4][DATA][34] , \latches_out_f[4][DATA][33] ,
         \latches_out_f[4][DATA][32] , \latches_out_f[4][DATA][31] ,
         \latches_out_f[4][DATA][30] , \latches_out_f[4][DATA][29] ,
         \latches_out_f[4][DATA][28] , \latches_out_f[4][DATA][27] ,
         \latches_out_f[4][DATA][26] , \latches_out_f[4][DATA][25] ,
         \latches_out_f[4][DATA][24] , \latches_out_f[4][DATA][23] ,
         \latches_out_f[4][DATA][22] , \latches_out_f[4][DATA][21] ,
         \latches_out_f[4][DATA][20] , \latches_out_f[4][DATA][19] ,
         \latches_out_f[4][DATA][18] , \latches_out_f[4][DATA][17] ,
         \latches_out_f[4][DATA][16] , \latches_out_f[4][DATA][15] ,
         \latches_out_f[4][DATA][14] , \latches_out_f[4][DATA][13] ,
         \latches_out_f[4][DATA][12] , \latches_out_f[4][DATA][11] ,
         \latches_out_f[4][DATA][10] , \latches_out_f[4][DATA][9] ,
         \latches_out_f[4][DATA][8] , \latches_out_f[4][DATA][7] ,
         \latches_out_f[4][DATA][6] , \latches_out_f[4][DATA][5] ,
         \latches_out_f[4][DATA][4] , \latches_out_f[4][DATA][3] ,
         \latches_out_f[4][DATA][2] , \latches_out_f[4][DATA][1] ,
         \latches_out_f[4][DATA][0] , \latches_out_f[3][REQ] ,
         \latches_out_f[3][DATA][34] , \latches_out_f[3][DATA][33] ,
         \latches_out_f[3][DATA][32] , \latches_out_f[3][DATA][31] ,
         \latches_out_f[3][DATA][30] , \latches_out_f[3][DATA][29] ,
         \latches_out_f[3][DATA][28] , \latches_out_f[3][DATA][27] ,
         \latches_out_f[3][DATA][26] , \latches_out_f[3][DATA][25] ,
         \latches_out_f[3][DATA][24] , \latches_out_f[3][DATA][23] ,
         \latches_out_f[3][DATA][22] , \latches_out_f[3][DATA][21] ,
         \latches_out_f[3][DATA][20] , \latches_out_f[3][DATA][19] ,
         \latches_out_f[3][DATA][18] , \latches_out_f[3][DATA][17] ,
         \latches_out_f[3][DATA][16] , \latches_out_f[3][DATA][15] ,
         \latches_out_f[3][DATA][14] , \latches_out_f[3][DATA][13] ,
         \latches_out_f[3][DATA][12] , \latches_out_f[3][DATA][11] ,
         \latches_out_f[3][DATA][10] , \latches_out_f[3][DATA][9] ,
         \latches_out_f[3][DATA][8] , \latches_out_f[3][DATA][7] ,
         \latches_out_f[3][DATA][6] , \latches_out_f[3][DATA][5] ,
         \latches_out_f[3][DATA][4] , \latches_out_f[3][DATA][3] ,
         \latches_out_f[3][DATA][2] , \latches_out_f[3][DATA][1] ,
         \latches_out_f[3][DATA][0] , \latches_out_f[2][REQ] ,
         \latches_out_f[2][DATA][34] , \latches_out_f[2][DATA][33] ,
         \latches_out_f[2][DATA][32] , \latches_out_f[2][DATA][31] ,
         \latches_out_f[2][DATA][30] , \latches_out_f[2][DATA][29] ,
         \latches_out_f[2][DATA][28] , \latches_out_f[2][DATA][27] ,
         \latches_out_f[2][DATA][26] , \latches_out_f[2][DATA][25] ,
         \latches_out_f[2][DATA][24] , \latches_out_f[2][DATA][23] ,
         \latches_out_f[2][DATA][22] , \latches_out_f[2][DATA][21] ,
         \latches_out_f[2][DATA][20] , \latches_out_f[2][DATA][19] ,
         \latches_out_f[2][DATA][18] , \latches_out_f[2][DATA][17] ,
         \latches_out_f[2][DATA][16] , \latches_out_f[2][DATA][15] ,
         \latches_out_f[2][DATA][14] , \latches_out_f[2][DATA][13] ,
         \latches_out_f[2][DATA][12] , \latches_out_f[2][DATA][11] ,
         \latches_out_f[2][DATA][10] , \latches_out_f[2][DATA][9] ,
         \latches_out_f[2][DATA][8] , \latches_out_f[2][DATA][7] ,
         \latches_out_f[2][DATA][6] , \latches_out_f[2][DATA][5] ,
         \latches_out_f[2][DATA][4] , \latches_out_f[2][DATA][3] ,
         \latches_out_f[2][DATA][2] , \latches_out_f[2][DATA][1] ,
         \latches_out_f[2][DATA][0] , \latches_out_f[1][REQ] ,
         \latches_out_f[1][DATA][34] , \latches_out_f[1][DATA][33] ,
         \latches_out_f[1][DATA][32] , \latches_out_f[1][DATA][31] ,
         \latches_out_f[1][DATA][30] , \latches_out_f[1][DATA][29] ,
         \latches_out_f[1][DATA][28] , \latches_out_f[1][DATA][27] ,
         \latches_out_f[1][DATA][26] , \latches_out_f[1][DATA][25] ,
         \latches_out_f[1][DATA][24] , \latches_out_f[1][DATA][23] ,
         \latches_out_f[1][DATA][22] , \latches_out_f[1][DATA][21] ,
         \latches_out_f[1][DATA][20] , \latches_out_f[1][DATA][19] ,
         \latches_out_f[1][DATA][18] , \latches_out_f[1][DATA][17] ,
         \latches_out_f[1][DATA][16] , \latches_out_f[1][DATA][15] ,
         \latches_out_f[1][DATA][14] , \latches_out_f[1][DATA][13] ,
         \latches_out_f[1][DATA][12] , \latches_out_f[1][DATA][11] ,
         \latches_out_f[1][DATA][10] , \latches_out_f[1][DATA][9] ,
         \latches_out_f[1][DATA][8] , \latches_out_f[1][DATA][7] ,
         \latches_out_f[1][DATA][6] , \latches_out_f[1][DATA][5] ,
         \latches_out_f[1][DATA][4] , \latches_out_f[1][DATA][3] ,
         \latches_out_f[1][DATA][2] , \latches_out_f[1][DATA][1] ,
         \latches_out_f[1][DATA][0] , \latches_out_f[0][REQ] ,
         \latches_out_f[0][DATA][34] , \latches_out_f[0][DATA][33] ,
         \latches_out_f[0][DATA][32] , \latches_out_f[0][DATA][31] ,
         \latches_out_f[0][DATA][30] , \latches_out_f[0][DATA][29] ,
         \latches_out_f[0][DATA][28] , \latches_out_f[0][DATA][27] ,
         \latches_out_f[0][DATA][26] , \latches_out_f[0][DATA][25] ,
         \latches_out_f[0][DATA][24] , \latches_out_f[0][DATA][23] ,
         \latches_out_f[0][DATA][22] , \latches_out_f[0][DATA][21] ,
         \latches_out_f[0][DATA][20] , \latches_out_f[0][DATA][19] ,
         \latches_out_f[0][DATA][18] , \latches_out_f[0][DATA][17] ,
         \latches_out_f[0][DATA][16] , \latches_out_f[0][DATA][15] ,
         \latches_out_f[0][DATA][14] , \latches_out_f[0][DATA][13] ,
         \latches_out_f[0][DATA][12] , \latches_out_f[0][DATA][11] ,
         \latches_out_f[0][DATA][10] , \latches_out_f[0][DATA][9] ,
         \latches_out_f[0][DATA][8] , \latches_out_f[0][DATA][7] ,
         \latches_out_f[0][DATA][6] , \latches_out_f[0][DATA][5] ,
         \latches_out_f[0][DATA][4] , \latches_out_f[0][DATA][3] ,
         \latches_out_f[0][DATA][2] , \latches_out_f[0][DATA][1] ,
         \latches_out_f[0][DATA][0] ;
  wire   \latches_in_f[4][REQ] , \latches_in_f[4][DATA][34] ,
         \latches_in_f[4][DATA][33] , \latches_in_f[4][DATA][32] ,
         \latches_in_f[4][DATA][31] , \latches_in_f[4][DATA][30] ,
         \latches_in_f[4][DATA][29] , \latches_in_f[4][DATA][28] ,
         \latches_in_f[4][DATA][27] , \latches_in_f[4][DATA][26] ,
         \latches_in_f[4][DATA][25] , \latches_in_f[4][DATA][24] ,
         \latches_in_f[4][DATA][23] , \latches_in_f[4][DATA][22] ,
         \latches_in_f[4][DATA][21] , \latches_in_f[4][DATA][20] ,
         \latches_in_f[4][DATA][19] , \latches_in_f[4][DATA][18] ,
         \latches_in_f[4][DATA][17] , \latches_in_f[4][DATA][16] ,
         \latches_in_f[4][DATA][15] , \latches_in_f[4][DATA][14] ,
         \latches_in_f[4][DATA][13] , \latches_in_f[4][DATA][12] ,
         \latches_in_f[4][DATA][11] , \latches_in_f[4][DATA][10] ,
         \latches_in_f[4][DATA][9] , \latches_in_f[4][DATA][8] ,
         \latches_in_f[4][DATA][7] , \latches_in_f[4][DATA][6] ,
         \latches_in_f[4][DATA][5] , \latches_in_f[4][DATA][4] ,
         \latches_in_f[4][DATA][3] , \latches_in_f[4][DATA][2] ,
         \latches_in_f[4][DATA][1] , \latches_in_f[4][DATA][0] ,
         \latches_in_f[3][REQ] , \latches_in_f[3][DATA][34] ,
         \latches_in_f[3][DATA][33] , \latches_in_f[3][DATA][32] ,
         \latches_in_f[3][DATA][31] , \latches_in_f[3][DATA][30] ,
         \latches_in_f[3][DATA][29] , \latches_in_f[3][DATA][28] ,
         \latches_in_f[3][DATA][27] , \latches_in_f[3][DATA][26] ,
         \latches_in_f[3][DATA][25] , \latches_in_f[3][DATA][24] ,
         \latches_in_f[3][DATA][23] , \latches_in_f[3][DATA][22] ,
         \latches_in_f[3][DATA][21] , \latches_in_f[3][DATA][20] ,
         \latches_in_f[3][DATA][19] , \latches_in_f[3][DATA][18] ,
         \latches_in_f[3][DATA][17] , \latches_in_f[3][DATA][16] ,
         \latches_in_f[3][DATA][15] , \latches_in_f[3][DATA][14] ,
         \latches_in_f[3][DATA][13] , \latches_in_f[3][DATA][12] ,
         \latches_in_f[3][DATA][11] , \latches_in_f[3][DATA][10] ,
         \latches_in_f[3][DATA][9] , \latches_in_f[3][DATA][8] ,
         \latches_in_f[3][DATA][7] , \latches_in_f[3][DATA][6] ,
         \latches_in_f[3][DATA][5] , \latches_in_f[3][DATA][4] ,
         \latches_in_f[3][DATA][3] , \latches_in_f[3][DATA][2] ,
         \latches_in_f[3][DATA][1] , \latches_in_f[3][DATA][0] ,
         \latches_in_f[2][REQ] , \latches_in_f[2][DATA][34] ,
         \latches_in_f[2][DATA][33] , \latches_in_f[2][DATA][32] ,
         \latches_in_f[2][DATA][31] , \latches_in_f[2][DATA][30] ,
         \latches_in_f[2][DATA][29] , \latches_in_f[2][DATA][28] ,
         \latches_in_f[2][DATA][27] , \latches_in_f[2][DATA][26] ,
         \latches_in_f[2][DATA][25] , \latches_in_f[2][DATA][24] ,
         \latches_in_f[2][DATA][23] , \latches_in_f[2][DATA][22] ,
         \latches_in_f[2][DATA][21] , \latches_in_f[2][DATA][20] ,
         \latches_in_f[2][DATA][19] , \latches_in_f[2][DATA][18] ,
         \latches_in_f[2][DATA][17] , \latches_in_f[2][DATA][16] ,
         \latches_in_f[2][DATA][15] , \latches_in_f[2][DATA][14] ,
         \latches_in_f[2][DATA][13] , \latches_in_f[2][DATA][12] ,
         \latches_in_f[2][DATA][11] , \latches_in_f[2][DATA][10] ,
         \latches_in_f[2][DATA][9] , \latches_in_f[2][DATA][8] ,
         \latches_in_f[2][DATA][7] , \latches_in_f[2][DATA][6] ,
         \latches_in_f[2][DATA][5] , \latches_in_f[2][DATA][4] ,
         \latches_in_f[2][DATA][3] , \latches_in_f[2][DATA][2] ,
         \latches_in_f[2][DATA][1] , \latches_in_f[2][DATA][0] ,
         \latches_in_f[1][REQ] , \latches_in_f[1][DATA][34] ,
         \latches_in_f[1][DATA][33] , \latches_in_f[1][DATA][32] ,
         \latches_in_f[1][DATA][31] , \latches_in_f[1][DATA][30] ,
         \latches_in_f[1][DATA][29] , \latches_in_f[1][DATA][28] ,
         \latches_in_f[1][DATA][27] , \latches_in_f[1][DATA][26] ,
         \latches_in_f[1][DATA][25] , \latches_in_f[1][DATA][24] ,
         \latches_in_f[1][DATA][23] , \latches_in_f[1][DATA][22] ,
         \latches_in_f[1][DATA][21] , \latches_in_f[1][DATA][20] ,
         \latches_in_f[1][DATA][19] , \latches_in_f[1][DATA][18] ,
         \latches_in_f[1][DATA][17] , \latches_in_f[1][DATA][16] ,
         \latches_in_f[1][DATA][15] , \latches_in_f[1][DATA][14] ,
         \latches_in_f[1][DATA][13] , \latches_in_f[1][DATA][12] ,
         \latches_in_f[1][DATA][11] , \latches_in_f[1][DATA][10] ,
         \latches_in_f[1][DATA][9] , \latches_in_f[1][DATA][8] ,
         \latches_in_f[1][DATA][7] , \latches_in_f[1][DATA][6] ,
         \latches_in_f[1][DATA][5] , \latches_in_f[1][DATA][4] ,
         \latches_in_f[1][DATA][3] , \latches_in_f[1][DATA][2] ,
         \latches_in_f[1][DATA][1] , \latches_in_f[1][DATA][0] ,
         \latches_in_f[0][REQ] , \latches_in_f[0][DATA][34] ,
         \latches_in_f[0][DATA][33] , \latches_in_f[0][DATA][32] ,
         \latches_in_f[0][DATA][31] , \latches_in_f[0][DATA][30] ,
         \latches_in_f[0][DATA][29] , \latches_in_f[0][DATA][28] ,
         \latches_in_f[0][DATA][27] , \latches_in_f[0][DATA][26] ,
         \latches_in_f[0][DATA][25] , \latches_in_f[0][DATA][24] ,
         \latches_in_f[0][DATA][23] , \latches_in_f[0][DATA][22] ,
         \latches_in_f[0][DATA][21] , \latches_in_f[0][DATA][20] ,
         \latches_in_f[0][DATA][19] , \latches_in_f[0][DATA][18] ,
         \latches_in_f[0][DATA][17] , \latches_in_f[0][DATA][16] ,
         \latches_in_f[0][DATA][15] , \latches_in_f[0][DATA][14] ,
         \latches_in_f[0][DATA][13] , \latches_in_f[0][DATA][12] ,
         \latches_in_f[0][DATA][11] , \latches_in_f[0][DATA][10] ,
         \latches_in_f[0][DATA][9] , \latches_in_f[0][DATA][8] ,
         \latches_in_f[0][DATA][7] , \latches_in_f[0][DATA][6] ,
         \latches_in_f[0][DATA][5] , \latches_in_f[0][DATA][4] ,
         \latches_in_f[0][DATA][3] , \latches_in_f[0][DATA][2] ,
         \latches_in_f[0][DATA][1] , \latches_in_f[0][DATA][0] ,
         \latches_in_b[4][ACK] , \latches_in_b[3][ACK] ,
         \latches_in_b[2][ACK] , \latches_in_b[1][ACK] ,
         \latches_in_b[0][ACK] , n1;

  crossbar_2 crossbar ( .preset(n1), .switch_sel({\switch_sel[4][4] , 
        \switch_sel[4][3] , \switch_sel[4][2] , \switch_sel[4][1] , 
        \switch_sel[4][0] , \switch_sel[3][4] , \switch_sel[3][3] , 
        \switch_sel[3][2] , \switch_sel[3][1] , \switch_sel[3][0] , 
        \switch_sel[2][4] , \switch_sel[2][3] , \switch_sel[2][2] , 
        \switch_sel[2][1] , \switch_sel[2][0] , \switch_sel[1][4] , 
        \switch_sel[1][3] , \switch_sel[1][2] , \switch_sel[1][1] , 
        \switch_sel[1][0] , \switch_sel[0][4] , \switch_sel[0][3] , 
        \switch_sel[0][2] , \switch_sel[0][1] , \switch_sel[0][0] }), 
        .chs_in_f({\chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] , 
        \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] , 
        \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] , 
        \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] , 
        \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] , 
        \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] , 
        \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] , 
        \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] , 
        \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] , 
        \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] , 
        \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] , 
        \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] , 
        \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] , 
        \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] , \chs_in_f[4][DATA][7] , 
        \chs_in_f[4][DATA][6] , \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] , 
        \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] , \chs_in_f[4][DATA][1] , 
        \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] , \chs_in_f[3][DATA][34] , 
        \chs_in_f[3][DATA][33] , \chs_in_f[3][DATA][32] , 
        \chs_in_f[3][DATA][31] , \chs_in_f[3][DATA][30] , 
        \chs_in_f[3][DATA][29] , \chs_in_f[3][DATA][28] , 
        \chs_in_f[3][DATA][27] , \chs_in_f[3][DATA][26] , 
        \chs_in_f[3][DATA][25] , \chs_in_f[3][DATA][24] , 
        \chs_in_f[3][DATA][23] , \chs_in_f[3][DATA][22] , 
        \chs_in_f[3][DATA][21] , \chs_in_f[3][DATA][20] , 
        \chs_in_f[3][DATA][19] , \chs_in_f[3][DATA][18] , 
        \chs_in_f[3][DATA][17] , \chs_in_f[3][DATA][16] , 
        \chs_in_f[3][DATA][15] , \chs_in_f[3][DATA][14] , 
        \chs_in_f[3][DATA][13] , \chs_in_f[3][DATA][12] , 
        \chs_in_f[3][DATA][11] , \chs_in_f[3][DATA][10] , 
        \chs_in_f[3][DATA][9] , \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] , 
        \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] , \chs_in_f[3][DATA][4] , 
        \chs_in_f[3][DATA][3] , \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] , 
        \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] , 
        \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] , 
        \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] , 
        \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] , 
        \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] , 
        \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] , 
        \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] , 
        \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] , 
        \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] , 
        \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] , 
        \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] , 
        \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] , 
        \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] , 
        \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] , \chs_in_f[2][DATA][7] , 
        \chs_in_f[2][DATA][6] , \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] , 
        \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] , \chs_in_f[2][DATA][1] , 
        \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] , \chs_in_f[1][DATA][34] , 
        \chs_in_f[1][DATA][33] , \chs_in_f[1][DATA][32] , 
        \chs_in_f[1][DATA][31] , \chs_in_f[1][DATA][30] , 
        \chs_in_f[1][DATA][29] , \chs_in_f[1][DATA][28] , 
        \chs_in_f[1][DATA][27] , \chs_in_f[1][DATA][26] , 
        \chs_in_f[1][DATA][25] , \chs_in_f[1][DATA][24] , 
        \chs_in_f[1][DATA][23] , \chs_in_f[1][DATA][22] , 
        \chs_in_f[1][DATA][21] , \chs_in_f[1][DATA][20] , 
        \chs_in_f[1][DATA][19] , \chs_in_f[1][DATA][18] , 
        \chs_in_f[1][DATA][17] , \chs_in_f[1][DATA][16] , 
        \chs_in_f[1][DATA][15] , \chs_in_f[1][DATA][14] , 
        \chs_in_f[1][DATA][13] , \chs_in_f[1][DATA][12] , 
        \chs_in_f[1][DATA][11] , \chs_in_f[1][DATA][10] , 
        \chs_in_f[1][DATA][9] , \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] , 
        \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] , \chs_in_f[1][DATA][4] , 
        \chs_in_f[1][DATA][3] , \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] , 
        \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] , 
        \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] , 
        \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] , 
        \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] , 
        \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] , 
        \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] , 
        \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] , 
        \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] , 
        \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] , 
        \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] , 
        \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] , 
        \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] , 
        \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] , 
        \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] , \chs_in_f[0][DATA][7] , 
        \chs_in_f[0][DATA][6] , \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] , 
        \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] , \chs_in_f[0][DATA][1] , 
        \chs_in_f[0][DATA][0] }), .chs_in_b({\chs_in_b[4][ACK] , 
        \chs_in_b[3][ACK] , \chs_in_b[2][ACK] , \chs_in_b[1][ACK] , 
        \chs_in_b[0][ACK] }), .chs_out_f({\latches_in_f[4][REQ] , 
        \latches_in_f[4][DATA][34] , \latches_in_f[4][DATA][33] , 
        \latches_in_f[4][DATA][32] , \latches_in_f[4][DATA][31] , 
        \latches_in_f[4][DATA][30] , \latches_in_f[4][DATA][29] , 
        \latches_in_f[4][DATA][28] , \latches_in_f[4][DATA][27] , 
        \latches_in_f[4][DATA][26] , \latches_in_f[4][DATA][25] , 
        \latches_in_f[4][DATA][24] , \latches_in_f[4][DATA][23] , 
        \latches_in_f[4][DATA][22] , \latches_in_f[4][DATA][21] , 
        \latches_in_f[4][DATA][20] , \latches_in_f[4][DATA][19] , 
        \latches_in_f[4][DATA][18] , \latches_in_f[4][DATA][17] , 
        \latches_in_f[4][DATA][16] , \latches_in_f[4][DATA][15] , 
        \latches_in_f[4][DATA][14] , \latches_in_f[4][DATA][13] , 
        \latches_in_f[4][DATA][12] , \latches_in_f[4][DATA][11] , 
        \latches_in_f[4][DATA][10] , \latches_in_f[4][DATA][9] , 
        \latches_in_f[4][DATA][8] , \latches_in_f[4][DATA][7] , 
        \latches_in_f[4][DATA][6] , \latches_in_f[4][DATA][5] , 
        \latches_in_f[4][DATA][4] , \latches_in_f[4][DATA][3] , 
        \latches_in_f[4][DATA][2] , \latches_in_f[4][DATA][1] , 
        \latches_in_f[4][DATA][0] , \latches_in_f[3][REQ] , 
        \latches_in_f[3][DATA][34] , \latches_in_f[3][DATA][33] , 
        \latches_in_f[3][DATA][32] , \latches_in_f[3][DATA][31] , 
        \latches_in_f[3][DATA][30] , \latches_in_f[3][DATA][29] , 
        \latches_in_f[3][DATA][28] , \latches_in_f[3][DATA][27] , 
        \latches_in_f[3][DATA][26] , \latches_in_f[3][DATA][25] , 
        \latches_in_f[3][DATA][24] , \latches_in_f[3][DATA][23] , 
        \latches_in_f[3][DATA][22] , \latches_in_f[3][DATA][21] , 
        \latches_in_f[3][DATA][20] , \latches_in_f[3][DATA][19] , 
        \latches_in_f[3][DATA][18] , \latches_in_f[3][DATA][17] , 
        \latches_in_f[3][DATA][16] , \latches_in_f[3][DATA][15] , 
        \latches_in_f[3][DATA][14] , \latches_in_f[3][DATA][13] , 
        \latches_in_f[3][DATA][12] , \latches_in_f[3][DATA][11] , 
        \latches_in_f[3][DATA][10] , \latches_in_f[3][DATA][9] , 
        \latches_in_f[3][DATA][8] , \latches_in_f[3][DATA][7] , 
        \latches_in_f[3][DATA][6] , \latches_in_f[3][DATA][5] , 
        \latches_in_f[3][DATA][4] , \latches_in_f[3][DATA][3] , 
        \latches_in_f[3][DATA][2] , \latches_in_f[3][DATA][1] , 
        \latches_in_f[3][DATA][0] , \latches_in_f[2][REQ] , 
        \latches_in_f[2][DATA][34] , \latches_in_f[2][DATA][33] , 
        \latches_in_f[2][DATA][32] , \latches_in_f[2][DATA][31] , 
        \latches_in_f[2][DATA][30] , \latches_in_f[2][DATA][29] , 
        \latches_in_f[2][DATA][28] , \latches_in_f[2][DATA][27] , 
        \latches_in_f[2][DATA][26] , \latches_in_f[2][DATA][25] , 
        \latches_in_f[2][DATA][24] , \latches_in_f[2][DATA][23] , 
        \latches_in_f[2][DATA][22] , \latches_in_f[2][DATA][21] , 
        \latches_in_f[2][DATA][20] , \latches_in_f[2][DATA][19] , 
        \latches_in_f[2][DATA][18] , \latches_in_f[2][DATA][17] , 
        \latches_in_f[2][DATA][16] , \latches_in_f[2][DATA][15] , 
        \latches_in_f[2][DATA][14] , \latches_in_f[2][DATA][13] , 
        \latches_in_f[2][DATA][12] , \latches_in_f[2][DATA][11] , 
        \latches_in_f[2][DATA][10] , \latches_in_f[2][DATA][9] , 
        \latches_in_f[2][DATA][8] , \latches_in_f[2][DATA][7] , 
        \latches_in_f[2][DATA][6] , \latches_in_f[2][DATA][5] , 
        \latches_in_f[2][DATA][4] , \latches_in_f[2][DATA][3] , 
        \latches_in_f[2][DATA][2] , \latches_in_f[2][DATA][1] , 
        \latches_in_f[2][DATA][0] , \latches_in_f[1][REQ] , 
        \latches_in_f[1][DATA][34] , \latches_in_f[1][DATA][33] , 
        \latches_in_f[1][DATA][32] , \latches_in_f[1][DATA][31] , 
        \latches_in_f[1][DATA][30] , \latches_in_f[1][DATA][29] , 
        \latches_in_f[1][DATA][28] , \latches_in_f[1][DATA][27] , 
        \latches_in_f[1][DATA][26] , \latches_in_f[1][DATA][25] , 
        \latches_in_f[1][DATA][24] , \latches_in_f[1][DATA][23] , 
        \latches_in_f[1][DATA][22] , \latches_in_f[1][DATA][21] , 
        \latches_in_f[1][DATA][20] , \latches_in_f[1][DATA][19] , 
        \latches_in_f[1][DATA][18] , \latches_in_f[1][DATA][17] , 
        \latches_in_f[1][DATA][16] , \latches_in_f[1][DATA][15] , 
        \latches_in_f[1][DATA][14] , \latches_in_f[1][DATA][13] , 
        \latches_in_f[1][DATA][12] , \latches_in_f[1][DATA][11] , 
        \latches_in_f[1][DATA][10] , \latches_in_f[1][DATA][9] , 
        \latches_in_f[1][DATA][8] , \latches_in_f[1][DATA][7] , 
        \latches_in_f[1][DATA][6] , \latches_in_f[1][DATA][5] , 
        \latches_in_f[1][DATA][4] , \latches_in_f[1][DATA][3] , 
        \latches_in_f[1][DATA][2] , \latches_in_f[1][DATA][1] , 
        \latches_in_f[1][DATA][0] , \latches_in_f[0][REQ] , 
        \latches_in_f[0][DATA][34] , \latches_in_f[0][DATA][33] , 
        \latches_in_f[0][DATA][32] , \latches_in_f[0][DATA][31] , 
        \latches_in_f[0][DATA][30] , \latches_in_f[0][DATA][29] , 
        \latches_in_f[0][DATA][28] , \latches_in_f[0][DATA][27] , 
        \latches_in_f[0][DATA][26] , \latches_in_f[0][DATA][25] , 
        \latches_in_f[0][DATA][24] , \latches_in_f[0][DATA][23] , 
        \latches_in_f[0][DATA][22] , \latches_in_f[0][DATA][21] , 
        \latches_in_f[0][DATA][20] , \latches_in_f[0][DATA][19] , 
        \latches_in_f[0][DATA][18] , \latches_in_f[0][DATA][17] , 
        \latches_in_f[0][DATA][16] , \latches_in_f[0][DATA][15] , 
        \latches_in_f[0][DATA][14] , \latches_in_f[0][DATA][13] , 
        \latches_in_f[0][DATA][12] , \latches_in_f[0][DATA][11] , 
        \latches_in_f[0][DATA][10] , \latches_in_f[0][DATA][9] , 
        \latches_in_f[0][DATA][8] , \latches_in_f[0][DATA][7] , 
        \latches_in_f[0][DATA][6] , \latches_in_f[0][DATA][5] , 
        \latches_in_f[0][DATA][4] , \latches_in_f[0][DATA][3] , 
        \latches_in_f[0][DATA][2] , \latches_in_f[0][DATA][1] , 
        \latches_in_f[0][DATA][0] }), .chs_out_b({\latches_in_b[4][ACK] , 
        \latches_in_b[3][ACK] , \latches_in_b[2][ACK] , \latches_in_b[1][ACK] , 
        \latches_in_b[0][ACK] }) );
  channel_latch_0_000000000_10 ch_latch_4 ( .preset(n1), .left_in({
        \latches_in_f[4][REQ] , \latches_in_f[4][DATA][34] , 
        \latches_in_f[4][DATA][33] , \latches_in_f[4][DATA][32] , 
        \latches_in_f[4][DATA][31] , \latches_in_f[4][DATA][30] , 
        \latches_in_f[4][DATA][29] , \latches_in_f[4][DATA][28] , 
        \latches_in_f[4][DATA][27] , \latches_in_f[4][DATA][26] , 
        \latches_in_f[4][DATA][25] , \latches_in_f[4][DATA][24] , 
        \latches_in_f[4][DATA][23] , \latches_in_f[4][DATA][22] , 
        \latches_in_f[4][DATA][21] , \latches_in_f[4][DATA][20] , 
        \latches_in_f[4][DATA][19] , \latches_in_f[4][DATA][18] , 
        \latches_in_f[4][DATA][17] , \latches_in_f[4][DATA][16] , 
        \latches_in_f[4][DATA][15] , \latches_in_f[4][DATA][14] , 
        \latches_in_f[4][DATA][13] , \latches_in_f[4][DATA][12] , 
        \latches_in_f[4][DATA][11] , \latches_in_f[4][DATA][10] , 
        \latches_in_f[4][DATA][9] , \latches_in_f[4][DATA][8] , 
        \latches_in_f[4][DATA][7] , \latches_in_f[4][DATA][6] , 
        \latches_in_f[4][DATA][5] , \latches_in_f[4][DATA][4] , 
        \latches_in_f[4][DATA][3] , \latches_in_f[4][DATA][2] , 
        \latches_in_f[4][DATA][1] , \latches_in_f[4][DATA][0] }), .left_out(
        \latches_in_b[4][ACK] ), .right_out({\latches_out_f[4][REQ] , 
        \latches_out_f[4][DATA][34] , \latches_out_f[4][DATA][33] , 
        \latches_out_f[4][DATA][32] , \latches_out_f[4][DATA][31] , 
        \latches_out_f[4][DATA][30] , \latches_out_f[4][DATA][29] , 
        \latches_out_f[4][DATA][28] , \latches_out_f[4][DATA][27] , 
        \latches_out_f[4][DATA][26] , \latches_out_f[4][DATA][25] , 
        \latches_out_f[4][DATA][24] , \latches_out_f[4][DATA][23] , 
        \latches_out_f[4][DATA][22] , \latches_out_f[4][DATA][21] , 
        \latches_out_f[4][DATA][20] , \latches_out_f[4][DATA][19] , 
        \latches_out_f[4][DATA][18] , \latches_out_f[4][DATA][17] , 
        \latches_out_f[4][DATA][16] , \latches_out_f[4][DATA][15] , 
        \latches_out_f[4][DATA][14] , \latches_out_f[4][DATA][13] , 
        \latches_out_f[4][DATA][12] , \latches_out_f[4][DATA][11] , 
        \latches_out_f[4][DATA][10] , \latches_out_f[4][DATA][9] , 
        \latches_out_f[4][DATA][8] , \latches_out_f[4][DATA][7] , 
        \latches_out_f[4][DATA][6] , \latches_out_f[4][DATA][5] , 
        \latches_out_f[4][DATA][4] , \latches_out_f[4][DATA][3] , 
        \latches_out_f[4][DATA][2] , \latches_out_f[4][DATA][1] , 
        \latches_out_f[4][DATA][0] }), .right_in(\latches_out_b[4][ACK] ) );
  channel_latch_0_000000000_9 ch_latch_3 ( .preset(n1), .left_in({
        \latches_in_f[3][REQ] , \latches_in_f[3][DATA][34] , 
        \latches_in_f[3][DATA][33] , \latches_in_f[3][DATA][32] , 
        \latches_in_f[3][DATA][31] , \latches_in_f[3][DATA][30] , 
        \latches_in_f[3][DATA][29] , \latches_in_f[3][DATA][28] , 
        \latches_in_f[3][DATA][27] , \latches_in_f[3][DATA][26] , 
        \latches_in_f[3][DATA][25] , \latches_in_f[3][DATA][24] , 
        \latches_in_f[3][DATA][23] , \latches_in_f[3][DATA][22] , 
        \latches_in_f[3][DATA][21] , \latches_in_f[3][DATA][20] , 
        \latches_in_f[3][DATA][19] , \latches_in_f[3][DATA][18] , 
        \latches_in_f[3][DATA][17] , \latches_in_f[3][DATA][16] , 
        \latches_in_f[3][DATA][15] , \latches_in_f[3][DATA][14] , 
        \latches_in_f[3][DATA][13] , \latches_in_f[3][DATA][12] , 
        \latches_in_f[3][DATA][11] , \latches_in_f[3][DATA][10] , 
        \latches_in_f[3][DATA][9] , \latches_in_f[3][DATA][8] , 
        \latches_in_f[3][DATA][7] , \latches_in_f[3][DATA][6] , 
        \latches_in_f[3][DATA][5] , \latches_in_f[3][DATA][4] , 
        \latches_in_f[3][DATA][3] , \latches_in_f[3][DATA][2] , 
        \latches_in_f[3][DATA][1] , \latches_in_f[3][DATA][0] }), .left_out(
        \latches_in_b[3][ACK] ), .right_out({\latches_out_f[3][REQ] , 
        \latches_out_f[3][DATA][34] , \latches_out_f[3][DATA][33] , 
        \latches_out_f[3][DATA][32] , \latches_out_f[3][DATA][31] , 
        \latches_out_f[3][DATA][30] , \latches_out_f[3][DATA][29] , 
        \latches_out_f[3][DATA][28] , \latches_out_f[3][DATA][27] , 
        \latches_out_f[3][DATA][26] , \latches_out_f[3][DATA][25] , 
        \latches_out_f[3][DATA][24] , \latches_out_f[3][DATA][23] , 
        \latches_out_f[3][DATA][22] , \latches_out_f[3][DATA][21] , 
        \latches_out_f[3][DATA][20] , \latches_out_f[3][DATA][19] , 
        \latches_out_f[3][DATA][18] , \latches_out_f[3][DATA][17] , 
        \latches_out_f[3][DATA][16] , \latches_out_f[3][DATA][15] , 
        \latches_out_f[3][DATA][14] , \latches_out_f[3][DATA][13] , 
        \latches_out_f[3][DATA][12] , \latches_out_f[3][DATA][11] , 
        \latches_out_f[3][DATA][10] , \latches_out_f[3][DATA][9] , 
        \latches_out_f[3][DATA][8] , \latches_out_f[3][DATA][7] , 
        \latches_out_f[3][DATA][6] , \latches_out_f[3][DATA][5] , 
        \latches_out_f[3][DATA][4] , \latches_out_f[3][DATA][3] , 
        \latches_out_f[3][DATA][2] , \latches_out_f[3][DATA][1] , 
        \latches_out_f[3][DATA][0] }), .right_in(\latches_out_b[3][ACK] ) );
  channel_latch_0_000000000_8 ch_latch_2 ( .preset(n1), .left_in({
        \latches_in_f[2][REQ] , \latches_in_f[2][DATA][34] , 
        \latches_in_f[2][DATA][33] , \latches_in_f[2][DATA][32] , 
        \latches_in_f[2][DATA][31] , \latches_in_f[2][DATA][30] , 
        \latches_in_f[2][DATA][29] , \latches_in_f[2][DATA][28] , 
        \latches_in_f[2][DATA][27] , \latches_in_f[2][DATA][26] , 
        \latches_in_f[2][DATA][25] , \latches_in_f[2][DATA][24] , 
        \latches_in_f[2][DATA][23] , \latches_in_f[2][DATA][22] , 
        \latches_in_f[2][DATA][21] , \latches_in_f[2][DATA][20] , 
        \latches_in_f[2][DATA][19] , \latches_in_f[2][DATA][18] , 
        \latches_in_f[2][DATA][17] , \latches_in_f[2][DATA][16] , 
        \latches_in_f[2][DATA][15] , \latches_in_f[2][DATA][14] , 
        \latches_in_f[2][DATA][13] , \latches_in_f[2][DATA][12] , 
        \latches_in_f[2][DATA][11] , \latches_in_f[2][DATA][10] , 
        \latches_in_f[2][DATA][9] , \latches_in_f[2][DATA][8] , 
        \latches_in_f[2][DATA][7] , \latches_in_f[2][DATA][6] , 
        \latches_in_f[2][DATA][5] , \latches_in_f[2][DATA][4] , 
        \latches_in_f[2][DATA][3] , \latches_in_f[2][DATA][2] , 
        \latches_in_f[2][DATA][1] , \latches_in_f[2][DATA][0] }), .left_out(
        \latches_in_b[2][ACK] ), .right_out({\latches_out_f[2][REQ] , 
        \latches_out_f[2][DATA][34] , \latches_out_f[2][DATA][33] , 
        \latches_out_f[2][DATA][32] , \latches_out_f[2][DATA][31] , 
        \latches_out_f[2][DATA][30] , \latches_out_f[2][DATA][29] , 
        \latches_out_f[2][DATA][28] , \latches_out_f[2][DATA][27] , 
        \latches_out_f[2][DATA][26] , \latches_out_f[2][DATA][25] , 
        \latches_out_f[2][DATA][24] , \latches_out_f[2][DATA][23] , 
        \latches_out_f[2][DATA][22] , \latches_out_f[2][DATA][21] , 
        \latches_out_f[2][DATA][20] , \latches_out_f[2][DATA][19] , 
        \latches_out_f[2][DATA][18] , \latches_out_f[2][DATA][17] , 
        \latches_out_f[2][DATA][16] , \latches_out_f[2][DATA][15] , 
        \latches_out_f[2][DATA][14] , \latches_out_f[2][DATA][13] , 
        \latches_out_f[2][DATA][12] , \latches_out_f[2][DATA][11] , 
        \latches_out_f[2][DATA][10] , \latches_out_f[2][DATA][9] , 
        \latches_out_f[2][DATA][8] , \latches_out_f[2][DATA][7] , 
        \latches_out_f[2][DATA][6] , \latches_out_f[2][DATA][5] , 
        \latches_out_f[2][DATA][4] , \latches_out_f[2][DATA][3] , 
        \latches_out_f[2][DATA][2] , \latches_out_f[2][DATA][1] , 
        \latches_out_f[2][DATA][0] }), .right_in(\latches_out_b[2][ACK] ) );
  channel_latch_0_000000000_7 ch_latch_1 ( .preset(n1), .left_in({
        \latches_in_f[1][REQ] , \latches_in_f[1][DATA][34] , 
        \latches_in_f[1][DATA][33] , \latches_in_f[1][DATA][32] , 
        \latches_in_f[1][DATA][31] , \latches_in_f[1][DATA][30] , 
        \latches_in_f[1][DATA][29] , \latches_in_f[1][DATA][28] , 
        \latches_in_f[1][DATA][27] , \latches_in_f[1][DATA][26] , 
        \latches_in_f[1][DATA][25] , \latches_in_f[1][DATA][24] , 
        \latches_in_f[1][DATA][23] , \latches_in_f[1][DATA][22] , 
        \latches_in_f[1][DATA][21] , \latches_in_f[1][DATA][20] , 
        \latches_in_f[1][DATA][19] , \latches_in_f[1][DATA][18] , 
        \latches_in_f[1][DATA][17] , \latches_in_f[1][DATA][16] , 
        \latches_in_f[1][DATA][15] , \latches_in_f[1][DATA][14] , 
        \latches_in_f[1][DATA][13] , \latches_in_f[1][DATA][12] , 
        \latches_in_f[1][DATA][11] , \latches_in_f[1][DATA][10] , 
        \latches_in_f[1][DATA][9] , \latches_in_f[1][DATA][8] , 
        \latches_in_f[1][DATA][7] , \latches_in_f[1][DATA][6] , 
        \latches_in_f[1][DATA][5] , \latches_in_f[1][DATA][4] , 
        \latches_in_f[1][DATA][3] , \latches_in_f[1][DATA][2] , 
        \latches_in_f[1][DATA][1] , \latches_in_f[1][DATA][0] }), .left_out(
        \latches_in_b[1][ACK] ), .right_out({\latches_out_f[1][REQ] , 
        \latches_out_f[1][DATA][34] , \latches_out_f[1][DATA][33] , 
        \latches_out_f[1][DATA][32] , \latches_out_f[1][DATA][31] , 
        \latches_out_f[1][DATA][30] , \latches_out_f[1][DATA][29] , 
        \latches_out_f[1][DATA][28] , \latches_out_f[1][DATA][27] , 
        \latches_out_f[1][DATA][26] , \latches_out_f[1][DATA][25] , 
        \latches_out_f[1][DATA][24] , \latches_out_f[1][DATA][23] , 
        \latches_out_f[1][DATA][22] , \latches_out_f[1][DATA][21] , 
        \latches_out_f[1][DATA][20] , \latches_out_f[1][DATA][19] , 
        \latches_out_f[1][DATA][18] , \latches_out_f[1][DATA][17] , 
        \latches_out_f[1][DATA][16] , \latches_out_f[1][DATA][15] , 
        \latches_out_f[1][DATA][14] , \latches_out_f[1][DATA][13] , 
        \latches_out_f[1][DATA][12] , \latches_out_f[1][DATA][11] , 
        \latches_out_f[1][DATA][10] , \latches_out_f[1][DATA][9] , 
        \latches_out_f[1][DATA][8] , \latches_out_f[1][DATA][7] , 
        \latches_out_f[1][DATA][6] , \latches_out_f[1][DATA][5] , 
        \latches_out_f[1][DATA][4] , \latches_out_f[1][DATA][3] , 
        \latches_out_f[1][DATA][2] , \latches_out_f[1][DATA][1] , 
        \latches_out_f[1][DATA][0] }), .right_in(\latches_out_b[1][ACK] ) );
  channel_latch_0_000000000_6 ch_latch_0 ( .preset(n1), .left_in({
        \latches_in_f[0][REQ] , \latches_in_f[0][DATA][34] , 
        \latches_in_f[0][DATA][33] , \latches_in_f[0][DATA][32] , 
        \latches_in_f[0][DATA][31] , \latches_in_f[0][DATA][30] , 
        \latches_in_f[0][DATA][29] , \latches_in_f[0][DATA][28] , 
        \latches_in_f[0][DATA][27] , \latches_in_f[0][DATA][26] , 
        \latches_in_f[0][DATA][25] , \latches_in_f[0][DATA][24] , 
        \latches_in_f[0][DATA][23] , \latches_in_f[0][DATA][22] , 
        \latches_in_f[0][DATA][21] , \latches_in_f[0][DATA][20] , 
        \latches_in_f[0][DATA][19] , \latches_in_f[0][DATA][18] , 
        \latches_in_f[0][DATA][17] , \latches_in_f[0][DATA][16] , 
        \latches_in_f[0][DATA][15] , \latches_in_f[0][DATA][14] , 
        \latches_in_f[0][DATA][13] , \latches_in_f[0][DATA][12] , 
        \latches_in_f[0][DATA][11] , \latches_in_f[0][DATA][10] , 
        \latches_in_f[0][DATA][9] , \latches_in_f[0][DATA][8] , 
        \latches_in_f[0][DATA][7] , \latches_in_f[0][DATA][6] , 
        \latches_in_f[0][DATA][5] , \latches_in_f[0][DATA][4] , 
        \latches_in_f[0][DATA][3] , \latches_in_f[0][DATA][2] , 
        \latches_in_f[0][DATA][1] , \latches_in_f[0][DATA][0] }), .left_out(
        \latches_in_b[0][ACK] ), .right_out({\latches_out_f[0][REQ] , 
        \latches_out_f[0][DATA][34] , \latches_out_f[0][DATA][33] , 
        \latches_out_f[0][DATA][32] , \latches_out_f[0][DATA][31] , 
        \latches_out_f[0][DATA][30] , \latches_out_f[0][DATA][29] , 
        \latches_out_f[0][DATA][28] , \latches_out_f[0][DATA][27] , 
        \latches_out_f[0][DATA][26] , \latches_out_f[0][DATA][25] , 
        \latches_out_f[0][DATA][24] , \latches_out_f[0][DATA][23] , 
        \latches_out_f[0][DATA][22] , \latches_out_f[0][DATA][21] , 
        \latches_out_f[0][DATA][20] , \latches_out_f[0][DATA][19] , 
        \latches_out_f[0][DATA][18] , \latches_out_f[0][DATA][17] , 
        \latches_out_f[0][DATA][16] , \latches_out_f[0][DATA][15] , 
        \latches_out_f[0][DATA][14] , \latches_out_f[0][DATA][13] , 
        \latches_out_f[0][DATA][12] , \latches_out_f[0][DATA][11] , 
        \latches_out_f[0][DATA][10] , \latches_out_f[0][DATA][9] , 
        \latches_out_f[0][DATA][8] , \latches_out_f[0][DATA][7] , 
        \latches_out_f[0][DATA][6] , \latches_out_f[0][DATA][5] , 
        \latches_out_f[0][DATA][4] , \latches_out_f[0][DATA][3] , 
        \latches_out_f[0][DATA][2] , \latches_out_f[0][DATA][1] , 
        \latches_out_f[0][DATA][0] }), .right_in(\latches_out_b[0][ACK] ) );
  HS65_LS_BFX9 U1 ( .A(preset), .Z(n1) );
endmodule


module noc_switch_2 ( preset, .north_in_f({\north_in_f[REQ] , 
        \north_in_f[DATA][34] , \north_in_f[DATA][33] , \north_in_f[DATA][32] , 
        \north_in_f[DATA][31] , \north_in_f[DATA][30] , \north_in_f[DATA][29] , 
        \north_in_f[DATA][28] , \north_in_f[DATA][27] , \north_in_f[DATA][26] , 
        \north_in_f[DATA][25] , \north_in_f[DATA][24] , \north_in_f[DATA][23] , 
        \north_in_f[DATA][22] , \north_in_f[DATA][21] , \north_in_f[DATA][20] , 
        \north_in_f[DATA][19] , \north_in_f[DATA][18] , \north_in_f[DATA][17] , 
        \north_in_f[DATA][16] , \north_in_f[DATA][15] , \north_in_f[DATA][14] , 
        \north_in_f[DATA][13] , \north_in_f[DATA][12] , \north_in_f[DATA][11] , 
        \north_in_f[DATA][10] , \north_in_f[DATA][9] , \north_in_f[DATA][8] , 
        \north_in_f[DATA][7] , \north_in_f[DATA][6] , \north_in_f[DATA][5] , 
        \north_in_f[DATA][4] , \north_in_f[DATA][3] , \north_in_f[DATA][2] , 
        \north_in_f[DATA][1] , \north_in_f[DATA][0] }), .north_in_b(
        \north_in_b[ACK] ), .east_in_f({\east_in_f[REQ] , 
        \east_in_f[DATA][34] , \east_in_f[DATA][33] , \east_in_f[DATA][32] , 
        \east_in_f[DATA][31] , \east_in_f[DATA][30] , \east_in_f[DATA][29] , 
        \east_in_f[DATA][28] , \east_in_f[DATA][27] , \east_in_f[DATA][26] , 
        \east_in_f[DATA][25] , \east_in_f[DATA][24] , \east_in_f[DATA][23] , 
        \east_in_f[DATA][22] , \east_in_f[DATA][21] , \east_in_f[DATA][20] , 
        \east_in_f[DATA][19] , \east_in_f[DATA][18] , \east_in_f[DATA][17] , 
        \east_in_f[DATA][16] , \east_in_f[DATA][15] , \east_in_f[DATA][14] , 
        \east_in_f[DATA][13] , \east_in_f[DATA][12] , \east_in_f[DATA][11] , 
        \east_in_f[DATA][10] , \east_in_f[DATA][9] , \east_in_f[DATA][8] , 
        \east_in_f[DATA][7] , \east_in_f[DATA][6] , \east_in_f[DATA][5] , 
        \east_in_f[DATA][4] , \east_in_f[DATA][3] , \east_in_f[DATA][2] , 
        \east_in_f[DATA][1] , \east_in_f[DATA][0] }), .east_in_b(
        \east_in_b[ACK] ), .south_in_f({\south_in_f[REQ] , 
        \south_in_f[DATA][34] , \south_in_f[DATA][33] , \south_in_f[DATA][32] , 
        \south_in_f[DATA][31] , \south_in_f[DATA][30] , \south_in_f[DATA][29] , 
        \south_in_f[DATA][28] , \south_in_f[DATA][27] , \south_in_f[DATA][26] , 
        \south_in_f[DATA][25] , \south_in_f[DATA][24] , \south_in_f[DATA][23] , 
        \south_in_f[DATA][22] , \south_in_f[DATA][21] , \south_in_f[DATA][20] , 
        \south_in_f[DATA][19] , \south_in_f[DATA][18] , \south_in_f[DATA][17] , 
        \south_in_f[DATA][16] , \south_in_f[DATA][15] , \south_in_f[DATA][14] , 
        \south_in_f[DATA][13] , \south_in_f[DATA][12] , \south_in_f[DATA][11] , 
        \south_in_f[DATA][10] , \south_in_f[DATA][9] , \south_in_f[DATA][8] , 
        \south_in_f[DATA][7] , \south_in_f[DATA][6] , \south_in_f[DATA][5] , 
        \south_in_f[DATA][4] , \south_in_f[DATA][3] , \south_in_f[DATA][2] , 
        \south_in_f[DATA][1] , \south_in_f[DATA][0] }), .south_in_b(
        \south_in_b[ACK] ), .west_in_f({\west_in_f[REQ] , 
        \west_in_f[DATA][34] , \west_in_f[DATA][33] , \west_in_f[DATA][32] , 
        \west_in_f[DATA][31] , \west_in_f[DATA][30] , \west_in_f[DATA][29] , 
        \west_in_f[DATA][28] , \west_in_f[DATA][27] , \west_in_f[DATA][26] , 
        \west_in_f[DATA][25] , \west_in_f[DATA][24] , \west_in_f[DATA][23] , 
        \west_in_f[DATA][22] , \west_in_f[DATA][21] , \west_in_f[DATA][20] , 
        \west_in_f[DATA][19] , \west_in_f[DATA][18] , \west_in_f[DATA][17] , 
        \west_in_f[DATA][16] , \west_in_f[DATA][15] , \west_in_f[DATA][14] , 
        \west_in_f[DATA][13] , \west_in_f[DATA][12] , \west_in_f[DATA][11] , 
        \west_in_f[DATA][10] , \west_in_f[DATA][9] , \west_in_f[DATA][8] , 
        \west_in_f[DATA][7] , \west_in_f[DATA][6] , \west_in_f[DATA][5] , 
        \west_in_f[DATA][4] , \west_in_f[DATA][3] , \west_in_f[DATA][2] , 
        \west_in_f[DATA][1] , \west_in_f[DATA][0] }), .west_in_b(
        \west_in_b[ACK] ), .resource_in_f({\resource_in_f[REQ] , 
        \resource_in_f[DATA][34] , \resource_in_f[DATA][33] , 
        \resource_in_f[DATA][32] , \resource_in_f[DATA][31] , 
        \resource_in_f[DATA][30] , \resource_in_f[DATA][29] , 
        \resource_in_f[DATA][28] , \resource_in_f[DATA][27] , 
        \resource_in_f[DATA][26] , \resource_in_f[DATA][25] , 
        \resource_in_f[DATA][24] , \resource_in_f[DATA][23] , 
        \resource_in_f[DATA][22] , \resource_in_f[DATA][21] , 
        \resource_in_f[DATA][20] , \resource_in_f[DATA][19] , 
        \resource_in_f[DATA][18] , \resource_in_f[DATA][17] , 
        \resource_in_f[DATA][16] , \resource_in_f[DATA][15] , 
        \resource_in_f[DATA][14] , \resource_in_f[DATA][13] , 
        \resource_in_f[DATA][12] , \resource_in_f[DATA][11] , 
        \resource_in_f[DATA][10] , \resource_in_f[DATA][9] , 
        \resource_in_f[DATA][8] , \resource_in_f[DATA][7] , 
        \resource_in_f[DATA][6] , \resource_in_f[DATA][5] , 
        \resource_in_f[DATA][4] , \resource_in_f[DATA][3] , 
        \resource_in_f[DATA][2] , \resource_in_f[DATA][1] , 
        \resource_in_f[DATA][0] }), .resource_in_b(\resource_in_b[ACK] ), 
    .north_out_f({\north_out_f[REQ] , \north_out_f[DATA][34] , 
        \north_out_f[DATA][33] , \north_out_f[DATA][32] , 
        \north_out_f[DATA][31] , \north_out_f[DATA][30] , 
        \north_out_f[DATA][29] , \north_out_f[DATA][28] , 
        \north_out_f[DATA][27] , \north_out_f[DATA][26] , 
        \north_out_f[DATA][25] , \north_out_f[DATA][24] , 
        \north_out_f[DATA][23] , \north_out_f[DATA][22] , 
        \north_out_f[DATA][21] , \north_out_f[DATA][20] , 
        \north_out_f[DATA][19] , \north_out_f[DATA][18] , 
        \north_out_f[DATA][17] , \north_out_f[DATA][16] , 
        \north_out_f[DATA][15] , \north_out_f[DATA][14] , 
        \north_out_f[DATA][13] , \north_out_f[DATA][12] , 
        \north_out_f[DATA][11] , \north_out_f[DATA][10] , 
        \north_out_f[DATA][9] , \north_out_f[DATA][8] , \north_out_f[DATA][7] , 
        \north_out_f[DATA][6] , \north_out_f[DATA][5] , \north_out_f[DATA][4] , 
        \north_out_f[DATA][3] , \north_out_f[DATA][2] , \north_out_f[DATA][1] , 
        \north_out_f[DATA][0] }), .north_out_b(\north_out_b[ACK] ), 
    .east_out_f({\east_out_f[REQ] , \east_out_f[DATA][34] , 
        \east_out_f[DATA][33] , \east_out_f[DATA][32] , \east_out_f[DATA][31] , 
        \east_out_f[DATA][30] , \east_out_f[DATA][29] , \east_out_f[DATA][28] , 
        \east_out_f[DATA][27] , \east_out_f[DATA][26] , \east_out_f[DATA][25] , 
        \east_out_f[DATA][24] , \east_out_f[DATA][23] , \east_out_f[DATA][22] , 
        \east_out_f[DATA][21] , \east_out_f[DATA][20] , \east_out_f[DATA][19] , 
        \east_out_f[DATA][18] , \east_out_f[DATA][17] , \east_out_f[DATA][16] , 
        \east_out_f[DATA][15] , \east_out_f[DATA][14] , \east_out_f[DATA][13] , 
        \east_out_f[DATA][12] , \east_out_f[DATA][11] , \east_out_f[DATA][10] , 
        \east_out_f[DATA][9] , \east_out_f[DATA][8] , \east_out_f[DATA][7] , 
        \east_out_f[DATA][6] , \east_out_f[DATA][5] , \east_out_f[DATA][4] , 
        \east_out_f[DATA][3] , \east_out_f[DATA][2] , \east_out_f[DATA][1] , 
        \east_out_f[DATA][0] }), .east_out_b(\east_out_b[ACK] ), 
    .south_out_f({\south_out_f[REQ] , \south_out_f[DATA][34] , 
        \south_out_f[DATA][33] , \south_out_f[DATA][32] , 
        \south_out_f[DATA][31] , \south_out_f[DATA][30] , 
        \south_out_f[DATA][29] , \south_out_f[DATA][28] , 
        \south_out_f[DATA][27] , \south_out_f[DATA][26] , 
        \south_out_f[DATA][25] , \south_out_f[DATA][24] , 
        \south_out_f[DATA][23] , \south_out_f[DATA][22] , 
        \south_out_f[DATA][21] , \south_out_f[DATA][20] , 
        \south_out_f[DATA][19] , \south_out_f[DATA][18] , 
        \south_out_f[DATA][17] , \south_out_f[DATA][16] , 
        \south_out_f[DATA][15] , \south_out_f[DATA][14] , 
        \south_out_f[DATA][13] , \south_out_f[DATA][12] , 
        \south_out_f[DATA][11] , \south_out_f[DATA][10] , 
        \south_out_f[DATA][9] , \south_out_f[DATA][8] , \south_out_f[DATA][7] , 
        \south_out_f[DATA][6] , \south_out_f[DATA][5] , \south_out_f[DATA][4] , 
        \south_out_f[DATA][3] , \south_out_f[DATA][2] , \south_out_f[DATA][1] , 
        \south_out_f[DATA][0] }), .south_out_b(\south_out_b[ACK] ), 
    .west_out_f({\west_out_f[REQ] , \west_out_f[DATA][34] , 
        \west_out_f[DATA][33] , \west_out_f[DATA][32] , \west_out_f[DATA][31] , 
        \west_out_f[DATA][30] , \west_out_f[DATA][29] , \west_out_f[DATA][28] , 
        \west_out_f[DATA][27] , \west_out_f[DATA][26] , \west_out_f[DATA][25] , 
        \west_out_f[DATA][24] , \west_out_f[DATA][23] , \west_out_f[DATA][22] , 
        \west_out_f[DATA][21] , \west_out_f[DATA][20] , \west_out_f[DATA][19] , 
        \west_out_f[DATA][18] , \west_out_f[DATA][17] , \west_out_f[DATA][16] , 
        \west_out_f[DATA][15] , \west_out_f[DATA][14] , \west_out_f[DATA][13] , 
        \west_out_f[DATA][12] , \west_out_f[DATA][11] , \west_out_f[DATA][10] , 
        \west_out_f[DATA][9] , \west_out_f[DATA][8] , \west_out_f[DATA][7] , 
        \west_out_f[DATA][6] , \west_out_f[DATA][5] , \west_out_f[DATA][4] , 
        \west_out_f[DATA][3] , \west_out_f[DATA][2] , \west_out_f[DATA][1] , 
        \west_out_f[DATA][0] }), .west_out_b(\west_out_b[ACK] ), 
    .resource_out_f({\resource_out_f[REQ] , \resource_out_f[DATA][34] , 
        \resource_out_f[DATA][33] , \resource_out_f[DATA][32] , 
        \resource_out_f[DATA][31] , \resource_out_f[DATA][30] , 
        \resource_out_f[DATA][29] , \resource_out_f[DATA][28] , 
        \resource_out_f[DATA][27] , \resource_out_f[DATA][26] , 
        \resource_out_f[DATA][25] , \resource_out_f[DATA][24] , 
        \resource_out_f[DATA][23] , \resource_out_f[DATA][22] , 
        \resource_out_f[DATA][21] , \resource_out_f[DATA][20] , 
        \resource_out_f[DATA][19] , \resource_out_f[DATA][18] , 
        \resource_out_f[DATA][17] , \resource_out_f[DATA][16] , 
        \resource_out_f[DATA][15] , \resource_out_f[DATA][14] , 
        \resource_out_f[DATA][13] , \resource_out_f[DATA][12] , 
        \resource_out_f[DATA][11] , \resource_out_f[DATA][10] , 
        \resource_out_f[DATA][9] , \resource_out_f[DATA][8] , 
        \resource_out_f[DATA][7] , \resource_out_f[DATA][6] , 
        \resource_out_f[DATA][5] , \resource_out_f[DATA][4] , 
        \resource_out_f[DATA][3] , \resource_out_f[DATA][2] , 
        \resource_out_f[DATA][1] , \resource_out_f[DATA][0] }), 
    .resource_out_b(\resource_out_b[ACK] ) );
  input preset, \north_in_f[REQ] , \north_in_f[DATA][34] ,
         \north_in_f[DATA][33] , \north_in_f[DATA][32] ,
         \north_in_f[DATA][31] , \north_in_f[DATA][30] ,
         \north_in_f[DATA][29] , \north_in_f[DATA][28] ,
         \north_in_f[DATA][27] , \north_in_f[DATA][26] ,
         \north_in_f[DATA][25] , \north_in_f[DATA][24] ,
         \north_in_f[DATA][23] , \north_in_f[DATA][22] ,
         \north_in_f[DATA][21] , \north_in_f[DATA][20] ,
         \north_in_f[DATA][19] , \north_in_f[DATA][18] ,
         \north_in_f[DATA][17] , \north_in_f[DATA][16] ,
         \north_in_f[DATA][15] , \north_in_f[DATA][14] ,
         \north_in_f[DATA][13] , \north_in_f[DATA][12] ,
         \north_in_f[DATA][11] , \north_in_f[DATA][10] , \north_in_f[DATA][9] ,
         \north_in_f[DATA][8] , \north_in_f[DATA][7] , \north_in_f[DATA][6] ,
         \north_in_f[DATA][5] , \north_in_f[DATA][4] , \north_in_f[DATA][3] ,
         \north_in_f[DATA][2] , \north_in_f[DATA][1] , \north_in_f[DATA][0] ,
         \east_in_f[REQ] , \east_in_f[DATA][34] , \east_in_f[DATA][33] ,
         \east_in_f[DATA][32] , \east_in_f[DATA][31] , \east_in_f[DATA][30] ,
         \east_in_f[DATA][29] , \east_in_f[DATA][28] , \east_in_f[DATA][27] ,
         \east_in_f[DATA][26] , \east_in_f[DATA][25] , \east_in_f[DATA][24] ,
         \east_in_f[DATA][23] , \east_in_f[DATA][22] , \east_in_f[DATA][21] ,
         \east_in_f[DATA][20] , \east_in_f[DATA][19] , \east_in_f[DATA][18] ,
         \east_in_f[DATA][17] , \east_in_f[DATA][16] , \east_in_f[DATA][15] ,
         \east_in_f[DATA][14] , \east_in_f[DATA][13] , \east_in_f[DATA][12] ,
         \east_in_f[DATA][11] , \east_in_f[DATA][10] , \east_in_f[DATA][9] ,
         \east_in_f[DATA][8] , \east_in_f[DATA][7] , \east_in_f[DATA][6] ,
         \east_in_f[DATA][5] , \east_in_f[DATA][4] , \east_in_f[DATA][3] ,
         \east_in_f[DATA][2] , \east_in_f[DATA][1] , \east_in_f[DATA][0] ,
         \south_in_f[REQ] , \south_in_f[DATA][34] , \south_in_f[DATA][33] ,
         \south_in_f[DATA][32] , \south_in_f[DATA][31] ,
         \south_in_f[DATA][30] , \south_in_f[DATA][29] ,
         \south_in_f[DATA][28] , \south_in_f[DATA][27] ,
         \south_in_f[DATA][26] , \south_in_f[DATA][25] ,
         \south_in_f[DATA][24] , \south_in_f[DATA][23] ,
         \south_in_f[DATA][22] , \south_in_f[DATA][21] ,
         \south_in_f[DATA][20] , \south_in_f[DATA][19] ,
         \south_in_f[DATA][18] , \south_in_f[DATA][17] ,
         \south_in_f[DATA][16] , \south_in_f[DATA][15] ,
         \south_in_f[DATA][14] , \south_in_f[DATA][13] ,
         \south_in_f[DATA][12] , \south_in_f[DATA][11] ,
         \south_in_f[DATA][10] , \south_in_f[DATA][9] , \south_in_f[DATA][8] ,
         \south_in_f[DATA][7] , \south_in_f[DATA][6] , \south_in_f[DATA][5] ,
         \south_in_f[DATA][4] , \south_in_f[DATA][3] , \south_in_f[DATA][2] ,
         \south_in_f[DATA][1] , \south_in_f[DATA][0] , \west_in_f[REQ] ,
         \west_in_f[DATA][34] , \west_in_f[DATA][33] , \west_in_f[DATA][32] ,
         \west_in_f[DATA][31] , \west_in_f[DATA][30] , \west_in_f[DATA][29] ,
         \west_in_f[DATA][28] , \west_in_f[DATA][27] , \west_in_f[DATA][26] ,
         \west_in_f[DATA][25] , \west_in_f[DATA][24] , \west_in_f[DATA][23] ,
         \west_in_f[DATA][22] , \west_in_f[DATA][21] , \west_in_f[DATA][20] ,
         \west_in_f[DATA][19] , \west_in_f[DATA][18] , \west_in_f[DATA][17] ,
         \west_in_f[DATA][16] , \west_in_f[DATA][15] , \west_in_f[DATA][14] ,
         \west_in_f[DATA][13] , \west_in_f[DATA][12] , \west_in_f[DATA][11] ,
         \west_in_f[DATA][10] , \west_in_f[DATA][9] , \west_in_f[DATA][8] ,
         \west_in_f[DATA][7] , \west_in_f[DATA][6] , \west_in_f[DATA][5] ,
         \west_in_f[DATA][4] , \west_in_f[DATA][3] , \west_in_f[DATA][2] ,
         \west_in_f[DATA][1] , \west_in_f[DATA][0] , \resource_in_f[REQ] ,
         \resource_in_f[DATA][34] , \resource_in_f[DATA][33] ,
         \resource_in_f[DATA][32] , \resource_in_f[DATA][31] ,
         \resource_in_f[DATA][30] , \resource_in_f[DATA][29] ,
         \resource_in_f[DATA][28] , \resource_in_f[DATA][27] ,
         \resource_in_f[DATA][26] , \resource_in_f[DATA][25] ,
         \resource_in_f[DATA][24] , \resource_in_f[DATA][23] ,
         \resource_in_f[DATA][22] , \resource_in_f[DATA][21] ,
         \resource_in_f[DATA][20] , \resource_in_f[DATA][19] ,
         \resource_in_f[DATA][18] , \resource_in_f[DATA][17] ,
         \resource_in_f[DATA][16] , \resource_in_f[DATA][15] ,
         \resource_in_f[DATA][14] , \resource_in_f[DATA][13] ,
         \resource_in_f[DATA][12] , \resource_in_f[DATA][11] ,
         \resource_in_f[DATA][10] , \resource_in_f[DATA][9] ,
         \resource_in_f[DATA][8] , \resource_in_f[DATA][7] ,
         \resource_in_f[DATA][6] , \resource_in_f[DATA][5] ,
         \resource_in_f[DATA][4] , \resource_in_f[DATA][3] ,
         \resource_in_f[DATA][2] , \resource_in_f[DATA][1] ,
         \resource_in_f[DATA][0] , \north_out_b[ACK] , \east_out_b[ACK] ,
         \south_out_b[ACK] , \west_out_b[ACK] , \resource_out_b[ACK] ;
  output \north_in_b[ACK] , \east_in_b[ACK] , \south_in_b[ACK] ,
         \west_in_b[ACK] , \resource_in_b[ACK] , \north_out_f[REQ] ,
         \north_out_f[DATA][34] , \north_out_f[DATA][33] ,
         \north_out_f[DATA][32] , \north_out_f[DATA][31] ,
         \north_out_f[DATA][30] , \north_out_f[DATA][29] ,
         \north_out_f[DATA][28] , \north_out_f[DATA][27] ,
         \north_out_f[DATA][26] , \north_out_f[DATA][25] ,
         \north_out_f[DATA][24] , \north_out_f[DATA][23] ,
         \north_out_f[DATA][22] , \north_out_f[DATA][21] ,
         \north_out_f[DATA][20] , \north_out_f[DATA][19] ,
         \north_out_f[DATA][18] , \north_out_f[DATA][17] ,
         \north_out_f[DATA][16] , \north_out_f[DATA][15] ,
         \north_out_f[DATA][14] , \north_out_f[DATA][13] ,
         \north_out_f[DATA][12] , \north_out_f[DATA][11] ,
         \north_out_f[DATA][10] , \north_out_f[DATA][9] ,
         \north_out_f[DATA][8] , \north_out_f[DATA][7] ,
         \north_out_f[DATA][6] , \north_out_f[DATA][5] ,
         \north_out_f[DATA][4] , \north_out_f[DATA][3] ,
         \north_out_f[DATA][2] , \north_out_f[DATA][1] ,
         \north_out_f[DATA][0] , \east_out_f[REQ] , \east_out_f[DATA][34] ,
         \east_out_f[DATA][33] , \east_out_f[DATA][32] ,
         \east_out_f[DATA][31] , \east_out_f[DATA][30] ,
         \east_out_f[DATA][29] , \east_out_f[DATA][28] ,
         \east_out_f[DATA][27] , \east_out_f[DATA][26] ,
         \east_out_f[DATA][25] , \east_out_f[DATA][24] ,
         \east_out_f[DATA][23] , \east_out_f[DATA][22] ,
         \east_out_f[DATA][21] , \east_out_f[DATA][20] ,
         \east_out_f[DATA][19] , \east_out_f[DATA][18] ,
         \east_out_f[DATA][17] , \east_out_f[DATA][16] ,
         \east_out_f[DATA][15] , \east_out_f[DATA][14] ,
         \east_out_f[DATA][13] , \east_out_f[DATA][12] ,
         \east_out_f[DATA][11] , \east_out_f[DATA][10] , \east_out_f[DATA][9] ,
         \east_out_f[DATA][8] , \east_out_f[DATA][7] , \east_out_f[DATA][6] ,
         \east_out_f[DATA][5] , \east_out_f[DATA][4] , \east_out_f[DATA][3] ,
         \east_out_f[DATA][2] , \east_out_f[DATA][1] , \east_out_f[DATA][0] ,
         \south_out_f[REQ] , \south_out_f[DATA][34] , \south_out_f[DATA][33] ,
         \south_out_f[DATA][32] , \south_out_f[DATA][31] ,
         \south_out_f[DATA][30] , \south_out_f[DATA][29] ,
         \south_out_f[DATA][28] , \south_out_f[DATA][27] ,
         \south_out_f[DATA][26] , \south_out_f[DATA][25] ,
         \south_out_f[DATA][24] , \south_out_f[DATA][23] ,
         \south_out_f[DATA][22] , \south_out_f[DATA][21] ,
         \south_out_f[DATA][20] , \south_out_f[DATA][19] ,
         \south_out_f[DATA][18] , \south_out_f[DATA][17] ,
         \south_out_f[DATA][16] , \south_out_f[DATA][15] ,
         \south_out_f[DATA][14] , \south_out_f[DATA][13] ,
         \south_out_f[DATA][12] , \south_out_f[DATA][11] ,
         \south_out_f[DATA][10] , \south_out_f[DATA][9] ,
         \south_out_f[DATA][8] , \south_out_f[DATA][7] ,
         \south_out_f[DATA][6] , \south_out_f[DATA][5] ,
         \south_out_f[DATA][4] , \south_out_f[DATA][3] ,
         \south_out_f[DATA][2] , \south_out_f[DATA][1] ,
         \south_out_f[DATA][0] , \west_out_f[REQ] , \west_out_f[DATA][34] ,
         \west_out_f[DATA][33] , \west_out_f[DATA][32] ,
         \west_out_f[DATA][31] , \west_out_f[DATA][30] ,
         \west_out_f[DATA][29] , \west_out_f[DATA][28] ,
         \west_out_f[DATA][27] , \west_out_f[DATA][26] ,
         \west_out_f[DATA][25] , \west_out_f[DATA][24] ,
         \west_out_f[DATA][23] , \west_out_f[DATA][22] ,
         \west_out_f[DATA][21] , \west_out_f[DATA][20] ,
         \west_out_f[DATA][19] , \west_out_f[DATA][18] ,
         \west_out_f[DATA][17] , \west_out_f[DATA][16] ,
         \west_out_f[DATA][15] , \west_out_f[DATA][14] ,
         \west_out_f[DATA][13] , \west_out_f[DATA][12] ,
         \west_out_f[DATA][11] , \west_out_f[DATA][10] , \west_out_f[DATA][9] ,
         \west_out_f[DATA][8] , \west_out_f[DATA][7] , \west_out_f[DATA][6] ,
         \west_out_f[DATA][5] , \west_out_f[DATA][4] , \west_out_f[DATA][3] ,
         \west_out_f[DATA][2] , \west_out_f[DATA][1] , \west_out_f[DATA][0] ,
         \resource_out_f[REQ] , \resource_out_f[DATA][34] ,
         \resource_out_f[DATA][33] , \resource_out_f[DATA][32] ,
         \resource_out_f[DATA][31] , \resource_out_f[DATA][30] ,
         \resource_out_f[DATA][29] , \resource_out_f[DATA][28] ,
         \resource_out_f[DATA][27] , \resource_out_f[DATA][26] ,
         \resource_out_f[DATA][25] , \resource_out_f[DATA][24] ,
         \resource_out_f[DATA][23] , \resource_out_f[DATA][22] ,
         \resource_out_f[DATA][21] , \resource_out_f[DATA][20] ,
         \resource_out_f[DATA][19] , \resource_out_f[DATA][18] ,
         \resource_out_f[DATA][17] , \resource_out_f[DATA][16] ,
         \resource_out_f[DATA][15] , \resource_out_f[DATA][14] ,
         \resource_out_f[DATA][13] , \resource_out_f[DATA][12] ,
         \resource_out_f[DATA][11] , \resource_out_f[DATA][10] ,
         \resource_out_f[DATA][9] , \resource_out_f[DATA][8] ,
         \resource_out_f[DATA][7] , \resource_out_f[DATA][6] ,
         \resource_out_f[DATA][5] , \resource_out_f[DATA][4] ,
         \resource_out_f[DATA][3] , \resource_out_f[DATA][2] ,
         \resource_out_f[DATA][1] , \resource_out_f[DATA][0] ;
  wire   \north_hpu_f[REQ] , \north_hpu_f[DATA][34] , \north_hpu_f[DATA][33] ,
         \north_hpu_f[DATA][32] , \north_hpu_f[DATA][31] ,
         \north_hpu_f[DATA][30] , \north_hpu_f[DATA][29] ,
         \north_hpu_f[DATA][28] , \north_hpu_f[DATA][27] ,
         \north_hpu_f[DATA][26] , \north_hpu_f[DATA][25] ,
         \north_hpu_f[DATA][24] , \north_hpu_f[DATA][23] ,
         \north_hpu_f[DATA][22] , \north_hpu_f[DATA][21] ,
         \north_hpu_f[DATA][20] , \north_hpu_f[DATA][19] ,
         \north_hpu_f[DATA][18] , \north_hpu_f[DATA][17] ,
         \north_hpu_f[DATA][16] , \north_hpu_f[DATA][15] ,
         \north_hpu_f[DATA][14] , \north_hpu_f[DATA][13] ,
         \north_hpu_f[DATA][12] , \north_hpu_f[DATA][11] ,
         \north_hpu_f[DATA][10] , \north_hpu_f[DATA][9] ,
         \north_hpu_f[DATA][8] , \north_hpu_f[DATA][7] ,
         \north_hpu_f[DATA][6] , \north_hpu_f[DATA][5] ,
         \north_hpu_f[DATA][4] , \north_hpu_f[DATA][3] ,
         \north_hpu_f[DATA][2] , \north_hpu_f[DATA][1] ,
         \north_hpu_f[DATA][0] , \north_hpu_b[ACK] , \south_hpu_f[REQ] ,
         \south_hpu_f[DATA][34] , \south_hpu_f[DATA][33] ,
         \south_hpu_f[DATA][32] , \south_hpu_f[DATA][31] ,
         \south_hpu_f[DATA][30] , \south_hpu_f[DATA][29] ,
         \south_hpu_f[DATA][28] , \south_hpu_f[DATA][27] ,
         \south_hpu_f[DATA][26] , \south_hpu_f[DATA][25] ,
         \south_hpu_f[DATA][24] , \south_hpu_f[DATA][23] ,
         \south_hpu_f[DATA][22] , \south_hpu_f[DATA][21] ,
         \south_hpu_f[DATA][20] , \south_hpu_f[DATA][19] ,
         \south_hpu_f[DATA][18] , \south_hpu_f[DATA][17] ,
         \south_hpu_f[DATA][16] , \south_hpu_f[DATA][15] ,
         \south_hpu_f[DATA][14] , \south_hpu_f[DATA][13] ,
         \south_hpu_f[DATA][12] , \south_hpu_f[DATA][11] ,
         \south_hpu_f[DATA][10] , \south_hpu_f[DATA][9] ,
         \south_hpu_f[DATA][8] , \south_hpu_f[DATA][7] ,
         \south_hpu_f[DATA][6] , \south_hpu_f[DATA][5] ,
         \south_hpu_f[DATA][4] , \south_hpu_f[DATA][3] ,
         \south_hpu_f[DATA][2] , \south_hpu_f[DATA][1] ,
         \south_hpu_f[DATA][0] , \south_hpu_b[ACK] , \east_hpu_f[REQ] ,
         \east_hpu_f[DATA][34] , \east_hpu_f[DATA][33] ,
         \east_hpu_f[DATA][32] , \east_hpu_f[DATA][31] ,
         \east_hpu_f[DATA][30] , \east_hpu_f[DATA][29] ,
         \east_hpu_f[DATA][28] , \east_hpu_f[DATA][27] ,
         \east_hpu_f[DATA][26] , \east_hpu_f[DATA][25] ,
         \east_hpu_f[DATA][24] , \east_hpu_f[DATA][23] ,
         \east_hpu_f[DATA][22] , \east_hpu_f[DATA][21] ,
         \east_hpu_f[DATA][20] , \east_hpu_f[DATA][19] ,
         \east_hpu_f[DATA][18] , \east_hpu_f[DATA][17] ,
         \east_hpu_f[DATA][16] , \east_hpu_f[DATA][15] ,
         \east_hpu_f[DATA][14] , \east_hpu_f[DATA][13] ,
         \east_hpu_f[DATA][12] , \east_hpu_f[DATA][11] ,
         \east_hpu_f[DATA][10] , \east_hpu_f[DATA][9] , \east_hpu_f[DATA][8] ,
         \east_hpu_f[DATA][7] , \east_hpu_f[DATA][6] , \east_hpu_f[DATA][5] ,
         \east_hpu_f[DATA][4] , \east_hpu_f[DATA][3] , \east_hpu_f[DATA][2] ,
         \east_hpu_f[DATA][1] , \east_hpu_f[DATA][0] , \east_hpu_b[ACK] ,
         \west_hpu_f[REQ] , \west_hpu_f[DATA][34] , \west_hpu_f[DATA][33] ,
         \west_hpu_f[DATA][32] , \west_hpu_f[DATA][31] ,
         \west_hpu_f[DATA][30] , \west_hpu_f[DATA][29] ,
         \west_hpu_f[DATA][28] , \west_hpu_f[DATA][27] ,
         \west_hpu_f[DATA][26] , \west_hpu_f[DATA][25] ,
         \west_hpu_f[DATA][24] , \west_hpu_f[DATA][23] ,
         \west_hpu_f[DATA][22] , \west_hpu_f[DATA][21] ,
         \west_hpu_f[DATA][20] , \west_hpu_f[DATA][19] ,
         \west_hpu_f[DATA][18] , \west_hpu_f[DATA][17] ,
         \west_hpu_f[DATA][16] , \west_hpu_f[DATA][15] ,
         \west_hpu_f[DATA][14] , \west_hpu_f[DATA][13] ,
         \west_hpu_f[DATA][12] , \west_hpu_f[DATA][11] ,
         \west_hpu_f[DATA][10] , \west_hpu_f[DATA][9] , \west_hpu_f[DATA][8] ,
         \west_hpu_f[DATA][7] , \west_hpu_f[DATA][6] , \west_hpu_f[DATA][5] ,
         \west_hpu_f[DATA][4] , \west_hpu_f[DATA][3] , \west_hpu_f[DATA][2] ,
         \west_hpu_f[DATA][1] , \west_hpu_f[DATA][0] , \west_hpu_b[ACK] ,
         \resource_hpu_f[REQ] , \resource_hpu_f[DATA][34] ,
         \resource_hpu_f[DATA][33] , \resource_hpu_f[DATA][32] ,
         \resource_hpu_f[DATA][31] , \resource_hpu_f[DATA][30] ,
         \resource_hpu_f[DATA][29] , \resource_hpu_f[DATA][28] ,
         \resource_hpu_f[DATA][27] , \resource_hpu_f[DATA][26] ,
         \resource_hpu_f[DATA][25] , \resource_hpu_f[DATA][24] ,
         \resource_hpu_f[DATA][23] , \resource_hpu_f[DATA][22] ,
         \resource_hpu_f[DATA][21] , \resource_hpu_f[DATA][20] ,
         \resource_hpu_f[DATA][19] , \resource_hpu_f[DATA][18] ,
         \resource_hpu_f[DATA][17] , \resource_hpu_f[DATA][16] ,
         \resource_hpu_f[DATA][15] , \resource_hpu_f[DATA][14] ,
         \resource_hpu_f[DATA][13] , \resource_hpu_f[DATA][12] ,
         \resource_hpu_f[DATA][11] , \resource_hpu_f[DATA][10] ,
         \resource_hpu_f[DATA][9] , \resource_hpu_f[DATA][8] ,
         \resource_hpu_f[DATA][7] , \resource_hpu_f[DATA][6] ,
         \resource_hpu_f[DATA][5] , \resource_hpu_f[DATA][4] ,
         \resource_hpu_f[DATA][3] , \resource_hpu_f[DATA][2] ,
         \resource_hpu_f[DATA][1] , \resource_hpu_f[DATA][0] ,
         \resource_hpu_b[ACK] , \chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] ,
         \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] ,
         \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] ,
         \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] ,
         \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] ,
         \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] ,
         \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] ,
         \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] ,
         \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] ,
         \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] ,
         \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] ,
         \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] ,
         \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] ,
         \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] ,
         \chs_in_f[4][DATA][7] , \chs_in_f[4][DATA][6] ,
         \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] ,
         \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] ,
         \chs_in_f[4][DATA][1] , \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] ,
         \chs_in_f[3][DATA][34] , \chs_in_f[3][DATA][33] ,
         \chs_in_f[3][DATA][32] , \chs_in_f[3][DATA][31] ,
         \chs_in_f[3][DATA][30] , \chs_in_f[3][DATA][29] ,
         \chs_in_f[3][DATA][28] , \chs_in_f[3][DATA][27] ,
         \chs_in_f[3][DATA][26] , \chs_in_f[3][DATA][25] ,
         \chs_in_f[3][DATA][24] , \chs_in_f[3][DATA][23] ,
         \chs_in_f[3][DATA][22] , \chs_in_f[3][DATA][21] ,
         \chs_in_f[3][DATA][20] , \chs_in_f[3][DATA][19] ,
         \chs_in_f[3][DATA][18] , \chs_in_f[3][DATA][17] ,
         \chs_in_f[3][DATA][16] , \chs_in_f[3][DATA][15] ,
         \chs_in_f[3][DATA][14] , \chs_in_f[3][DATA][13] ,
         \chs_in_f[3][DATA][12] , \chs_in_f[3][DATA][11] ,
         \chs_in_f[3][DATA][10] , \chs_in_f[3][DATA][9] ,
         \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] ,
         \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] ,
         \chs_in_f[3][DATA][4] , \chs_in_f[3][DATA][3] ,
         \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] ,
         \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] ,
         \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] ,
         \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] ,
         \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] ,
         \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] ,
         \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] ,
         \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] ,
         \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] ,
         \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] ,
         \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] ,
         \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] ,
         \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] ,
         \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] ,
         \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] ,
         \chs_in_f[2][DATA][7] , \chs_in_f[2][DATA][6] ,
         \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] ,
         \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] ,
         \chs_in_f[2][DATA][1] , \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] ,
         \chs_in_f[1][DATA][34] , \chs_in_f[1][DATA][33] ,
         \chs_in_f[1][DATA][32] , \chs_in_f[1][DATA][31] ,
         \chs_in_f[1][DATA][30] , \chs_in_f[1][DATA][29] ,
         \chs_in_f[1][DATA][28] , \chs_in_f[1][DATA][27] ,
         \chs_in_f[1][DATA][26] , \chs_in_f[1][DATA][25] ,
         \chs_in_f[1][DATA][24] , \chs_in_f[1][DATA][23] ,
         \chs_in_f[1][DATA][22] , \chs_in_f[1][DATA][21] ,
         \chs_in_f[1][DATA][20] , \chs_in_f[1][DATA][19] ,
         \chs_in_f[1][DATA][18] , \chs_in_f[1][DATA][17] ,
         \chs_in_f[1][DATA][16] , \chs_in_f[1][DATA][15] ,
         \chs_in_f[1][DATA][14] , \chs_in_f[1][DATA][13] ,
         \chs_in_f[1][DATA][12] , \chs_in_f[1][DATA][11] ,
         \chs_in_f[1][DATA][10] , \chs_in_f[1][DATA][9] ,
         \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] ,
         \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] ,
         \chs_in_f[1][DATA][4] , \chs_in_f[1][DATA][3] ,
         \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] ,
         \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] ,
         \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] ,
         \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] ,
         \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] ,
         \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] ,
         \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] ,
         \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] ,
         \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] ,
         \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] ,
         \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] ,
         \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] ,
         \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] ,
         \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] ,
         \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] ,
         \chs_in_f[0][DATA][7] , \chs_in_f[0][DATA][6] ,
         \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] ,
         \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] ,
         \chs_in_f[0][DATA][1] , \chs_in_f[0][DATA][0] , \chs_in_b[4][ACK] ,
         \chs_in_b[3][ACK] , \chs_in_b[2][ACK] , \chs_in_b[1][ACK] ,
         \chs_in_b[0][ACK] , \switch_sel[4][4] , \switch_sel[4][3] ,
         \switch_sel[4][2] , \switch_sel[4][1] , \switch_sel[4][0] ,
         \switch_sel[3][4] , \switch_sel[3][3] , \switch_sel[3][2] ,
         \switch_sel[3][1] , \switch_sel[3][0] , \switch_sel[2][4] ,
         \switch_sel[2][3] , \switch_sel[2][2] , \switch_sel[2][1] ,
         \switch_sel[2][0] , \switch_sel[1][4] , \switch_sel[1][3] ,
         \switch_sel[1][2] , \switch_sel[1][1] , \switch_sel[1][0] ,
         \switch_sel[0][4] , \switch_sel[0][3] , \switch_sel[0][2] ,
         \switch_sel[0][1] , \switch_sel[0][0] , n2, n3;

  channel_latch_1_xxxxxxxxx_30 north_in_latch ( .preset(n3), .left_in({
        \north_in_f[REQ] , \north_in_f[DATA][34] , \north_in_f[DATA][33] , 
        \north_in_f[DATA][32] , \north_in_f[DATA][31] , \north_in_f[DATA][30] , 
        \north_in_f[DATA][29] , \north_in_f[DATA][28] , \north_in_f[DATA][27] , 
        \north_in_f[DATA][26] , \north_in_f[DATA][25] , \north_in_f[DATA][24] , 
        \north_in_f[DATA][23] , \north_in_f[DATA][22] , \north_in_f[DATA][21] , 
        \north_in_f[DATA][20] , \north_in_f[DATA][19] , \north_in_f[DATA][18] , 
        \north_in_f[DATA][17] , \north_in_f[DATA][16] , \north_in_f[DATA][15] , 
        \north_in_f[DATA][14] , \north_in_f[DATA][13] , \north_in_f[DATA][12] , 
        \north_in_f[DATA][11] , \north_in_f[DATA][10] , \north_in_f[DATA][9] , 
        \north_in_f[DATA][8] , \north_in_f[DATA][7] , \north_in_f[DATA][6] , 
        \north_in_f[DATA][5] , \north_in_f[DATA][4] , \north_in_f[DATA][3] , 
        \north_in_f[DATA][2] , \north_in_f[DATA][1] , \north_in_f[DATA][0] }), 
        .left_out(\north_in_b[ACK] ), .right_out({\north_hpu_f[REQ] , 
        \north_hpu_f[DATA][34] , \north_hpu_f[DATA][33] , 
        \north_hpu_f[DATA][32] , \north_hpu_f[DATA][31] , 
        \north_hpu_f[DATA][30] , \north_hpu_f[DATA][29] , 
        \north_hpu_f[DATA][28] , \north_hpu_f[DATA][27] , 
        \north_hpu_f[DATA][26] , \north_hpu_f[DATA][25] , 
        \north_hpu_f[DATA][24] , \north_hpu_f[DATA][23] , 
        \north_hpu_f[DATA][22] , \north_hpu_f[DATA][21] , 
        \north_hpu_f[DATA][20] , \north_hpu_f[DATA][19] , 
        \north_hpu_f[DATA][18] , \north_hpu_f[DATA][17] , 
        \north_hpu_f[DATA][16] , \north_hpu_f[DATA][15] , 
        \north_hpu_f[DATA][14] , \north_hpu_f[DATA][13] , 
        \north_hpu_f[DATA][12] , \north_hpu_f[DATA][11] , 
        \north_hpu_f[DATA][10] , \north_hpu_f[DATA][9] , 
        \north_hpu_f[DATA][8] , \north_hpu_f[DATA][7] , \north_hpu_f[DATA][6] , 
        \north_hpu_f[DATA][5] , \north_hpu_f[DATA][4] , \north_hpu_f[DATA][3] , 
        \north_hpu_f[DATA][2] , \north_hpu_f[DATA][1] , \north_hpu_f[DATA][0] }), .right_in(\north_hpu_b[ACK] ) );
  channel_latch_1_xxxxxxxxx_29 south_in_latch ( .preset(n3), .left_in({
        \south_in_f[REQ] , \south_in_f[DATA][34] , \south_in_f[DATA][33] , 
        \south_in_f[DATA][32] , \south_in_f[DATA][31] , \south_in_f[DATA][30] , 
        \south_in_f[DATA][29] , \south_in_f[DATA][28] , \south_in_f[DATA][27] , 
        \south_in_f[DATA][26] , \south_in_f[DATA][25] , \south_in_f[DATA][24] , 
        \south_in_f[DATA][23] , \south_in_f[DATA][22] , \south_in_f[DATA][21] , 
        \south_in_f[DATA][20] , \south_in_f[DATA][19] , \south_in_f[DATA][18] , 
        \south_in_f[DATA][17] , \south_in_f[DATA][16] , \south_in_f[DATA][15] , 
        \south_in_f[DATA][14] , \south_in_f[DATA][13] , \south_in_f[DATA][12] , 
        \south_in_f[DATA][11] , \south_in_f[DATA][10] , \south_in_f[DATA][9] , 
        \south_in_f[DATA][8] , \south_in_f[DATA][7] , \south_in_f[DATA][6] , 
        \south_in_f[DATA][5] , \south_in_f[DATA][4] , \south_in_f[DATA][3] , 
        \south_in_f[DATA][2] , \south_in_f[DATA][1] , \south_in_f[DATA][0] }), 
        .left_out(\south_in_b[ACK] ), .right_out({\south_hpu_f[REQ] , 
        \south_hpu_f[DATA][34] , \south_hpu_f[DATA][33] , 
        \south_hpu_f[DATA][32] , \south_hpu_f[DATA][31] , 
        \south_hpu_f[DATA][30] , \south_hpu_f[DATA][29] , 
        \south_hpu_f[DATA][28] , \south_hpu_f[DATA][27] , 
        \south_hpu_f[DATA][26] , \south_hpu_f[DATA][25] , 
        \south_hpu_f[DATA][24] , \south_hpu_f[DATA][23] , 
        \south_hpu_f[DATA][22] , \south_hpu_f[DATA][21] , 
        \south_hpu_f[DATA][20] , \south_hpu_f[DATA][19] , 
        \south_hpu_f[DATA][18] , \south_hpu_f[DATA][17] , 
        \south_hpu_f[DATA][16] , \south_hpu_f[DATA][15] , 
        \south_hpu_f[DATA][14] , \south_hpu_f[DATA][13] , 
        \south_hpu_f[DATA][12] , \south_hpu_f[DATA][11] , 
        \south_hpu_f[DATA][10] , \south_hpu_f[DATA][9] , 
        \south_hpu_f[DATA][8] , \south_hpu_f[DATA][7] , \south_hpu_f[DATA][6] , 
        \south_hpu_f[DATA][5] , \south_hpu_f[DATA][4] , \south_hpu_f[DATA][3] , 
        \south_hpu_f[DATA][2] , \south_hpu_f[DATA][1] , \south_hpu_f[DATA][0] }), .right_in(\south_hpu_b[ACK] ) );
  channel_latch_1_xxxxxxxxx_28 east_in_latch ( .preset(n3), .left_in({
        \east_in_f[REQ] , \east_in_f[DATA][34] , \east_in_f[DATA][33] , 
        \east_in_f[DATA][32] , \east_in_f[DATA][31] , \east_in_f[DATA][30] , 
        \east_in_f[DATA][29] , \east_in_f[DATA][28] , \east_in_f[DATA][27] , 
        \east_in_f[DATA][26] , \east_in_f[DATA][25] , \east_in_f[DATA][24] , 
        \east_in_f[DATA][23] , \east_in_f[DATA][22] , \east_in_f[DATA][21] , 
        \east_in_f[DATA][20] , \east_in_f[DATA][19] , \east_in_f[DATA][18] , 
        \east_in_f[DATA][17] , \east_in_f[DATA][16] , \east_in_f[DATA][15] , 
        \east_in_f[DATA][14] , \east_in_f[DATA][13] , \east_in_f[DATA][12] , 
        \east_in_f[DATA][11] , \east_in_f[DATA][10] , \east_in_f[DATA][9] , 
        \east_in_f[DATA][8] , \east_in_f[DATA][7] , \east_in_f[DATA][6] , 
        \east_in_f[DATA][5] , \east_in_f[DATA][4] , \east_in_f[DATA][3] , 
        \east_in_f[DATA][2] , \east_in_f[DATA][1] , \east_in_f[DATA][0] }), 
        .left_out(\east_in_b[ACK] ), .right_out({\east_hpu_f[REQ] , 
        \east_hpu_f[DATA][34] , \east_hpu_f[DATA][33] , \east_hpu_f[DATA][32] , 
        \east_hpu_f[DATA][31] , \east_hpu_f[DATA][30] , \east_hpu_f[DATA][29] , 
        \east_hpu_f[DATA][28] , \east_hpu_f[DATA][27] , \east_hpu_f[DATA][26] , 
        \east_hpu_f[DATA][25] , \east_hpu_f[DATA][24] , \east_hpu_f[DATA][23] , 
        \east_hpu_f[DATA][22] , \east_hpu_f[DATA][21] , \east_hpu_f[DATA][20] , 
        \east_hpu_f[DATA][19] , \east_hpu_f[DATA][18] , \east_hpu_f[DATA][17] , 
        \east_hpu_f[DATA][16] , \east_hpu_f[DATA][15] , \east_hpu_f[DATA][14] , 
        \east_hpu_f[DATA][13] , \east_hpu_f[DATA][12] , \east_hpu_f[DATA][11] , 
        \east_hpu_f[DATA][10] , \east_hpu_f[DATA][9] , \east_hpu_f[DATA][8] , 
        \east_hpu_f[DATA][7] , \east_hpu_f[DATA][6] , \east_hpu_f[DATA][5] , 
        \east_hpu_f[DATA][4] , \east_hpu_f[DATA][3] , \east_hpu_f[DATA][2] , 
        \east_hpu_f[DATA][1] , \east_hpu_f[DATA][0] }), .right_in(
        \east_hpu_b[ACK] ) );
  channel_latch_1_xxxxxxxxx_27 west_in_latch ( .preset(n3), .left_in({
        \west_in_f[REQ] , \west_in_f[DATA][34] , \west_in_f[DATA][33] , 
        \west_in_f[DATA][32] , \west_in_f[DATA][31] , \west_in_f[DATA][30] , 
        \west_in_f[DATA][29] , \west_in_f[DATA][28] , \west_in_f[DATA][27] , 
        \west_in_f[DATA][26] , \west_in_f[DATA][25] , \west_in_f[DATA][24] , 
        \west_in_f[DATA][23] , \west_in_f[DATA][22] , \west_in_f[DATA][21] , 
        \west_in_f[DATA][20] , \west_in_f[DATA][19] , \west_in_f[DATA][18] , 
        \west_in_f[DATA][17] , \west_in_f[DATA][16] , \west_in_f[DATA][15] , 
        \west_in_f[DATA][14] , \west_in_f[DATA][13] , \west_in_f[DATA][12] , 
        \west_in_f[DATA][11] , \west_in_f[DATA][10] , \west_in_f[DATA][9] , 
        \west_in_f[DATA][8] , \west_in_f[DATA][7] , \west_in_f[DATA][6] , 
        \west_in_f[DATA][5] , \west_in_f[DATA][4] , \west_in_f[DATA][3] , 
        \west_in_f[DATA][2] , \west_in_f[DATA][1] , \west_in_f[DATA][0] }), 
        .left_out(\west_in_b[ACK] ), .right_out({\west_hpu_f[REQ] , 
        \west_hpu_f[DATA][34] , \west_hpu_f[DATA][33] , \west_hpu_f[DATA][32] , 
        \west_hpu_f[DATA][31] , \west_hpu_f[DATA][30] , \west_hpu_f[DATA][29] , 
        \west_hpu_f[DATA][28] , \west_hpu_f[DATA][27] , \west_hpu_f[DATA][26] , 
        \west_hpu_f[DATA][25] , \west_hpu_f[DATA][24] , \west_hpu_f[DATA][23] , 
        \west_hpu_f[DATA][22] , \west_hpu_f[DATA][21] , \west_hpu_f[DATA][20] , 
        \west_hpu_f[DATA][19] , \west_hpu_f[DATA][18] , \west_hpu_f[DATA][17] , 
        \west_hpu_f[DATA][16] , \west_hpu_f[DATA][15] , \west_hpu_f[DATA][14] , 
        \west_hpu_f[DATA][13] , \west_hpu_f[DATA][12] , \west_hpu_f[DATA][11] , 
        \west_hpu_f[DATA][10] , \west_hpu_f[DATA][9] , \west_hpu_f[DATA][8] , 
        \west_hpu_f[DATA][7] , \west_hpu_f[DATA][6] , \west_hpu_f[DATA][5] , 
        \west_hpu_f[DATA][4] , \west_hpu_f[DATA][3] , \west_hpu_f[DATA][2] , 
        \west_hpu_f[DATA][1] , \west_hpu_f[DATA][0] }), .right_in(
        \west_hpu_b[ACK] ) );
  channel_latch_1_xxxxxxxxx_26 resource_in_latch ( .preset(n3), .left_in({
        \resource_in_f[REQ] , \resource_in_f[DATA][34] , 
        \resource_in_f[DATA][33] , \resource_in_f[DATA][32] , 
        \resource_in_f[DATA][31] , \resource_in_f[DATA][30] , 
        \resource_in_f[DATA][29] , \resource_in_f[DATA][28] , 
        \resource_in_f[DATA][27] , \resource_in_f[DATA][26] , 
        \resource_in_f[DATA][25] , \resource_in_f[DATA][24] , 
        \resource_in_f[DATA][23] , \resource_in_f[DATA][22] , 
        \resource_in_f[DATA][21] , \resource_in_f[DATA][20] , 
        \resource_in_f[DATA][19] , \resource_in_f[DATA][18] , 
        \resource_in_f[DATA][17] , \resource_in_f[DATA][16] , 
        \resource_in_f[DATA][15] , \resource_in_f[DATA][14] , 
        \resource_in_f[DATA][13] , \resource_in_f[DATA][12] , 
        \resource_in_f[DATA][11] , \resource_in_f[DATA][10] , 
        \resource_in_f[DATA][9] , \resource_in_f[DATA][8] , 
        \resource_in_f[DATA][7] , \resource_in_f[DATA][6] , 
        \resource_in_f[DATA][5] , \resource_in_f[DATA][4] , 
        \resource_in_f[DATA][3] , \resource_in_f[DATA][2] , 
        \resource_in_f[DATA][1] , \resource_in_f[DATA][0] }), .left_out(
        \resource_in_b[ACK] ), .right_out({\resource_hpu_f[REQ] , 
        \resource_hpu_f[DATA][34] , \resource_hpu_f[DATA][33] , 
        \resource_hpu_f[DATA][32] , \resource_hpu_f[DATA][31] , 
        \resource_hpu_f[DATA][30] , \resource_hpu_f[DATA][29] , 
        \resource_hpu_f[DATA][28] , \resource_hpu_f[DATA][27] , 
        \resource_hpu_f[DATA][26] , \resource_hpu_f[DATA][25] , 
        \resource_hpu_f[DATA][24] , \resource_hpu_f[DATA][23] , 
        \resource_hpu_f[DATA][22] , \resource_hpu_f[DATA][21] , 
        \resource_hpu_f[DATA][20] , \resource_hpu_f[DATA][19] , 
        \resource_hpu_f[DATA][18] , \resource_hpu_f[DATA][17] , 
        \resource_hpu_f[DATA][16] , \resource_hpu_f[DATA][15] , 
        \resource_hpu_f[DATA][14] , \resource_hpu_f[DATA][13] , 
        \resource_hpu_f[DATA][12] , \resource_hpu_f[DATA][11] , 
        \resource_hpu_f[DATA][10] , \resource_hpu_f[DATA][9] , 
        \resource_hpu_f[DATA][8] , \resource_hpu_f[DATA][7] , 
        \resource_hpu_f[DATA][6] , \resource_hpu_f[DATA][5] , 
        \resource_hpu_f[DATA][4] , \resource_hpu_f[DATA][3] , 
        \resource_hpu_f[DATA][2] , \resource_hpu_f[DATA][1] , 
        \resource_hpu_f[DATA][0] }), .right_in(\resource_hpu_b[ACK] ) );
  hpu_0_0_2 north_hpu ( .preset(n2), .chan_in_f({\north_hpu_f[REQ] , 
        \north_hpu_f[DATA][34] , \north_hpu_f[DATA][33] , 
        \north_hpu_f[DATA][32] , \north_hpu_f[DATA][31] , 
        \north_hpu_f[DATA][30] , \north_hpu_f[DATA][29] , 
        \north_hpu_f[DATA][28] , \north_hpu_f[DATA][27] , 
        \north_hpu_f[DATA][26] , \north_hpu_f[DATA][25] , 
        \north_hpu_f[DATA][24] , \north_hpu_f[DATA][23] , 
        \north_hpu_f[DATA][22] , \north_hpu_f[DATA][21] , 
        \north_hpu_f[DATA][20] , \north_hpu_f[DATA][19] , 
        \north_hpu_f[DATA][18] , \north_hpu_f[DATA][17] , 
        \north_hpu_f[DATA][16] , \north_hpu_f[DATA][15] , 
        \north_hpu_f[DATA][14] , \north_hpu_f[DATA][13] , 
        \north_hpu_f[DATA][12] , \north_hpu_f[DATA][11] , 
        \north_hpu_f[DATA][10] , \north_hpu_f[DATA][9] , 
        \north_hpu_f[DATA][8] , \north_hpu_f[DATA][7] , \north_hpu_f[DATA][6] , 
        \north_hpu_f[DATA][5] , \north_hpu_f[DATA][4] , \north_hpu_f[DATA][3] , 
        \north_hpu_f[DATA][2] , \north_hpu_f[DATA][1] , \north_hpu_f[DATA][0] }), .chan_in_b(\north_hpu_b[ACK] ), .chan_out_f({\chs_in_f[0][REQ] , 
        \chs_in_f[0][DATA][34] , \chs_in_f[0][DATA][33] , 
        \chs_in_f[0][DATA][32] , \chs_in_f[0][DATA][31] , 
        \chs_in_f[0][DATA][30] , \chs_in_f[0][DATA][29] , 
        \chs_in_f[0][DATA][28] , \chs_in_f[0][DATA][27] , 
        \chs_in_f[0][DATA][26] , \chs_in_f[0][DATA][25] , 
        \chs_in_f[0][DATA][24] , \chs_in_f[0][DATA][23] , 
        \chs_in_f[0][DATA][22] , \chs_in_f[0][DATA][21] , 
        \chs_in_f[0][DATA][20] , \chs_in_f[0][DATA][19] , 
        \chs_in_f[0][DATA][18] , \chs_in_f[0][DATA][17] , 
        \chs_in_f[0][DATA][16] , \chs_in_f[0][DATA][15] , 
        \chs_in_f[0][DATA][14] , \chs_in_f[0][DATA][13] , 
        \chs_in_f[0][DATA][12] , \chs_in_f[0][DATA][11] , 
        \chs_in_f[0][DATA][10] , \chs_in_f[0][DATA][9] , 
        \chs_in_f[0][DATA][8] , \chs_in_f[0][DATA][7] , \chs_in_f[0][DATA][6] , 
        \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] , \chs_in_f[0][DATA][3] , 
        \chs_in_f[0][DATA][2] , \chs_in_f[0][DATA][1] , \chs_in_f[0][DATA][0] }), .chan_out_b(\chs_in_b[0][ACK] ), .sel({\switch_sel[0][4] , 
        \switch_sel[0][3] , \switch_sel[0][2] , \switch_sel[0][1] , 
        \switch_sel[0][0] }) );
  hpu_0_2_2 south_hpu ( .preset(n2), .chan_in_f({\south_hpu_f[REQ] , 
        \south_hpu_f[DATA][34] , \south_hpu_f[DATA][33] , 
        \south_hpu_f[DATA][32] , \south_hpu_f[DATA][31] , 
        \south_hpu_f[DATA][30] , \south_hpu_f[DATA][29] , 
        \south_hpu_f[DATA][28] , \south_hpu_f[DATA][27] , 
        \south_hpu_f[DATA][26] , \south_hpu_f[DATA][25] , 
        \south_hpu_f[DATA][24] , \south_hpu_f[DATA][23] , 
        \south_hpu_f[DATA][22] , \south_hpu_f[DATA][21] , 
        \south_hpu_f[DATA][20] , \south_hpu_f[DATA][19] , 
        \south_hpu_f[DATA][18] , \south_hpu_f[DATA][17] , 
        \south_hpu_f[DATA][16] , \south_hpu_f[DATA][15] , 
        \south_hpu_f[DATA][14] , \south_hpu_f[DATA][13] , 
        \south_hpu_f[DATA][12] , \south_hpu_f[DATA][11] , 
        \south_hpu_f[DATA][10] , \south_hpu_f[DATA][9] , 
        \south_hpu_f[DATA][8] , \south_hpu_f[DATA][7] , \south_hpu_f[DATA][6] , 
        \south_hpu_f[DATA][5] , \south_hpu_f[DATA][4] , \south_hpu_f[DATA][3] , 
        \south_hpu_f[DATA][2] , \south_hpu_f[DATA][1] , \south_hpu_f[DATA][0] }), .chan_in_b(\south_hpu_b[ACK] ), .chan_out_f({\chs_in_f[2][REQ] , 
        \chs_in_f[2][DATA][34] , \chs_in_f[2][DATA][33] , 
        \chs_in_f[2][DATA][32] , \chs_in_f[2][DATA][31] , 
        \chs_in_f[2][DATA][30] , \chs_in_f[2][DATA][29] , 
        \chs_in_f[2][DATA][28] , \chs_in_f[2][DATA][27] , 
        \chs_in_f[2][DATA][26] , \chs_in_f[2][DATA][25] , 
        \chs_in_f[2][DATA][24] , \chs_in_f[2][DATA][23] , 
        \chs_in_f[2][DATA][22] , \chs_in_f[2][DATA][21] , 
        \chs_in_f[2][DATA][20] , \chs_in_f[2][DATA][19] , 
        \chs_in_f[2][DATA][18] , \chs_in_f[2][DATA][17] , 
        \chs_in_f[2][DATA][16] , \chs_in_f[2][DATA][15] , 
        \chs_in_f[2][DATA][14] , \chs_in_f[2][DATA][13] , 
        \chs_in_f[2][DATA][12] , \chs_in_f[2][DATA][11] , 
        \chs_in_f[2][DATA][10] , \chs_in_f[2][DATA][9] , 
        \chs_in_f[2][DATA][8] , \chs_in_f[2][DATA][7] , \chs_in_f[2][DATA][6] , 
        \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] , \chs_in_f[2][DATA][3] , 
        \chs_in_f[2][DATA][2] , \chs_in_f[2][DATA][1] , \chs_in_f[2][DATA][0] }), .chan_out_b(\chs_in_b[2][ACK] ), .sel({\switch_sel[2][4] , 
        \switch_sel[2][3] , \switch_sel[2][2] , \switch_sel[2][1] , 
        \switch_sel[2][0] }) );
  hpu_0_1_2 east_hpu ( .preset(n2), .chan_in_f({\east_hpu_f[REQ] , 
        \east_hpu_f[DATA][34] , \east_hpu_f[DATA][33] , \east_hpu_f[DATA][32] , 
        \east_hpu_f[DATA][31] , \east_hpu_f[DATA][30] , \east_hpu_f[DATA][29] , 
        \east_hpu_f[DATA][28] , \east_hpu_f[DATA][27] , \east_hpu_f[DATA][26] , 
        \east_hpu_f[DATA][25] , \east_hpu_f[DATA][24] , \east_hpu_f[DATA][23] , 
        \east_hpu_f[DATA][22] , \east_hpu_f[DATA][21] , \east_hpu_f[DATA][20] , 
        \east_hpu_f[DATA][19] , \east_hpu_f[DATA][18] , \east_hpu_f[DATA][17] , 
        \east_hpu_f[DATA][16] , \east_hpu_f[DATA][15] , \east_hpu_f[DATA][14] , 
        \east_hpu_f[DATA][13] , \east_hpu_f[DATA][12] , \east_hpu_f[DATA][11] , 
        \east_hpu_f[DATA][10] , \east_hpu_f[DATA][9] , \east_hpu_f[DATA][8] , 
        \east_hpu_f[DATA][7] , \east_hpu_f[DATA][6] , \east_hpu_f[DATA][5] , 
        \east_hpu_f[DATA][4] , \east_hpu_f[DATA][3] , \east_hpu_f[DATA][2] , 
        \east_hpu_f[DATA][1] , \east_hpu_f[DATA][0] }), .chan_in_b(
        \east_hpu_b[ACK] ), .chan_out_f({\chs_in_f[1][REQ] , 
        \chs_in_f[1][DATA][34] , \chs_in_f[1][DATA][33] , 
        \chs_in_f[1][DATA][32] , \chs_in_f[1][DATA][31] , 
        \chs_in_f[1][DATA][30] , \chs_in_f[1][DATA][29] , 
        \chs_in_f[1][DATA][28] , \chs_in_f[1][DATA][27] , 
        \chs_in_f[1][DATA][26] , \chs_in_f[1][DATA][25] , 
        \chs_in_f[1][DATA][24] , \chs_in_f[1][DATA][23] , 
        \chs_in_f[1][DATA][22] , \chs_in_f[1][DATA][21] , 
        \chs_in_f[1][DATA][20] , \chs_in_f[1][DATA][19] , 
        \chs_in_f[1][DATA][18] , \chs_in_f[1][DATA][17] , 
        \chs_in_f[1][DATA][16] , \chs_in_f[1][DATA][15] , 
        \chs_in_f[1][DATA][14] , \chs_in_f[1][DATA][13] , 
        \chs_in_f[1][DATA][12] , \chs_in_f[1][DATA][11] , 
        \chs_in_f[1][DATA][10] , \chs_in_f[1][DATA][9] , 
        \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] , \chs_in_f[1][DATA][6] , 
        \chs_in_f[1][DATA][5] , \chs_in_f[1][DATA][4] , \chs_in_f[1][DATA][3] , 
        \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] , \chs_in_f[1][DATA][0] }), .chan_out_b(\chs_in_b[1][ACK] ), .sel({\switch_sel[1][4] , 
        \switch_sel[1][3] , \switch_sel[1][2] , \switch_sel[1][1] , 
        \switch_sel[1][0] }) );
  hpu_0_3_2 west_hpu ( .preset(n2), .chan_in_f({\west_hpu_f[REQ] , 
        \west_hpu_f[DATA][34] , \west_hpu_f[DATA][33] , \west_hpu_f[DATA][32] , 
        \west_hpu_f[DATA][31] , \west_hpu_f[DATA][30] , \west_hpu_f[DATA][29] , 
        \west_hpu_f[DATA][28] , \west_hpu_f[DATA][27] , \west_hpu_f[DATA][26] , 
        \west_hpu_f[DATA][25] , \west_hpu_f[DATA][24] , \west_hpu_f[DATA][23] , 
        \west_hpu_f[DATA][22] , \west_hpu_f[DATA][21] , \west_hpu_f[DATA][20] , 
        \west_hpu_f[DATA][19] , \west_hpu_f[DATA][18] , \west_hpu_f[DATA][17] , 
        \west_hpu_f[DATA][16] , \west_hpu_f[DATA][15] , \west_hpu_f[DATA][14] , 
        \west_hpu_f[DATA][13] , \west_hpu_f[DATA][12] , \west_hpu_f[DATA][11] , 
        \west_hpu_f[DATA][10] , \west_hpu_f[DATA][9] , \west_hpu_f[DATA][8] , 
        \west_hpu_f[DATA][7] , \west_hpu_f[DATA][6] , \west_hpu_f[DATA][5] , 
        \west_hpu_f[DATA][4] , \west_hpu_f[DATA][3] , \west_hpu_f[DATA][2] , 
        \west_hpu_f[DATA][1] , \west_hpu_f[DATA][0] }), .chan_in_b(
        \west_hpu_b[ACK] ), .chan_out_f({\chs_in_f[3][REQ] , 
        \chs_in_f[3][DATA][34] , \chs_in_f[3][DATA][33] , 
        \chs_in_f[3][DATA][32] , \chs_in_f[3][DATA][31] , 
        \chs_in_f[3][DATA][30] , \chs_in_f[3][DATA][29] , 
        \chs_in_f[3][DATA][28] , \chs_in_f[3][DATA][27] , 
        \chs_in_f[3][DATA][26] , \chs_in_f[3][DATA][25] , 
        \chs_in_f[3][DATA][24] , \chs_in_f[3][DATA][23] , 
        \chs_in_f[3][DATA][22] , \chs_in_f[3][DATA][21] , 
        \chs_in_f[3][DATA][20] , \chs_in_f[3][DATA][19] , 
        \chs_in_f[3][DATA][18] , \chs_in_f[3][DATA][17] , 
        \chs_in_f[3][DATA][16] , \chs_in_f[3][DATA][15] , 
        \chs_in_f[3][DATA][14] , \chs_in_f[3][DATA][13] , 
        \chs_in_f[3][DATA][12] , \chs_in_f[3][DATA][11] , 
        \chs_in_f[3][DATA][10] , \chs_in_f[3][DATA][9] , 
        \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] , \chs_in_f[3][DATA][6] , 
        \chs_in_f[3][DATA][5] , \chs_in_f[3][DATA][4] , \chs_in_f[3][DATA][3] , 
        \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] , \chs_in_f[3][DATA][0] }), .chan_out_b(\chs_in_b[3][ACK] ), .sel({\switch_sel[3][4] , 
        \switch_sel[3][3] , \switch_sel[3][2] , \switch_sel[3][1] , 
        \switch_sel[3][0] }) );
  hpu_1_x_2 resource_hpu ( .preset(n2), .chan_in_f({\resource_hpu_f[REQ] , 
        \resource_hpu_f[DATA][34] , \resource_hpu_f[DATA][33] , 
        \resource_hpu_f[DATA][32] , \resource_hpu_f[DATA][31] , 
        \resource_hpu_f[DATA][30] , \resource_hpu_f[DATA][29] , 
        \resource_hpu_f[DATA][28] , \resource_hpu_f[DATA][27] , 
        \resource_hpu_f[DATA][26] , \resource_hpu_f[DATA][25] , 
        \resource_hpu_f[DATA][24] , \resource_hpu_f[DATA][23] , 
        \resource_hpu_f[DATA][22] , \resource_hpu_f[DATA][21] , 
        \resource_hpu_f[DATA][20] , \resource_hpu_f[DATA][19] , 
        \resource_hpu_f[DATA][18] , \resource_hpu_f[DATA][17] , 
        \resource_hpu_f[DATA][16] , \resource_hpu_f[DATA][15] , 
        \resource_hpu_f[DATA][14] , \resource_hpu_f[DATA][13] , 
        \resource_hpu_f[DATA][12] , \resource_hpu_f[DATA][11] , 
        \resource_hpu_f[DATA][10] , \resource_hpu_f[DATA][9] , 
        \resource_hpu_f[DATA][8] , \resource_hpu_f[DATA][7] , 
        \resource_hpu_f[DATA][6] , \resource_hpu_f[DATA][5] , 
        \resource_hpu_f[DATA][4] , \resource_hpu_f[DATA][3] , 
        \resource_hpu_f[DATA][2] , \resource_hpu_f[DATA][1] , 
        \resource_hpu_f[DATA][0] }), .chan_in_b(\resource_hpu_b[ACK] ), 
        .chan_out_f({\chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] , 
        \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] , 
        \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] , 
        \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] , 
        \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] , 
        \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] , 
        \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] , 
        \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] , 
        \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] , 
        \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] , 
        \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] , 
        \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] , 
        \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] , 
        \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] , \chs_in_f[4][DATA][7] , 
        \chs_in_f[4][DATA][6] , \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] , 
        \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] , \chs_in_f[4][DATA][1] , 
        \chs_in_f[4][DATA][0] }), .chan_out_b(\chs_in_b[4][ACK] ), .sel({
        \switch_sel[4][4] , \switch_sel[4][3] , \switch_sel[4][2] , 
        \switch_sel[4][1] , \switch_sel[4][0] }) );
  crossbar_stage_2 xbar_with_latches ( .preset(n3), .switch_sel({1'b0, 
        \switch_sel[4][3] , \switch_sel[4][2] , \switch_sel[4][1] , 
        \switch_sel[4][0] , \switch_sel[3][4] , 1'b0, \switch_sel[3][2] , 
        \switch_sel[3][1] , \switch_sel[3][0] , \switch_sel[2][4] , 
        \switch_sel[2][3] , 1'b0, \switch_sel[2][1] , \switch_sel[2][0] , 
        \switch_sel[1][4] , \switch_sel[1][3] , \switch_sel[1][2] , 1'b0, 
        \switch_sel[1][0] , \switch_sel[0][4] , \switch_sel[0][3] , 
        \switch_sel[0][2] , \switch_sel[0][1] , 1'b0}), .chs_in_f({
        \chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] , \chs_in_f[4][DATA][33] , 
        \chs_in_f[4][DATA][32] , \chs_in_f[4][DATA][31] , 
        \chs_in_f[4][DATA][30] , \chs_in_f[4][DATA][29] , 
        \chs_in_f[4][DATA][28] , \chs_in_f[4][DATA][27] , 
        \chs_in_f[4][DATA][26] , \chs_in_f[4][DATA][25] , 
        \chs_in_f[4][DATA][24] , \chs_in_f[4][DATA][23] , 
        \chs_in_f[4][DATA][22] , \chs_in_f[4][DATA][21] , 
        \chs_in_f[4][DATA][20] , \chs_in_f[4][DATA][19] , 
        \chs_in_f[4][DATA][18] , \chs_in_f[4][DATA][17] , 
        \chs_in_f[4][DATA][16] , \chs_in_f[4][DATA][15] , 
        \chs_in_f[4][DATA][14] , \chs_in_f[4][DATA][13] , 
        \chs_in_f[4][DATA][12] , \chs_in_f[4][DATA][11] , 
        \chs_in_f[4][DATA][10] , \chs_in_f[4][DATA][9] , 
        \chs_in_f[4][DATA][8] , \chs_in_f[4][DATA][7] , \chs_in_f[4][DATA][6] , 
        \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] , \chs_in_f[4][DATA][3] , 
        \chs_in_f[4][DATA][2] , \chs_in_f[4][DATA][1] , \chs_in_f[4][DATA][0] , 
        \chs_in_f[3][REQ] , \chs_in_f[3][DATA][34] , \chs_in_f[3][DATA][33] , 
        \chs_in_f[3][DATA][32] , \chs_in_f[3][DATA][31] , 
        \chs_in_f[3][DATA][30] , \chs_in_f[3][DATA][29] , 
        \chs_in_f[3][DATA][28] , \chs_in_f[3][DATA][27] , 
        \chs_in_f[3][DATA][26] , \chs_in_f[3][DATA][25] , 
        \chs_in_f[3][DATA][24] , \chs_in_f[3][DATA][23] , 
        \chs_in_f[3][DATA][22] , \chs_in_f[3][DATA][21] , 
        \chs_in_f[3][DATA][20] , \chs_in_f[3][DATA][19] , 
        \chs_in_f[3][DATA][18] , \chs_in_f[3][DATA][17] , 
        \chs_in_f[3][DATA][16] , \chs_in_f[3][DATA][15] , 
        \chs_in_f[3][DATA][14] , \chs_in_f[3][DATA][13] , 
        \chs_in_f[3][DATA][12] , \chs_in_f[3][DATA][11] , 
        \chs_in_f[3][DATA][10] , \chs_in_f[3][DATA][9] , 
        \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] , \chs_in_f[3][DATA][6] , 
        \chs_in_f[3][DATA][5] , \chs_in_f[3][DATA][4] , \chs_in_f[3][DATA][3] , 
        \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] , \chs_in_f[3][DATA][0] , 
        \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] , \chs_in_f[2][DATA][33] , 
        \chs_in_f[2][DATA][32] , \chs_in_f[2][DATA][31] , 
        \chs_in_f[2][DATA][30] , \chs_in_f[2][DATA][29] , 
        \chs_in_f[2][DATA][28] , \chs_in_f[2][DATA][27] , 
        \chs_in_f[2][DATA][26] , \chs_in_f[2][DATA][25] , 
        \chs_in_f[2][DATA][24] , \chs_in_f[2][DATA][23] , 
        \chs_in_f[2][DATA][22] , \chs_in_f[2][DATA][21] , 
        \chs_in_f[2][DATA][20] , \chs_in_f[2][DATA][19] , 
        \chs_in_f[2][DATA][18] , \chs_in_f[2][DATA][17] , 
        \chs_in_f[2][DATA][16] , \chs_in_f[2][DATA][15] , 
        \chs_in_f[2][DATA][14] , \chs_in_f[2][DATA][13] , 
        \chs_in_f[2][DATA][12] , \chs_in_f[2][DATA][11] , 
        \chs_in_f[2][DATA][10] , \chs_in_f[2][DATA][9] , 
        \chs_in_f[2][DATA][8] , \chs_in_f[2][DATA][7] , \chs_in_f[2][DATA][6] , 
        \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] , \chs_in_f[2][DATA][3] , 
        \chs_in_f[2][DATA][2] , \chs_in_f[2][DATA][1] , \chs_in_f[2][DATA][0] , 
        \chs_in_f[1][REQ] , \chs_in_f[1][DATA][34] , \chs_in_f[1][DATA][33] , 
        \chs_in_f[1][DATA][32] , \chs_in_f[1][DATA][31] , 
        \chs_in_f[1][DATA][30] , \chs_in_f[1][DATA][29] , 
        \chs_in_f[1][DATA][28] , \chs_in_f[1][DATA][27] , 
        \chs_in_f[1][DATA][26] , \chs_in_f[1][DATA][25] , 
        \chs_in_f[1][DATA][24] , \chs_in_f[1][DATA][23] , 
        \chs_in_f[1][DATA][22] , \chs_in_f[1][DATA][21] , 
        \chs_in_f[1][DATA][20] , \chs_in_f[1][DATA][19] , 
        \chs_in_f[1][DATA][18] , \chs_in_f[1][DATA][17] , 
        \chs_in_f[1][DATA][16] , \chs_in_f[1][DATA][15] , 
        \chs_in_f[1][DATA][14] , \chs_in_f[1][DATA][13] , 
        \chs_in_f[1][DATA][12] , \chs_in_f[1][DATA][11] , 
        \chs_in_f[1][DATA][10] , \chs_in_f[1][DATA][9] , 
        \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] , \chs_in_f[1][DATA][6] , 
        \chs_in_f[1][DATA][5] , \chs_in_f[1][DATA][4] , \chs_in_f[1][DATA][3] , 
        \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] , \chs_in_f[1][DATA][0] , 
        \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] , \chs_in_f[0][DATA][33] , 
        \chs_in_f[0][DATA][32] , \chs_in_f[0][DATA][31] , 
        \chs_in_f[0][DATA][30] , \chs_in_f[0][DATA][29] , 
        \chs_in_f[0][DATA][28] , \chs_in_f[0][DATA][27] , 
        \chs_in_f[0][DATA][26] , \chs_in_f[0][DATA][25] , 
        \chs_in_f[0][DATA][24] , \chs_in_f[0][DATA][23] , 
        \chs_in_f[0][DATA][22] , \chs_in_f[0][DATA][21] , 
        \chs_in_f[0][DATA][20] , \chs_in_f[0][DATA][19] , 
        \chs_in_f[0][DATA][18] , \chs_in_f[0][DATA][17] , 
        \chs_in_f[0][DATA][16] , \chs_in_f[0][DATA][15] , 
        \chs_in_f[0][DATA][14] , \chs_in_f[0][DATA][13] , 
        \chs_in_f[0][DATA][12] , \chs_in_f[0][DATA][11] , 
        \chs_in_f[0][DATA][10] , \chs_in_f[0][DATA][9] , 
        \chs_in_f[0][DATA][8] , \chs_in_f[0][DATA][7] , \chs_in_f[0][DATA][6] , 
        \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] , \chs_in_f[0][DATA][3] , 
        \chs_in_f[0][DATA][2] , \chs_in_f[0][DATA][1] , \chs_in_f[0][DATA][0] }), .chs_in_b({\chs_in_b[4][ACK] , \chs_in_b[3][ACK] , \chs_in_b[2][ACK] , 
        \chs_in_b[1][ACK] , \chs_in_b[0][ACK] }), .latches_out_f({
        \resource_out_f[REQ] , \resource_out_f[DATA][34] , 
        \resource_out_f[DATA][33] , \resource_out_f[DATA][32] , 
        \resource_out_f[DATA][31] , \resource_out_f[DATA][30] , 
        \resource_out_f[DATA][29] , \resource_out_f[DATA][28] , 
        \resource_out_f[DATA][27] , \resource_out_f[DATA][26] , 
        \resource_out_f[DATA][25] , \resource_out_f[DATA][24] , 
        \resource_out_f[DATA][23] , \resource_out_f[DATA][22] , 
        \resource_out_f[DATA][21] , \resource_out_f[DATA][20] , 
        \resource_out_f[DATA][19] , \resource_out_f[DATA][18] , 
        \resource_out_f[DATA][17] , \resource_out_f[DATA][16] , 
        \resource_out_f[DATA][15] , \resource_out_f[DATA][14] , 
        \resource_out_f[DATA][13] , \resource_out_f[DATA][12] , 
        \resource_out_f[DATA][11] , \resource_out_f[DATA][10] , 
        \resource_out_f[DATA][9] , \resource_out_f[DATA][8] , 
        \resource_out_f[DATA][7] , \resource_out_f[DATA][6] , 
        \resource_out_f[DATA][5] , \resource_out_f[DATA][4] , 
        \resource_out_f[DATA][3] , \resource_out_f[DATA][2] , 
        \resource_out_f[DATA][1] , \resource_out_f[DATA][0] , 
        \west_out_f[REQ] , \west_out_f[DATA][34] , \west_out_f[DATA][33] , 
        \west_out_f[DATA][32] , \west_out_f[DATA][31] , \west_out_f[DATA][30] , 
        \west_out_f[DATA][29] , \west_out_f[DATA][28] , \west_out_f[DATA][27] , 
        \west_out_f[DATA][26] , \west_out_f[DATA][25] , \west_out_f[DATA][24] , 
        \west_out_f[DATA][23] , \west_out_f[DATA][22] , \west_out_f[DATA][21] , 
        \west_out_f[DATA][20] , \west_out_f[DATA][19] , \west_out_f[DATA][18] , 
        \west_out_f[DATA][17] , \west_out_f[DATA][16] , \west_out_f[DATA][15] , 
        \west_out_f[DATA][14] , \west_out_f[DATA][13] , \west_out_f[DATA][12] , 
        \west_out_f[DATA][11] , \west_out_f[DATA][10] , \west_out_f[DATA][9] , 
        \west_out_f[DATA][8] , \west_out_f[DATA][7] , \west_out_f[DATA][6] , 
        \west_out_f[DATA][5] , \west_out_f[DATA][4] , \west_out_f[DATA][3] , 
        \west_out_f[DATA][2] , \west_out_f[DATA][1] , \west_out_f[DATA][0] , 
        \south_out_f[REQ] , \south_out_f[DATA][34] , \south_out_f[DATA][33] , 
        \south_out_f[DATA][32] , \south_out_f[DATA][31] , 
        \south_out_f[DATA][30] , \south_out_f[DATA][29] , 
        \south_out_f[DATA][28] , \south_out_f[DATA][27] , 
        \south_out_f[DATA][26] , \south_out_f[DATA][25] , 
        \south_out_f[DATA][24] , \south_out_f[DATA][23] , 
        \south_out_f[DATA][22] , \south_out_f[DATA][21] , 
        \south_out_f[DATA][20] , \south_out_f[DATA][19] , 
        \south_out_f[DATA][18] , \south_out_f[DATA][17] , 
        \south_out_f[DATA][16] , \south_out_f[DATA][15] , 
        \south_out_f[DATA][14] , \south_out_f[DATA][13] , 
        \south_out_f[DATA][12] , \south_out_f[DATA][11] , 
        \south_out_f[DATA][10] , \south_out_f[DATA][9] , 
        \south_out_f[DATA][8] , \south_out_f[DATA][7] , \south_out_f[DATA][6] , 
        \south_out_f[DATA][5] , \south_out_f[DATA][4] , \south_out_f[DATA][3] , 
        \south_out_f[DATA][2] , \south_out_f[DATA][1] , \south_out_f[DATA][0] , 
        \east_out_f[REQ] , \east_out_f[DATA][34] , \east_out_f[DATA][33] , 
        \east_out_f[DATA][32] , \east_out_f[DATA][31] , \east_out_f[DATA][30] , 
        \east_out_f[DATA][29] , \east_out_f[DATA][28] , \east_out_f[DATA][27] , 
        \east_out_f[DATA][26] , \east_out_f[DATA][25] , \east_out_f[DATA][24] , 
        \east_out_f[DATA][23] , \east_out_f[DATA][22] , \east_out_f[DATA][21] , 
        \east_out_f[DATA][20] , \east_out_f[DATA][19] , \east_out_f[DATA][18] , 
        \east_out_f[DATA][17] , \east_out_f[DATA][16] , \east_out_f[DATA][15] , 
        \east_out_f[DATA][14] , \east_out_f[DATA][13] , \east_out_f[DATA][12] , 
        \east_out_f[DATA][11] , \east_out_f[DATA][10] , \east_out_f[DATA][9] , 
        \east_out_f[DATA][8] , \east_out_f[DATA][7] , \east_out_f[DATA][6] , 
        \east_out_f[DATA][5] , \east_out_f[DATA][4] , \east_out_f[DATA][3] , 
        \east_out_f[DATA][2] , \east_out_f[DATA][1] , \east_out_f[DATA][0] , 
        \north_out_f[REQ] , \north_out_f[DATA][34] , \north_out_f[DATA][33] , 
        \north_out_f[DATA][32] , \north_out_f[DATA][31] , 
        \north_out_f[DATA][30] , \north_out_f[DATA][29] , 
        \north_out_f[DATA][28] , \north_out_f[DATA][27] , 
        \north_out_f[DATA][26] , \north_out_f[DATA][25] , 
        \north_out_f[DATA][24] , \north_out_f[DATA][23] , 
        \north_out_f[DATA][22] , \north_out_f[DATA][21] , 
        \north_out_f[DATA][20] , \north_out_f[DATA][19] , 
        \north_out_f[DATA][18] , \north_out_f[DATA][17] , 
        \north_out_f[DATA][16] , \north_out_f[DATA][15] , 
        \north_out_f[DATA][14] , \north_out_f[DATA][13] , 
        \north_out_f[DATA][12] , \north_out_f[DATA][11] , 
        \north_out_f[DATA][10] , \north_out_f[DATA][9] , 
        \north_out_f[DATA][8] , \north_out_f[DATA][7] , \north_out_f[DATA][6] , 
        \north_out_f[DATA][5] , \north_out_f[DATA][4] , \north_out_f[DATA][3] , 
        \north_out_f[DATA][2] , \north_out_f[DATA][1] , \north_out_f[DATA][0] }), .latches_out_b({\resource_out_b[ACK] , \west_out_b[ACK] , 
        \south_out_b[ACK] , \east_out_b[ACK] , \north_out_b[ACK] }) );
  HS65_LS_BFX9 U1 ( .A(preset), .Z(n3) );
  HS65_LS_BFX9 U2 ( .A(preset), .Z(n2) );
endmodule


module noc_node_2 ( p_clk, n_clk, reset, .proc_in({\proc_in[MCMD][1] , 
        \proc_in[MCMD][0] , \proc_in[MADDR][31] , \proc_in[MADDR][30] , 
        \proc_in[MADDR][29] , \proc_in[MADDR][28] , \proc_in[MADDR][27] , 
        \proc_in[MADDR][26] , \proc_in[MADDR][25] , \proc_in[MADDR][24] , 
        \proc_in[MADDR][23] , \proc_in[MADDR][22] , \proc_in[MADDR][21] , 
        \proc_in[MADDR][20] , \proc_in[MADDR][19] , \proc_in[MADDR][18] , 
        \proc_in[MADDR][17] , \proc_in[MADDR][16] , \proc_in[MADDR][15] , 
        \proc_in[MADDR][14] , \proc_in[MADDR][13] , \proc_in[MADDR][12] , 
        \proc_in[MADDR][11] , \proc_in[MADDR][10] , \proc_in[MADDR][9] , 
        \proc_in[MADDR][8] , \proc_in[MADDR][7] , \proc_in[MADDR][6] , 
        \proc_in[MADDR][5] , \proc_in[MADDR][4] , \proc_in[MADDR][3] , 
        \proc_in[MADDR][2] , \proc_in[MADDR][1] , \proc_in[MADDR][0] , 
        \proc_in[MDATA][31] , \proc_in[MDATA][30] , \proc_in[MDATA][29] , 
        \proc_in[MDATA][28] , \proc_in[MDATA][27] , \proc_in[MDATA][26] , 
        \proc_in[MDATA][25] , \proc_in[MDATA][24] , \proc_in[MDATA][23] , 
        \proc_in[MDATA][22] , \proc_in[MDATA][21] , \proc_in[MDATA][20] , 
        \proc_in[MDATA][19] , \proc_in[MDATA][18] , \proc_in[MDATA][17] , 
        \proc_in[MDATA][16] , \proc_in[MDATA][15] , \proc_in[MDATA][14] , 
        \proc_in[MDATA][13] , \proc_in[MDATA][12] , \proc_in[MDATA][11] , 
        \proc_in[MDATA][10] , \proc_in[MDATA][9] , \proc_in[MDATA][8] , 
        \proc_in[MDATA][7] , \proc_in[MDATA][6] , \proc_in[MDATA][5] , 
        \proc_in[MDATA][4] , \proc_in[MDATA][3] , \proc_in[MDATA][2] , 
        \proc_in[MDATA][1] , \proc_in[MDATA][0] }), .proc_out({
        \proc_out[SCMDACCEPT] , \proc_out[SRESP] , \proc_out[SDATA][31] , 
        \proc_out[SDATA][30] , \proc_out[SDATA][29] , \proc_out[SDATA][28] , 
        \proc_out[SDATA][27] , \proc_out[SDATA][26] , \proc_out[SDATA][25] , 
        \proc_out[SDATA][24] , \proc_out[SDATA][23] , \proc_out[SDATA][22] , 
        \proc_out[SDATA][21] , \proc_out[SDATA][20] , \proc_out[SDATA][19] , 
        \proc_out[SDATA][18] , \proc_out[SDATA][17] , \proc_out[SDATA][16] , 
        \proc_out[SDATA][15] , \proc_out[SDATA][14] , \proc_out[SDATA][13] , 
        \proc_out[SDATA][12] , \proc_out[SDATA][11] , \proc_out[SDATA][10] , 
        \proc_out[SDATA][9] , \proc_out[SDATA][8] , \proc_out[SDATA][7] , 
        \proc_out[SDATA][6] , \proc_out[SDATA][5] , \proc_out[SDATA][4] , 
        \proc_out[SDATA][3] , \proc_out[SDATA][2] , \proc_out[SDATA][1] , 
        \proc_out[SDATA][0] }), .spm_in({\spm_in[SCMDACCEPT] , \spm_in[SRESP] , 
        \spm_in[SDATA][63] , \spm_in[SDATA][62] , \spm_in[SDATA][61] , 
        \spm_in[SDATA][60] , \spm_in[SDATA][59] , \spm_in[SDATA][58] , 
        \spm_in[SDATA][57] , \spm_in[SDATA][56] , \spm_in[SDATA][55] , 
        \spm_in[SDATA][54] , \spm_in[SDATA][53] , \spm_in[SDATA][52] , 
        \spm_in[SDATA][51] , \spm_in[SDATA][50] , \spm_in[SDATA][49] , 
        \spm_in[SDATA][48] , \spm_in[SDATA][47] , \spm_in[SDATA][46] , 
        \spm_in[SDATA][45] , \spm_in[SDATA][44] , \spm_in[SDATA][43] , 
        \spm_in[SDATA][42] , \spm_in[SDATA][41] , \spm_in[SDATA][40] , 
        \spm_in[SDATA][39] , \spm_in[SDATA][38] , \spm_in[SDATA][37] , 
        \spm_in[SDATA][36] , \spm_in[SDATA][35] , \spm_in[SDATA][34] , 
        \spm_in[SDATA][33] , \spm_in[SDATA][32] , \spm_in[SDATA][31] , 
        \spm_in[SDATA][30] , \spm_in[SDATA][29] , \spm_in[SDATA][28] , 
        \spm_in[SDATA][27] , \spm_in[SDATA][26] , \spm_in[SDATA][25] , 
        \spm_in[SDATA][24] , \spm_in[SDATA][23] , \spm_in[SDATA][22] , 
        \spm_in[SDATA][21] , \spm_in[SDATA][20] , \spm_in[SDATA][19] , 
        \spm_in[SDATA][18] , \spm_in[SDATA][17] , \spm_in[SDATA][16] , 
        \spm_in[SDATA][15] , \spm_in[SDATA][14] , \spm_in[SDATA][13] , 
        \spm_in[SDATA][12] , \spm_in[SDATA][11] , \spm_in[SDATA][10] , 
        \spm_in[SDATA][9] , \spm_in[SDATA][8] , \spm_in[SDATA][7] , 
        \spm_in[SDATA][6] , \spm_in[SDATA][5] , \spm_in[SDATA][4] , 
        \spm_in[SDATA][3] , \spm_in[SDATA][2] , \spm_in[SDATA][1] , 
        \spm_in[SDATA][0] }), .spm_out({\spm_out[MCMD][1] , \spm_out[MCMD][0] , 
        \spm_out[MADDR][31] , \spm_out[MADDR][30] , \spm_out[MADDR][29] , 
        \spm_out[MADDR][28] , \spm_out[MADDR][27] , \spm_out[MADDR][26] , 
        \spm_out[MADDR][25] , \spm_out[MADDR][24] , \spm_out[MADDR][23] , 
        \spm_out[MADDR][22] , \spm_out[MADDR][21] , \spm_out[MADDR][20] , 
        \spm_out[MADDR][19] , \spm_out[MADDR][18] , \spm_out[MADDR][17] , 
        \spm_out[MADDR][16] , \spm_out[MADDR][15] , \spm_out[MADDR][14] , 
        \spm_out[MADDR][13] , \spm_out[MADDR][12] , \spm_out[MADDR][11] , 
        \spm_out[MADDR][10] , \spm_out[MADDR][9] , \spm_out[MADDR][8] , 
        \spm_out[MADDR][7] , \spm_out[MADDR][6] , \spm_out[MADDR][5] , 
        \spm_out[MADDR][4] , \spm_out[MADDR][3] , \spm_out[MADDR][2] , 
        \spm_out[MADDR][1] , \spm_out[MADDR][0] , \spm_out[MDATA][63] , 
        \spm_out[MDATA][62] , \spm_out[MDATA][61] , \spm_out[MDATA][60] , 
        \spm_out[MDATA][59] , \spm_out[MDATA][58] , \spm_out[MDATA][57] , 
        \spm_out[MDATA][56] , \spm_out[MDATA][55] , \spm_out[MDATA][54] , 
        \spm_out[MDATA][53] , \spm_out[MDATA][52] , \spm_out[MDATA][51] , 
        \spm_out[MDATA][50] , \spm_out[MDATA][49] , \spm_out[MDATA][48] , 
        \spm_out[MDATA][47] , \spm_out[MDATA][46] , \spm_out[MDATA][45] , 
        \spm_out[MDATA][44] , \spm_out[MDATA][43] , \spm_out[MDATA][42] , 
        \spm_out[MDATA][41] , \spm_out[MDATA][40] , \spm_out[MDATA][39] , 
        \spm_out[MDATA][38] , \spm_out[MDATA][37] , \spm_out[MDATA][36] , 
        \spm_out[MDATA][35] , \spm_out[MDATA][34] , \spm_out[MDATA][33] , 
        \spm_out[MDATA][32] , \spm_out[MDATA][31] , \spm_out[MDATA][30] , 
        \spm_out[MDATA][29] , \spm_out[MDATA][28] , \spm_out[MDATA][27] , 
        \spm_out[MDATA][26] , \spm_out[MDATA][25] , \spm_out[MDATA][24] , 
        \spm_out[MDATA][23] , \spm_out[MDATA][22] , \spm_out[MDATA][21] , 
        \spm_out[MDATA][20] , \spm_out[MDATA][19] , \spm_out[MDATA][18] , 
        \spm_out[MDATA][17] , \spm_out[MDATA][16] , \spm_out[MDATA][15] , 
        \spm_out[MDATA][14] , \spm_out[MDATA][13] , \spm_out[MDATA][12] , 
        \spm_out[MDATA][11] , \spm_out[MDATA][10] , \spm_out[MDATA][9] , 
        \spm_out[MDATA][8] , \spm_out[MDATA][7] , \spm_out[MDATA][6] , 
        \spm_out[MDATA][5] , \spm_out[MDATA][4] , \spm_out[MDATA][3] , 
        \spm_out[MDATA][2] , \spm_out[MDATA][1] , \spm_out[MDATA][0] }), 
    .north_in_f({\north_in_f[REQ] , \north_in_f[DATA][34] , 
        \north_in_f[DATA][33] , \north_in_f[DATA][32] , \north_in_f[DATA][31] , 
        \north_in_f[DATA][30] , \north_in_f[DATA][29] , \north_in_f[DATA][28] , 
        \north_in_f[DATA][27] , \north_in_f[DATA][26] , \north_in_f[DATA][25] , 
        \north_in_f[DATA][24] , \north_in_f[DATA][23] , \north_in_f[DATA][22] , 
        \north_in_f[DATA][21] , \north_in_f[DATA][20] , \north_in_f[DATA][19] , 
        \north_in_f[DATA][18] , \north_in_f[DATA][17] , \north_in_f[DATA][16] , 
        \north_in_f[DATA][15] , \north_in_f[DATA][14] , \north_in_f[DATA][13] , 
        \north_in_f[DATA][12] , \north_in_f[DATA][11] , \north_in_f[DATA][10] , 
        \north_in_f[DATA][9] , \north_in_f[DATA][8] , \north_in_f[DATA][7] , 
        \north_in_f[DATA][6] , \north_in_f[DATA][5] , \north_in_f[DATA][4] , 
        \north_in_f[DATA][3] , \north_in_f[DATA][2] , \north_in_f[DATA][1] , 
        \north_in_f[DATA][0] }), .north_in_b(\north_in_b[ACK] ), .east_in_f({
        \east_in_f[REQ] , \east_in_f[DATA][34] , \east_in_f[DATA][33] , 
        \east_in_f[DATA][32] , \east_in_f[DATA][31] , \east_in_f[DATA][30] , 
        \east_in_f[DATA][29] , \east_in_f[DATA][28] , \east_in_f[DATA][27] , 
        \east_in_f[DATA][26] , \east_in_f[DATA][25] , \east_in_f[DATA][24] , 
        \east_in_f[DATA][23] , \east_in_f[DATA][22] , \east_in_f[DATA][21] , 
        \east_in_f[DATA][20] , \east_in_f[DATA][19] , \east_in_f[DATA][18] , 
        \east_in_f[DATA][17] , \east_in_f[DATA][16] , \east_in_f[DATA][15] , 
        \east_in_f[DATA][14] , \east_in_f[DATA][13] , \east_in_f[DATA][12] , 
        \east_in_f[DATA][11] , \east_in_f[DATA][10] , \east_in_f[DATA][9] , 
        \east_in_f[DATA][8] , \east_in_f[DATA][7] , \east_in_f[DATA][6] , 
        \east_in_f[DATA][5] , \east_in_f[DATA][4] , \east_in_f[DATA][3] , 
        \east_in_f[DATA][2] , \east_in_f[DATA][1] , \east_in_f[DATA][0] }), 
    .east_in_b(\east_in_b[ACK] ), .south_in_f({\south_in_f[REQ] , 
        \south_in_f[DATA][34] , \south_in_f[DATA][33] , \south_in_f[DATA][32] , 
        \south_in_f[DATA][31] , \south_in_f[DATA][30] , \south_in_f[DATA][29] , 
        \south_in_f[DATA][28] , \south_in_f[DATA][27] , \south_in_f[DATA][26] , 
        \south_in_f[DATA][25] , \south_in_f[DATA][24] , \south_in_f[DATA][23] , 
        \south_in_f[DATA][22] , \south_in_f[DATA][21] , \south_in_f[DATA][20] , 
        \south_in_f[DATA][19] , \south_in_f[DATA][18] , \south_in_f[DATA][17] , 
        \south_in_f[DATA][16] , \south_in_f[DATA][15] , \south_in_f[DATA][14] , 
        \south_in_f[DATA][13] , \south_in_f[DATA][12] , \south_in_f[DATA][11] , 
        \south_in_f[DATA][10] , \south_in_f[DATA][9] , \south_in_f[DATA][8] , 
        \south_in_f[DATA][7] , \south_in_f[DATA][6] , \south_in_f[DATA][5] , 
        \south_in_f[DATA][4] , \south_in_f[DATA][3] , \south_in_f[DATA][2] , 
        \south_in_f[DATA][1] , \south_in_f[DATA][0] }), .south_in_b(
        \south_in_b[ACK] ), .west_in_f({\west_in_f[REQ] , 
        \west_in_f[DATA][34] , \west_in_f[DATA][33] , \west_in_f[DATA][32] , 
        \west_in_f[DATA][31] , \west_in_f[DATA][30] , \west_in_f[DATA][29] , 
        \west_in_f[DATA][28] , \west_in_f[DATA][27] , \west_in_f[DATA][26] , 
        \west_in_f[DATA][25] , \west_in_f[DATA][24] , \west_in_f[DATA][23] , 
        \west_in_f[DATA][22] , \west_in_f[DATA][21] , \west_in_f[DATA][20] , 
        \west_in_f[DATA][19] , \west_in_f[DATA][18] , \west_in_f[DATA][17] , 
        \west_in_f[DATA][16] , \west_in_f[DATA][15] , \west_in_f[DATA][14] , 
        \west_in_f[DATA][13] , \west_in_f[DATA][12] , \west_in_f[DATA][11] , 
        \west_in_f[DATA][10] , \west_in_f[DATA][9] , \west_in_f[DATA][8] , 
        \west_in_f[DATA][7] , \west_in_f[DATA][6] , \west_in_f[DATA][5] , 
        \west_in_f[DATA][4] , \west_in_f[DATA][3] , \west_in_f[DATA][2] , 
        \west_in_f[DATA][1] , \west_in_f[DATA][0] }), .west_in_b(
        \west_in_b[ACK] ), .north_out_f({\north_out_f[REQ] , 
        \north_out_f[DATA][34] , \north_out_f[DATA][33] , 
        \north_out_f[DATA][32] , \north_out_f[DATA][31] , 
        \north_out_f[DATA][30] , \north_out_f[DATA][29] , 
        \north_out_f[DATA][28] , \north_out_f[DATA][27] , 
        \north_out_f[DATA][26] , \north_out_f[DATA][25] , 
        \north_out_f[DATA][24] , \north_out_f[DATA][23] , 
        \north_out_f[DATA][22] , \north_out_f[DATA][21] , 
        \north_out_f[DATA][20] , \north_out_f[DATA][19] , 
        \north_out_f[DATA][18] , \north_out_f[DATA][17] , 
        \north_out_f[DATA][16] , \north_out_f[DATA][15] , 
        \north_out_f[DATA][14] , \north_out_f[DATA][13] , 
        \north_out_f[DATA][12] , \north_out_f[DATA][11] , 
        \north_out_f[DATA][10] , \north_out_f[DATA][9] , 
        \north_out_f[DATA][8] , \north_out_f[DATA][7] , \north_out_f[DATA][6] , 
        \north_out_f[DATA][5] , \north_out_f[DATA][4] , \north_out_f[DATA][3] , 
        \north_out_f[DATA][2] , \north_out_f[DATA][1] , \north_out_f[DATA][0] 
        }), .north_out_b(\north_out_b[ACK] ), .east_out_f({\east_out_f[REQ] , 
        \east_out_f[DATA][34] , \east_out_f[DATA][33] , \east_out_f[DATA][32] , 
        \east_out_f[DATA][31] , \east_out_f[DATA][30] , \east_out_f[DATA][29] , 
        \east_out_f[DATA][28] , \east_out_f[DATA][27] , \east_out_f[DATA][26] , 
        \east_out_f[DATA][25] , \east_out_f[DATA][24] , \east_out_f[DATA][23] , 
        \east_out_f[DATA][22] , \east_out_f[DATA][21] , \east_out_f[DATA][20] , 
        \east_out_f[DATA][19] , \east_out_f[DATA][18] , \east_out_f[DATA][17] , 
        \east_out_f[DATA][16] , \east_out_f[DATA][15] , \east_out_f[DATA][14] , 
        \east_out_f[DATA][13] , \east_out_f[DATA][12] , \east_out_f[DATA][11] , 
        \east_out_f[DATA][10] , \east_out_f[DATA][9] , \east_out_f[DATA][8] , 
        \east_out_f[DATA][7] , \east_out_f[DATA][6] , \east_out_f[DATA][5] , 
        \east_out_f[DATA][4] , \east_out_f[DATA][3] , \east_out_f[DATA][2] , 
        \east_out_f[DATA][1] , \east_out_f[DATA][0] }), .east_out_b(
        \east_out_b[ACK] ), .south_out_f({\south_out_f[REQ] , 
        \south_out_f[DATA][34] , \south_out_f[DATA][33] , 
        \south_out_f[DATA][32] , \south_out_f[DATA][31] , 
        \south_out_f[DATA][30] , \south_out_f[DATA][29] , 
        \south_out_f[DATA][28] , \south_out_f[DATA][27] , 
        \south_out_f[DATA][26] , \south_out_f[DATA][25] , 
        \south_out_f[DATA][24] , \south_out_f[DATA][23] , 
        \south_out_f[DATA][22] , \south_out_f[DATA][21] , 
        \south_out_f[DATA][20] , \south_out_f[DATA][19] , 
        \south_out_f[DATA][18] , \south_out_f[DATA][17] , 
        \south_out_f[DATA][16] , \south_out_f[DATA][15] , 
        \south_out_f[DATA][14] , \south_out_f[DATA][13] , 
        \south_out_f[DATA][12] , \south_out_f[DATA][11] , 
        \south_out_f[DATA][10] , \south_out_f[DATA][9] , 
        \south_out_f[DATA][8] , \south_out_f[DATA][7] , \south_out_f[DATA][6] , 
        \south_out_f[DATA][5] , \south_out_f[DATA][4] , \south_out_f[DATA][3] , 
        \south_out_f[DATA][2] , \south_out_f[DATA][1] , \south_out_f[DATA][0] 
        }), .south_out_b(\south_out_b[ACK] ), .west_out_f({\west_out_f[REQ] , 
        \west_out_f[DATA][34] , \west_out_f[DATA][33] , \west_out_f[DATA][32] , 
        \west_out_f[DATA][31] , \west_out_f[DATA][30] , \west_out_f[DATA][29] , 
        \west_out_f[DATA][28] , \west_out_f[DATA][27] , \west_out_f[DATA][26] , 
        \west_out_f[DATA][25] , \west_out_f[DATA][24] , \west_out_f[DATA][23] , 
        \west_out_f[DATA][22] , \west_out_f[DATA][21] , \west_out_f[DATA][20] , 
        \west_out_f[DATA][19] , \west_out_f[DATA][18] , \west_out_f[DATA][17] , 
        \west_out_f[DATA][16] , \west_out_f[DATA][15] , \west_out_f[DATA][14] , 
        \west_out_f[DATA][13] , \west_out_f[DATA][12] , \west_out_f[DATA][11] , 
        \west_out_f[DATA][10] , \west_out_f[DATA][9] , \west_out_f[DATA][8] , 
        \west_out_f[DATA][7] , \west_out_f[DATA][6] , \west_out_f[DATA][5] , 
        \west_out_f[DATA][4] , \west_out_f[DATA][3] , \west_out_f[DATA][2] , 
        \west_out_f[DATA][1] , \west_out_f[DATA][0] }), .west_out_b(
        \west_out_b[ACK] ) );
  input p_clk, n_clk, reset, \proc_in[MCMD][1] , \proc_in[MCMD][0] ,
         \proc_in[MADDR][31] , \proc_in[MADDR][30] , \proc_in[MADDR][29] ,
         \proc_in[MADDR][28] , \proc_in[MADDR][27] , \proc_in[MADDR][26] ,
         \proc_in[MADDR][25] , \proc_in[MADDR][24] , \proc_in[MADDR][23] ,
         \proc_in[MADDR][22] , \proc_in[MADDR][21] , \proc_in[MADDR][20] ,
         \proc_in[MADDR][19] , \proc_in[MADDR][18] , \proc_in[MADDR][17] ,
         \proc_in[MADDR][16] , \proc_in[MADDR][15] , \proc_in[MADDR][14] ,
         \proc_in[MADDR][13] , \proc_in[MADDR][12] , \proc_in[MADDR][11] ,
         \proc_in[MADDR][10] , \proc_in[MADDR][9] , \proc_in[MADDR][8] ,
         \proc_in[MADDR][7] , \proc_in[MADDR][6] , \proc_in[MADDR][5] ,
         \proc_in[MADDR][4] , \proc_in[MADDR][3] , \proc_in[MADDR][2] ,
         \proc_in[MADDR][1] , \proc_in[MADDR][0] , \proc_in[MDATA][31] ,
         \proc_in[MDATA][30] , \proc_in[MDATA][29] , \proc_in[MDATA][28] ,
         \proc_in[MDATA][27] , \proc_in[MDATA][26] , \proc_in[MDATA][25] ,
         \proc_in[MDATA][24] , \proc_in[MDATA][23] , \proc_in[MDATA][22] ,
         \proc_in[MDATA][21] , \proc_in[MDATA][20] , \proc_in[MDATA][19] ,
         \proc_in[MDATA][18] , \proc_in[MDATA][17] , \proc_in[MDATA][16] ,
         \proc_in[MDATA][15] , \proc_in[MDATA][14] , \proc_in[MDATA][13] ,
         \proc_in[MDATA][12] , \proc_in[MDATA][11] , \proc_in[MDATA][10] ,
         \proc_in[MDATA][9] , \proc_in[MDATA][8] , \proc_in[MDATA][7] ,
         \proc_in[MDATA][6] , \proc_in[MDATA][5] , \proc_in[MDATA][4] ,
         \proc_in[MDATA][3] , \proc_in[MDATA][2] , \proc_in[MDATA][1] ,
         \proc_in[MDATA][0] , \spm_in[SCMDACCEPT] , \spm_in[SRESP] ,
         \spm_in[SDATA][63] , \spm_in[SDATA][62] , \spm_in[SDATA][61] ,
         \spm_in[SDATA][60] , \spm_in[SDATA][59] , \spm_in[SDATA][58] ,
         \spm_in[SDATA][57] , \spm_in[SDATA][56] , \spm_in[SDATA][55] ,
         \spm_in[SDATA][54] , \spm_in[SDATA][53] , \spm_in[SDATA][52] ,
         \spm_in[SDATA][51] , \spm_in[SDATA][50] , \spm_in[SDATA][49] ,
         \spm_in[SDATA][48] , \spm_in[SDATA][47] , \spm_in[SDATA][46] ,
         \spm_in[SDATA][45] , \spm_in[SDATA][44] , \spm_in[SDATA][43] ,
         \spm_in[SDATA][42] , \spm_in[SDATA][41] , \spm_in[SDATA][40] ,
         \spm_in[SDATA][39] , \spm_in[SDATA][38] , \spm_in[SDATA][37] ,
         \spm_in[SDATA][36] , \spm_in[SDATA][35] , \spm_in[SDATA][34] ,
         \spm_in[SDATA][33] , \spm_in[SDATA][32] , \spm_in[SDATA][31] ,
         \spm_in[SDATA][30] , \spm_in[SDATA][29] , \spm_in[SDATA][28] ,
         \spm_in[SDATA][27] , \spm_in[SDATA][26] , \spm_in[SDATA][25] ,
         \spm_in[SDATA][24] , \spm_in[SDATA][23] , \spm_in[SDATA][22] ,
         \spm_in[SDATA][21] , \spm_in[SDATA][20] , \spm_in[SDATA][19] ,
         \spm_in[SDATA][18] , \spm_in[SDATA][17] , \spm_in[SDATA][16] ,
         \spm_in[SDATA][15] , \spm_in[SDATA][14] , \spm_in[SDATA][13] ,
         \spm_in[SDATA][12] , \spm_in[SDATA][11] , \spm_in[SDATA][10] ,
         \spm_in[SDATA][9] , \spm_in[SDATA][8] , \spm_in[SDATA][7] ,
         \spm_in[SDATA][6] , \spm_in[SDATA][5] , \spm_in[SDATA][4] ,
         \spm_in[SDATA][3] , \spm_in[SDATA][2] , \spm_in[SDATA][1] ,
         \spm_in[SDATA][0] , \north_in_f[REQ] , \north_in_f[DATA][34] ,
         \north_in_f[DATA][33] , \north_in_f[DATA][32] ,
         \north_in_f[DATA][31] , \north_in_f[DATA][30] ,
         \north_in_f[DATA][29] , \north_in_f[DATA][28] ,
         \north_in_f[DATA][27] , \north_in_f[DATA][26] ,
         \north_in_f[DATA][25] , \north_in_f[DATA][24] ,
         \north_in_f[DATA][23] , \north_in_f[DATA][22] ,
         \north_in_f[DATA][21] , \north_in_f[DATA][20] ,
         \north_in_f[DATA][19] , \north_in_f[DATA][18] ,
         \north_in_f[DATA][17] , \north_in_f[DATA][16] ,
         \north_in_f[DATA][15] , \north_in_f[DATA][14] ,
         \north_in_f[DATA][13] , \north_in_f[DATA][12] ,
         \north_in_f[DATA][11] , \north_in_f[DATA][10] , \north_in_f[DATA][9] ,
         \north_in_f[DATA][8] , \north_in_f[DATA][7] , \north_in_f[DATA][6] ,
         \north_in_f[DATA][5] , \north_in_f[DATA][4] , \north_in_f[DATA][3] ,
         \north_in_f[DATA][2] , \north_in_f[DATA][1] , \north_in_f[DATA][0] ,
         \east_in_f[REQ] , \east_in_f[DATA][34] , \east_in_f[DATA][33] ,
         \east_in_f[DATA][32] , \east_in_f[DATA][31] , \east_in_f[DATA][30] ,
         \east_in_f[DATA][29] , \east_in_f[DATA][28] , \east_in_f[DATA][27] ,
         \east_in_f[DATA][26] , \east_in_f[DATA][25] , \east_in_f[DATA][24] ,
         \east_in_f[DATA][23] , \east_in_f[DATA][22] , \east_in_f[DATA][21] ,
         \east_in_f[DATA][20] , \east_in_f[DATA][19] , \east_in_f[DATA][18] ,
         \east_in_f[DATA][17] , \east_in_f[DATA][16] , \east_in_f[DATA][15] ,
         \east_in_f[DATA][14] , \east_in_f[DATA][13] , \east_in_f[DATA][12] ,
         \east_in_f[DATA][11] , \east_in_f[DATA][10] , \east_in_f[DATA][9] ,
         \east_in_f[DATA][8] , \east_in_f[DATA][7] , \east_in_f[DATA][6] ,
         \east_in_f[DATA][5] , \east_in_f[DATA][4] , \east_in_f[DATA][3] ,
         \east_in_f[DATA][2] , \east_in_f[DATA][1] , \east_in_f[DATA][0] ,
         \south_in_f[REQ] , \south_in_f[DATA][34] , \south_in_f[DATA][33] ,
         \south_in_f[DATA][32] , \south_in_f[DATA][31] ,
         \south_in_f[DATA][30] , \south_in_f[DATA][29] ,
         \south_in_f[DATA][28] , \south_in_f[DATA][27] ,
         \south_in_f[DATA][26] , \south_in_f[DATA][25] ,
         \south_in_f[DATA][24] , \south_in_f[DATA][23] ,
         \south_in_f[DATA][22] , \south_in_f[DATA][21] ,
         \south_in_f[DATA][20] , \south_in_f[DATA][19] ,
         \south_in_f[DATA][18] , \south_in_f[DATA][17] ,
         \south_in_f[DATA][16] , \south_in_f[DATA][15] ,
         \south_in_f[DATA][14] , \south_in_f[DATA][13] ,
         \south_in_f[DATA][12] , \south_in_f[DATA][11] ,
         \south_in_f[DATA][10] , \south_in_f[DATA][9] , \south_in_f[DATA][8] ,
         \south_in_f[DATA][7] , \south_in_f[DATA][6] , \south_in_f[DATA][5] ,
         \south_in_f[DATA][4] , \south_in_f[DATA][3] , \south_in_f[DATA][2] ,
         \south_in_f[DATA][1] , \south_in_f[DATA][0] , \west_in_f[REQ] ,
         \west_in_f[DATA][34] , \west_in_f[DATA][33] , \west_in_f[DATA][32] ,
         \west_in_f[DATA][31] , \west_in_f[DATA][30] , \west_in_f[DATA][29] ,
         \west_in_f[DATA][28] , \west_in_f[DATA][27] , \west_in_f[DATA][26] ,
         \west_in_f[DATA][25] , \west_in_f[DATA][24] , \west_in_f[DATA][23] ,
         \west_in_f[DATA][22] , \west_in_f[DATA][21] , \west_in_f[DATA][20] ,
         \west_in_f[DATA][19] , \west_in_f[DATA][18] , \west_in_f[DATA][17] ,
         \west_in_f[DATA][16] , \west_in_f[DATA][15] , \west_in_f[DATA][14] ,
         \west_in_f[DATA][13] , \west_in_f[DATA][12] , \west_in_f[DATA][11] ,
         \west_in_f[DATA][10] , \west_in_f[DATA][9] , \west_in_f[DATA][8] ,
         \west_in_f[DATA][7] , \west_in_f[DATA][6] , \west_in_f[DATA][5] ,
         \west_in_f[DATA][4] , \west_in_f[DATA][3] , \west_in_f[DATA][2] ,
         \west_in_f[DATA][1] , \west_in_f[DATA][0] , \north_out_b[ACK] ,
         \east_out_b[ACK] , \south_out_b[ACK] , \west_out_b[ACK] ;
  output \proc_out[SCMDACCEPT] , \proc_out[SRESP] , \proc_out[SDATA][31] ,
         \proc_out[SDATA][30] , \proc_out[SDATA][29] , \proc_out[SDATA][28] ,
         \proc_out[SDATA][27] , \proc_out[SDATA][26] , \proc_out[SDATA][25] ,
         \proc_out[SDATA][24] , \proc_out[SDATA][23] , \proc_out[SDATA][22] ,
         \proc_out[SDATA][21] , \proc_out[SDATA][20] , \proc_out[SDATA][19] ,
         \proc_out[SDATA][18] , \proc_out[SDATA][17] , \proc_out[SDATA][16] ,
         \proc_out[SDATA][15] , \proc_out[SDATA][14] , \proc_out[SDATA][13] ,
         \proc_out[SDATA][12] , \proc_out[SDATA][11] , \proc_out[SDATA][10] ,
         \proc_out[SDATA][9] , \proc_out[SDATA][8] , \proc_out[SDATA][7] ,
         \proc_out[SDATA][6] , \proc_out[SDATA][5] , \proc_out[SDATA][4] ,
         \proc_out[SDATA][3] , \proc_out[SDATA][2] , \proc_out[SDATA][1] ,
         \proc_out[SDATA][0] , \spm_out[MCMD][1] , \spm_out[MCMD][0] ,
         \spm_out[MADDR][31] , \spm_out[MADDR][30] , \spm_out[MADDR][29] ,
         \spm_out[MADDR][28] , \spm_out[MADDR][27] , \spm_out[MADDR][26] ,
         \spm_out[MADDR][25] , \spm_out[MADDR][24] , \spm_out[MADDR][23] ,
         \spm_out[MADDR][22] , \spm_out[MADDR][21] , \spm_out[MADDR][20] ,
         \spm_out[MADDR][19] , \spm_out[MADDR][18] , \spm_out[MADDR][17] ,
         \spm_out[MADDR][16] , \spm_out[MADDR][15] , \spm_out[MADDR][14] ,
         \spm_out[MADDR][13] , \spm_out[MADDR][12] , \spm_out[MADDR][11] ,
         \spm_out[MADDR][10] , \spm_out[MADDR][9] , \spm_out[MADDR][8] ,
         \spm_out[MADDR][7] , \spm_out[MADDR][6] , \spm_out[MADDR][5] ,
         \spm_out[MADDR][4] , \spm_out[MADDR][3] , \spm_out[MADDR][2] ,
         \spm_out[MADDR][1] , \spm_out[MADDR][0] , \spm_out[MDATA][63] ,
         \spm_out[MDATA][62] , \spm_out[MDATA][61] , \spm_out[MDATA][60] ,
         \spm_out[MDATA][59] , \spm_out[MDATA][58] , \spm_out[MDATA][57] ,
         \spm_out[MDATA][56] , \spm_out[MDATA][55] , \spm_out[MDATA][54] ,
         \spm_out[MDATA][53] , \spm_out[MDATA][52] , \spm_out[MDATA][51] ,
         \spm_out[MDATA][50] , \spm_out[MDATA][49] , \spm_out[MDATA][48] ,
         \spm_out[MDATA][47] , \spm_out[MDATA][46] , \spm_out[MDATA][45] ,
         \spm_out[MDATA][44] , \spm_out[MDATA][43] , \spm_out[MDATA][42] ,
         \spm_out[MDATA][41] , \spm_out[MDATA][40] , \spm_out[MDATA][39] ,
         \spm_out[MDATA][38] , \spm_out[MDATA][37] , \spm_out[MDATA][36] ,
         \spm_out[MDATA][35] , \spm_out[MDATA][34] , \spm_out[MDATA][33] ,
         \spm_out[MDATA][32] , \spm_out[MDATA][31] , \spm_out[MDATA][30] ,
         \spm_out[MDATA][29] , \spm_out[MDATA][28] , \spm_out[MDATA][27] ,
         \spm_out[MDATA][26] , \spm_out[MDATA][25] , \spm_out[MDATA][24] ,
         \spm_out[MDATA][23] , \spm_out[MDATA][22] , \spm_out[MDATA][21] ,
         \spm_out[MDATA][20] , \spm_out[MDATA][19] , \spm_out[MDATA][18] ,
         \spm_out[MDATA][17] , \spm_out[MDATA][16] , \spm_out[MDATA][15] ,
         \spm_out[MDATA][14] , \spm_out[MDATA][13] , \spm_out[MDATA][12] ,
         \spm_out[MDATA][11] , \spm_out[MDATA][10] , \spm_out[MDATA][9] ,
         \spm_out[MDATA][8] , \spm_out[MDATA][7] , \spm_out[MDATA][6] ,
         \spm_out[MDATA][5] , \spm_out[MDATA][4] , \spm_out[MDATA][3] ,
         \spm_out[MDATA][2] , \spm_out[MDATA][1] , \spm_out[MDATA][0] ,
         \north_in_b[ACK] , \east_in_b[ACK] , \south_in_b[ACK] ,
         \west_in_b[ACK] , \north_out_f[REQ] , \north_out_f[DATA][34] ,
         \north_out_f[DATA][33] , \north_out_f[DATA][32] ,
         \north_out_f[DATA][31] , \north_out_f[DATA][30] ,
         \north_out_f[DATA][29] , \north_out_f[DATA][28] ,
         \north_out_f[DATA][27] , \north_out_f[DATA][26] ,
         \north_out_f[DATA][25] , \north_out_f[DATA][24] ,
         \north_out_f[DATA][23] , \north_out_f[DATA][22] ,
         \north_out_f[DATA][21] , \north_out_f[DATA][20] ,
         \north_out_f[DATA][19] , \north_out_f[DATA][18] ,
         \north_out_f[DATA][17] , \north_out_f[DATA][16] ,
         \north_out_f[DATA][15] , \north_out_f[DATA][14] ,
         \north_out_f[DATA][13] , \north_out_f[DATA][12] ,
         \north_out_f[DATA][11] , \north_out_f[DATA][10] ,
         \north_out_f[DATA][9] , \north_out_f[DATA][8] ,
         \north_out_f[DATA][7] , \north_out_f[DATA][6] ,
         \north_out_f[DATA][5] , \north_out_f[DATA][4] ,
         \north_out_f[DATA][3] , \north_out_f[DATA][2] ,
         \north_out_f[DATA][1] , \north_out_f[DATA][0] , \east_out_f[REQ] ,
         \east_out_f[DATA][34] , \east_out_f[DATA][33] ,
         \east_out_f[DATA][32] , \east_out_f[DATA][31] ,
         \east_out_f[DATA][30] , \east_out_f[DATA][29] ,
         \east_out_f[DATA][28] , \east_out_f[DATA][27] ,
         \east_out_f[DATA][26] , \east_out_f[DATA][25] ,
         \east_out_f[DATA][24] , \east_out_f[DATA][23] ,
         \east_out_f[DATA][22] , \east_out_f[DATA][21] ,
         \east_out_f[DATA][20] , \east_out_f[DATA][19] ,
         \east_out_f[DATA][18] , \east_out_f[DATA][17] ,
         \east_out_f[DATA][16] , \east_out_f[DATA][15] ,
         \east_out_f[DATA][14] , \east_out_f[DATA][13] ,
         \east_out_f[DATA][12] , \east_out_f[DATA][11] ,
         \east_out_f[DATA][10] , \east_out_f[DATA][9] , \east_out_f[DATA][8] ,
         \east_out_f[DATA][7] , \east_out_f[DATA][6] , \east_out_f[DATA][5] ,
         \east_out_f[DATA][4] , \east_out_f[DATA][3] , \east_out_f[DATA][2] ,
         \east_out_f[DATA][1] , \east_out_f[DATA][0] , \south_out_f[REQ] ,
         \south_out_f[DATA][34] , \south_out_f[DATA][33] ,
         \south_out_f[DATA][32] , \south_out_f[DATA][31] ,
         \south_out_f[DATA][30] , \south_out_f[DATA][29] ,
         \south_out_f[DATA][28] , \south_out_f[DATA][27] ,
         \south_out_f[DATA][26] , \south_out_f[DATA][25] ,
         \south_out_f[DATA][24] , \south_out_f[DATA][23] ,
         \south_out_f[DATA][22] , \south_out_f[DATA][21] ,
         \south_out_f[DATA][20] , \south_out_f[DATA][19] ,
         \south_out_f[DATA][18] , \south_out_f[DATA][17] ,
         \south_out_f[DATA][16] , \south_out_f[DATA][15] ,
         \south_out_f[DATA][14] , \south_out_f[DATA][13] ,
         \south_out_f[DATA][12] , \south_out_f[DATA][11] ,
         \south_out_f[DATA][10] , \south_out_f[DATA][9] ,
         \south_out_f[DATA][8] , \south_out_f[DATA][7] ,
         \south_out_f[DATA][6] , \south_out_f[DATA][5] ,
         \south_out_f[DATA][4] , \south_out_f[DATA][3] ,
         \south_out_f[DATA][2] , \south_out_f[DATA][1] ,
         \south_out_f[DATA][0] , \west_out_f[REQ] , \west_out_f[DATA][34] ,
         \west_out_f[DATA][33] , \west_out_f[DATA][32] ,
         \west_out_f[DATA][31] , \west_out_f[DATA][30] ,
         \west_out_f[DATA][29] , \west_out_f[DATA][28] ,
         \west_out_f[DATA][27] , \west_out_f[DATA][26] ,
         \west_out_f[DATA][25] , \west_out_f[DATA][24] ,
         \west_out_f[DATA][23] , \west_out_f[DATA][22] ,
         \west_out_f[DATA][21] , \west_out_f[DATA][20] ,
         \west_out_f[DATA][19] , \west_out_f[DATA][18] ,
         \west_out_f[DATA][17] , \west_out_f[DATA][16] ,
         \west_out_f[DATA][15] , \west_out_f[DATA][14] ,
         \west_out_f[DATA][13] , \west_out_f[DATA][12] ,
         \west_out_f[DATA][11] , \west_out_f[DATA][10] , \west_out_f[DATA][9] ,
         \west_out_f[DATA][8] , \west_out_f[DATA][7] , \west_out_f[DATA][6] ,
         \west_out_f[DATA][5] , \west_out_f[DATA][4] , \west_out_f[DATA][3] ,
         \west_out_f[DATA][2] , \west_out_f[DATA][1] , \west_out_f[DATA][0] ;
  wire   del_half_clk0, \ip_to_net_f[REQ] , n1, n3, n4, n5, n6, n7, n8, n9,
         n10, n11;
  wire   [34:0] net_to_ip;
  wire   [34:0] ip_to_net;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17;
  assign \spm_out[MADDR][31]  = 1'b0;
  assign \spm_out[MADDR][30]  = 1'b0;
  assign \spm_out[MADDR][29]  = 1'b0;
  assign \spm_out[MADDR][28]  = 1'b0;
  assign \spm_out[MADDR][27]  = 1'b0;
  assign \spm_out[MADDR][26]  = 1'b0;
  assign \spm_out[MADDR][25]  = 1'b0;
  assign \spm_out[MADDR][24]  = 1'b0;
  assign \spm_out[MADDR][23]  = 1'b0;
  assign \spm_out[MADDR][22]  = 1'b0;
  assign \spm_out[MADDR][21]  = 1'b0;
  assign \spm_out[MADDR][20]  = 1'b0;
  assign \spm_out[MADDR][19]  = 1'b0;
  assign \spm_out[MADDR][18]  = 1'b0;
  assign \spm_out[MADDR][17]  = 1'b0;
  assign \spm_out[MADDR][16]  = 1'b0;
  assign \spm_out[MADDR][15]  = 1'b0;

  nAdapter_2 na ( .na_clk(n_clk), .na_reset(reset), .proc_in({
        \proc_in[MCMD][1] , \proc_in[MCMD][0] , \proc_in[MADDR][31] , 
        \proc_in[MADDR][30] , \proc_in[MADDR][29] , \proc_in[MADDR][28] , 
        \proc_in[MADDR][27] , \proc_in[MADDR][26] , \proc_in[MADDR][25] , 
        \proc_in[MADDR][24] , \proc_in[MADDR][23] , \proc_in[MADDR][22] , 
        \proc_in[MADDR][21] , \proc_in[MADDR][20] , \proc_in[MADDR][19] , 
        \proc_in[MADDR][18] , \proc_in[MADDR][17] , \proc_in[MADDR][16] , 
        \proc_in[MADDR][15] , \proc_in[MADDR][14] , \proc_in[MADDR][13] , 
        \proc_in[MADDR][12] , \proc_in[MADDR][11] , \proc_in[MADDR][10] , 
        \proc_in[MADDR][9] , \proc_in[MADDR][8] , \proc_in[MADDR][7] , 
        \proc_in[MADDR][6] , \proc_in[MADDR][5] , \proc_in[MADDR][4] , 
        \proc_in[MADDR][3] , \proc_in[MADDR][2] , \proc_in[MADDR][1] , 
        \proc_in[MADDR][0] , \proc_in[MDATA][31] , \proc_in[MDATA][30] , 
        \proc_in[MDATA][29] , \proc_in[MDATA][28] , \proc_in[MDATA][27] , 
        \proc_in[MDATA][26] , \proc_in[MDATA][25] , \proc_in[MDATA][24] , 
        \proc_in[MDATA][23] , \proc_in[MDATA][22] , \proc_in[MDATA][21] , 
        \proc_in[MDATA][20] , \proc_in[MDATA][19] , \proc_in[MDATA][18] , 
        \proc_in[MDATA][17] , \proc_in[MDATA][16] , \proc_in[MDATA][15] , 
        \proc_in[MDATA][14] , \proc_in[MDATA][13] , \proc_in[MDATA][12] , 
        \proc_in[MDATA][11] , \proc_in[MDATA][10] , \proc_in[MDATA][9] , 
        \proc_in[MDATA][8] , \proc_in[MDATA][7] , \proc_in[MDATA][6] , 
        \proc_in[MDATA][5] , \proc_in[MDATA][4] , \proc_in[MDATA][3] , 
        \proc_in[MDATA][2] , \proc_in[MDATA][1] , \proc_in[MDATA][0] }), 
        .proc_out({\proc_out[SCMDACCEPT] , \proc_out[SRESP] , 
        \proc_out[SDATA][31] , \proc_out[SDATA][30] , \proc_out[SDATA][29] , 
        \proc_out[SDATA][28] , \proc_out[SDATA][27] , \proc_out[SDATA][26] , 
        \proc_out[SDATA][25] , \proc_out[SDATA][24] , \proc_out[SDATA][23] , 
        \proc_out[SDATA][22] , \proc_out[SDATA][21] , \proc_out[SDATA][20] , 
        \proc_out[SDATA][19] , \proc_out[SDATA][18] , \proc_out[SDATA][17] , 
        \proc_out[SDATA][16] , \proc_out[SDATA][15] , \proc_out[SDATA][14] , 
        \proc_out[SDATA][13] , \proc_out[SDATA][12] , \proc_out[SDATA][11] , 
        \proc_out[SDATA][10] , \proc_out[SDATA][9] , \proc_out[SDATA][8] , 
        \proc_out[SDATA][7] , \proc_out[SDATA][6] , \proc_out[SDATA][5] , 
        \proc_out[SDATA][4] , \proc_out[SDATA][3] , \proc_out[SDATA][2] , 
        \proc_out[SDATA][1] , \proc_out[SDATA][0] }), .spm_in({
        \spm_in[SCMDACCEPT] , \spm_in[SRESP] , \spm_in[SDATA][63] , 
        \spm_in[SDATA][62] , \spm_in[SDATA][61] , \spm_in[SDATA][60] , 
        \spm_in[SDATA][59] , \spm_in[SDATA][58] , \spm_in[SDATA][57] , 
        \spm_in[SDATA][56] , \spm_in[SDATA][55] , \spm_in[SDATA][54] , 
        \spm_in[SDATA][53] , \spm_in[SDATA][52] , \spm_in[SDATA][51] , 
        \spm_in[SDATA][50] , \spm_in[SDATA][49] , \spm_in[SDATA][48] , 
        \spm_in[SDATA][47] , \spm_in[SDATA][46] , \spm_in[SDATA][45] , 
        \spm_in[SDATA][44] , \spm_in[SDATA][43] , \spm_in[SDATA][42] , 
        \spm_in[SDATA][41] , \spm_in[SDATA][40] , \spm_in[SDATA][39] , 
        \spm_in[SDATA][38] , \spm_in[SDATA][37] , \spm_in[SDATA][36] , 
        \spm_in[SDATA][35] , \spm_in[SDATA][34] , \spm_in[SDATA][33] , 
        \spm_in[SDATA][32] , \spm_in[SDATA][31] , \spm_in[SDATA][30] , 
        \spm_in[SDATA][29] , \spm_in[SDATA][28] , \spm_in[SDATA][27] , 
        \spm_in[SDATA][26] , \spm_in[SDATA][25] , \spm_in[SDATA][24] , 
        \spm_in[SDATA][23] , \spm_in[SDATA][22] , \spm_in[SDATA][21] , 
        \spm_in[SDATA][20] , \spm_in[SDATA][19] , \spm_in[SDATA][18] , 
        \spm_in[SDATA][17] , \spm_in[SDATA][16] , \spm_in[SDATA][15] , 
        \spm_in[SDATA][14] , \spm_in[SDATA][13] , \spm_in[SDATA][12] , 
        \spm_in[SDATA][11] , \spm_in[SDATA][10] , \spm_in[SDATA][9] , 
        \spm_in[SDATA][8] , \spm_in[SDATA][7] , \spm_in[SDATA][6] , 
        \spm_in[SDATA][5] , \spm_in[SDATA][4] , \spm_in[SDATA][3] , 
        \spm_in[SDATA][2] , \spm_in[SDATA][1] , \spm_in[SDATA][0] }), 
        .spm_out({\spm_out[MCMD][1] , \spm_out[MCMD][0] , 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, \spm_out[MADDR][14] , \spm_out[MADDR][13] , 
        \spm_out[MADDR][12] , \spm_out[MADDR][11] , \spm_out[MADDR][10] , 
        \spm_out[MADDR][9] , \spm_out[MADDR][8] , \spm_out[MADDR][7] , 
        \spm_out[MADDR][6] , \spm_out[MADDR][5] , \spm_out[MADDR][4] , 
        \spm_out[MADDR][3] , \spm_out[MADDR][2] , \spm_out[MADDR][1] , 
        \spm_out[MADDR][0] , \spm_out[MDATA][63] , \spm_out[MDATA][62] , 
        \spm_out[MDATA][61] , \spm_out[MDATA][60] , \spm_out[MDATA][59] , 
        \spm_out[MDATA][58] , \spm_out[MDATA][57] , \spm_out[MDATA][56] , 
        \spm_out[MDATA][55] , \spm_out[MDATA][54] , \spm_out[MDATA][53] , 
        \spm_out[MDATA][52] , \spm_out[MDATA][51] , \spm_out[MDATA][50] , 
        \spm_out[MDATA][49] , \spm_out[MDATA][48] , \spm_out[MDATA][47] , 
        \spm_out[MDATA][46] , \spm_out[MDATA][45] , \spm_out[MDATA][44] , 
        \spm_out[MDATA][43] , \spm_out[MDATA][42] , \spm_out[MDATA][41] , 
        \spm_out[MDATA][40] , \spm_out[MDATA][39] , \spm_out[MDATA][38] , 
        \spm_out[MDATA][37] , \spm_out[MDATA][36] , \spm_out[MDATA][35] , 
        \spm_out[MDATA][34] , \spm_out[MDATA][33] , \spm_out[MDATA][32] , 
        \spm_out[MDATA][31] , \spm_out[MDATA][30] , \spm_out[MDATA][29] , 
        \spm_out[MDATA][28] , \spm_out[MDATA][27] , \spm_out[MDATA][26] , 
        \spm_out[MDATA][25] , \spm_out[MDATA][24] , \spm_out[MDATA][23] , 
        \spm_out[MDATA][22] , \spm_out[MDATA][21] , \spm_out[MDATA][20] , 
        \spm_out[MDATA][19] , \spm_out[MDATA][18] , \spm_out[MDATA][17] , 
        \spm_out[MDATA][16] , \spm_out[MDATA][15] , \spm_out[MDATA][14] , 
        \spm_out[MDATA][13] , \spm_out[MDATA][12] , \spm_out[MDATA][11] , 
        \spm_out[MDATA][10] , \spm_out[MDATA][9] , \spm_out[MDATA][8] , 
        \spm_out[MDATA][7] , \spm_out[MDATA][6] , \spm_out[MDATA][5] , 
        \spm_out[MDATA][4] , \spm_out[MDATA][3] , \spm_out[MDATA][2] , 
        \spm_out[MDATA][1] , \spm_out[MDATA][0] }), .pkt_in(net_to_ip), 
        .pkt_out(ip_to_net) );
  noc_switch_2 r ( .preset(reset), .north_in_f({\north_in_f[REQ] , 
        \north_in_f[DATA][34] , \north_in_f[DATA][33] , \north_in_f[DATA][32] , 
        \north_in_f[DATA][31] , \north_in_f[DATA][30] , \north_in_f[DATA][29] , 
        \north_in_f[DATA][28] , \north_in_f[DATA][27] , \north_in_f[DATA][26] , 
        \north_in_f[DATA][25] , \north_in_f[DATA][24] , \north_in_f[DATA][23] , 
        \north_in_f[DATA][22] , \north_in_f[DATA][21] , \north_in_f[DATA][20] , 
        \north_in_f[DATA][19] , \north_in_f[DATA][18] , \north_in_f[DATA][17] , 
        \north_in_f[DATA][16] , \north_in_f[DATA][15] , \north_in_f[DATA][14] , 
        \north_in_f[DATA][13] , \north_in_f[DATA][12] , \north_in_f[DATA][11] , 
        \north_in_f[DATA][10] , \north_in_f[DATA][9] , \north_in_f[DATA][8] , 
        \north_in_f[DATA][7] , \north_in_f[DATA][6] , \north_in_f[DATA][5] , 
        \north_in_f[DATA][4] , \north_in_f[DATA][3] , \north_in_f[DATA][2] , 
        \north_in_f[DATA][1] , \north_in_f[DATA][0] }), .north_in_b(
        \north_in_b[ACK] ), .east_in_f({\east_in_f[REQ] , 
        \east_in_f[DATA][34] , \east_in_f[DATA][33] , \east_in_f[DATA][32] , 
        \east_in_f[DATA][31] , \east_in_f[DATA][30] , \east_in_f[DATA][29] , 
        \east_in_f[DATA][28] , \east_in_f[DATA][27] , \east_in_f[DATA][26] , 
        \east_in_f[DATA][25] , \east_in_f[DATA][24] , \east_in_f[DATA][23] , 
        \east_in_f[DATA][22] , \east_in_f[DATA][21] , \east_in_f[DATA][20] , 
        \east_in_f[DATA][19] , \east_in_f[DATA][18] , \east_in_f[DATA][17] , 
        \east_in_f[DATA][16] , \east_in_f[DATA][15] , \east_in_f[DATA][14] , 
        \east_in_f[DATA][13] , \east_in_f[DATA][12] , \east_in_f[DATA][11] , 
        \east_in_f[DATA][10] , \east_in_f[DATA][9] , \east_in_f[DATA][8] , 
        \east_in_f[DATA][7] , \east_in_f[DATA][6] , \east_in_f[DATA][5] , 
        \east_in_f[DATA][4] , \east_in_f[DATA][3] , \east_in_f[DATA][2] , 
        \east_in_f[DATA][1] , \east_in_f[DATA][0] }), .east_in_b(
        \east_in_b[ACK] ), .south_in_f({\south_in_f[REQ] , 
        \south_in_f[DATA][34] , \south_in_f[DATA][33] , \south_in_f[DATA][32] , 
        \south_in_f[DATA][31] , \south_in_f[DATA][30] , \south_in_f[DATA][29] , 
        \south_in_f[DATA][28] , \south_in_f[DATA][27] , \south_in_f[DATA][26] , 
        \south_in_f[DATA][25] , \south_in_f[DATA][24] , \south_in_f[DATA][23] , 
        \south_in_f[DATA][22] , \south_in_f[DATA][21] , \south_in_f[DATA][20] , 
        \south_in_f[DATA][19] , \south_in_f[DATA][18] , \south_in_f[DATA][17] , 
        \south_in_f[DATA][16] , \south_in_f[DATA][15] , \south_in_f[DATA][14] , 
        \south_in_f[DATA][13] , \south_in_f[DATA][12] , \south_in_f[DATA][11] , 
        \south_in_f[DATA][10] , \south_in_f[DATA][9] , \south_in_f[DATA][8] , 
        \south_in_f[DATA][7] , \south_in_f[DATA][6] , \south_in_f[DATA][5] , 
        \south_in_f[DATA][4] , \south_in_f[DATA][3] , \south_in_f[DATA][2] , 
        \south_in_f[DATA][1] , \south_in_f[DATA][0] }), .south_in_b(
        \south_in_b[ACK] ), .west_in_f({\west_in_f[REQ] , 
        \west_in_f[DATA][34] , \west_in_f[DATA][33] , \west_in_f[DATA][32] , 
        \west_in_f[DATA][31] , \west_in_f[DATA][30] , \west_in_f[DATA][29] , 
        \west_in_f[DATA][28] , \west_in_f[DATA][27] , \west_in_f[DATA][26] , 
        \west_in_f[DATA][25] , \west_in_f[DATA][24] , \west_in_f[DATA][23] , 
        \west_in_f[DATA][22] , \west_in_f[DATA][21] , \west_in_f[DATA][20] , 
        \west_in_f[DATA][19] , \west_in_f[DATA][18] , \west_in_f[DATA][17] , 
        \west_in_f[DATA][16] , \west_in_f[DATA][15] , \west_in_f[DATA][14] , 
        \west_in_f[DATA][13] , \west_in_f[DATA][12] , \west_in_f[DATA][11] , 
        \west_in_f[DATA][10] , \west_in_f[DATA][9] , \west_in_f[DATA][8] , 
        \west_in_f[DATA][7] , \west_in_f[DATA][6] , \west_in_f[DATA][5] , 
        \west_in_f[DATA][4] , \west_in_f[DATA][3] , \west_in_f[DATA][2] , 
        \west_in_f[DATA][1] , \west_in_f[DATA][0] }), .west_in_b(
        \west_in_b[ACK] ), .resource_in_f({\ip_to_net_f[REQ] , ip_to_net}), 
        .north_out_f({\north_out_f[REQ] , \north_out_f[DATA][34] , 
        \north_out_f[DATA][33] , \north_out_f[DATA][32] , 
        \north_out_f[DATA][31] , \north_out_f[DATA][30] , 
        \north_out_f[DATA][29] , \north_out_f[DATA][28] , 
        \north_out_f[DATA][27] , \north_out_f[DATA][26] , 
        \north_out_f[DATA][25] , \north_out_f[DATA][24] , 
        \north_out_f[DATA][23] , \north_out_f[DATA][22] , 
        \north_out_f[DATA][21] , \north_out_f[DATA][20] , 
        \north_out_f[DATA][19] , \north_out_f[DATA][18] , 
        \north_out_f[DATA][17] , \north_out_f[DATA][16] , 
        \north_out_f[DATA][15] , \north_out_f[DATA][14] , 
        \north_out_f[DATA][13] , \north_out_f[DATA][12] , 
        \north_out_f[DATA][11] , \north_out_f[DATA][10] , 
        \north_out_f[DATA][9] , \north_out_f[DATA][8] , \north_out_f[DATA][7] , 
        \north_out_f[DATA][6] , \north_out_f[DATA][5] , \north_out_f[DATA][4] , 
        \north_out_f[DATA][3] , \north_out_f[DATA][2] , \north_out_f[DATA][1] , 
        \north_out_f[DATA][0] }), .north_out_b(\north_out_b[ACK] ), 
        .east_out_f({\east_out_f[REQ] , \east_out_f[DATA][34] , 
        \east_out_f[DATA][33] , \east_out_f[DATA][32] , \east_out_f[DATA][31] , 
        \east_out_f[DATA][30] , \east_out_f[DATA][29] , \east_out_f[DATA][28] , 
        \east_out_f[DATA][27] , \east_out_f[DATA][26] , \east_out_f[DATA][25] , 
        \east_out_f[DATA][24] , \east_out_f[DATA][23] , \east_out_f[DATA][22] , 
        \east_out_f[DATA][21] , \east_out_f[DATA][20] , \east_out_f[DATA][19] , 
        \east_out_f[DATA][18] , \east_out_f[DATA][17] , \east_out_f[DATA][16] , 
        \east_out_f[DATA][15] , \east_out_f[DATA][14] , \east_out_f[DATA][13] , 
        \east_out_f[DATA][12] , \east_out_f[DATA][11] , \east_out_f[DATA][10] , 
        \east_out_f[DATA][9] , \east_out_f[DATA][8] , \east_out_f[DATA][7] , 
        \east_out_f[DATA][6] , \east_out_f[DATA][5] , \east_out_f[DATA][4] , 
        \east_out_f[DATA][3] , \east_out_f[DATA][2] , \east_out_f[DATA][1] , 
        \east_out_f[DATA][0] }), .east_out_b(\east_out_b[ACK] ), .south_out_f(
        {\south_out_f[REQ] , \south_out_f[DATA][34] , \south_out_f[DATA][33] , 
        \south_out_f[DATA][32] , \south_out_f[DATA][31] , 
        \south_out_f[DATA][30] , \south_out_f[DATA][29] , 
        \south_out_f[DATA][28] , \south_out_f[DATA][27] , 
        \south_out_f[DATA][26] , \south_out_f[DATA][25] , 
        \south_out_f[DATA][24] , \south_out_f[DATA][23] , 
        \south_out_f[DATA][22] , \south_out_f[DATA][21] , 
        \south_out_f[DATA][20] , \south_out_f[DATA][19] , 
        \south_out_f[DATA][18] , \south_out_f[DATA][17] , 
        \south_out_f[DATA][16] , \south_out_f[DATA][15] , 
        \south_out_f[DATA][14] , \south_out_f[DATA][13] , 
        \south_out_f[DATA][12] , \south_out_f[DATA][11] , 
        \south_out_f[DATA][10] , \south_out_f[DATA][9] , 
        \south_out_f[DATA][8] , \south_out_f[DATA][7] , \south_out_f[DATA][6] , 
        \south_out_f[DATA][5] , \south_out_f[DATA][4] , \south_out_f[DATA][3] , 
        \south_out_f[DATA][2] , \south_out_f[DATA][1] , \south_out_f[DATA][0] }), .south_out_b(\south_out_b[ACK] ), .west_out_f({\west_out_f[REQ] , 
        \west_out_f[DATA][34] , \west_out_f[DATA][33] , \west_out_f[DATA][32] , 
        \west_out_f[DATA][31] , \west_out_f[DATA][30] , \west_out_f[DATA][29] , 
        \west_out_f[DATA][28] , \west_out_f[DATA][27] , \west_out_f[DATA][26] , 
        \west_out_f[DATA][25] , \west_out_f[DATA][24] , \west_out_f[DATA][23] , 
        \west_out_f[DATA][22] , \west_out_f[DATA][21] , \west_out_f[DATA][20] , 
        \west_out_f[DATA][19] , \west_out_f[DATA][18] , \west_out_f[DATA][17] , 
        \west_out_f[DATA][16] , \west_out_f[DATA][15] , \west_out_f[DATA][14] , 
        \west_out_f[DATA][13] , \west_out_f[DATA][12] , \west_out_f[DATA][11] , 
        \west_out_f[DATA][10] , \west_out_f[DATA][9] , \west_out_f[DATA][8] , 
        \west_out_f[DATA][7] , \west_out_f[DATA][6] , \west_out_f[DATA][5] , 
        \west_out_f[DATA][4] , \west_out_f[DATA][3] , \west_out_f[DATA][2] , 
        \west_out_f[DATA][1] , \west_out_f[DATA][0] }), .west_out_b(
        \west_out_b[ACK] ), .resource_out_f({SYNOPSYS_UNCONNECTED__17, 
        net_to_ip}), .resource_out_b(n9) );
  HS65_LS_DFPRQNX9 half_clk_reg ( .D(n11), .CP(n_clk), .RN(n8), .QN(n11) );
  HS65_LS_IVX9 I_2 ( .A(n4), .Z(\ip_to_net_f[REQ] ) );
  HS65_LH_IVX2 I_1 ( .A(n10), .Z(del_half_clk0) );
  HS65_LS_IVX9 U3 ( .A(n11), .Z(n10) );
  HS65_LH_IVX2 U4 ( .A(n1), .Z(n3) );
  HS65_LS_IVX106 U5 ( .A(del_half_clk0), .Z(n1) );
  HS65_LS_BFX9 U6 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U7 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U8 ( .A(n7), .Z(n6) );
  HS65_LS_BFX9 U9 ( .A(n3), .Z(n7) );
  HS65_LS_IVX9 U10 ( .A(reset), .Z(n8) );
  HS65_LS_IVX9 U11 ( .A(del_half_clk0), .Z(n9) );
endmodule


module counter_WIDTH3_1 ( clk, reset, enable, cnt );
  output [2:0] cnt;
  input clk, reset, enable;
  wire   n1, n2, n3, n4, n5, n8, n9, n10, n11;

  HS65_LS_DFPRQX9 \reg_reg[0]  ( .D(n5), .CP(clk), .RN(n1), .Q(cnt[0]) );
  HS65_LS_DFPRQX9 \reg_reg[2]  ( .D(n8), .CP(clk), .RN(n1), .Q(cnt[2]) );
  HS65_LS_DFPRQX9 \reg_reg[1]  ( .D(n9), .CP(clk), .RN(n1), .Q(cnt[1]) );
  HS65_LS_IVX9 U3 ( .A(reset), .Z(n1) );
  HS65_LS_OAI32X5 U4 ( .A(n4), .B(n11), .C(n2), .D(enable), .E(n3), .Z(n8) );
  HS65_LS_NAND2X7 U5 ( .A(enable), .B(n3), .Z(n11) );
  HS65_LS_OAI32X5 U6 ( .A(n2), .B(cnt[1]), .C(n11), .D(n10), .E(n4), .Z(n9) );
  HS65_LS_OA12X9 U7 ( .A(cnt[0]), .B(cnt[2]), .C(enable), .Z(n10) );
  HS65_LS_OAI22X6 U8 ( .A(enable), .B(n2), .C(cnt[0]), .D(n11), .Z(n5) );
  HS65_LS_IVX9 U9 ( .A(cnt[0]), .Z(n2) );
  HS65_LS_IVX9 U10 ( .A(cnt[1]), .Z(n4) );
  HS65_LS_IVX9 U11 ( .A(cnt[2]), .Z(n3) );
endmodule


module bram_DATA16_ADDR2_2 ( clk, reset, rd_addr, wr_addr, wr_data, wr_ena, 
        rd_data );
  input [1:0] rd_addr;
  input [1:0] wr_addr;
  input [15:0] wr_data;
  output [15:0] rd_data;
  input clk, reset, wr_ena;
  wire   \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] ,
         \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][15] , \mem[1][14] , \mem[1][13] ,
         \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] , \mem[1][8] ,
         \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] ,
         \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][15] , \mem[0][14] ,
         \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] ,
         \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] ,
         \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, n1,
         n2, n3, n4, n5, n6, n7, n8, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162;

  HS65_LS_DFPRQX9 \mem_reg[3][15]  ( .D(n91), .CP(clk), .RN(n1), .Q(
        \mem[3][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][14]  ( .D(n92), .CP(clk), .RN(n1), .Q(
        \mem[3][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][13]  ( .D(n93), .CP(clk), .RN(n1), .Q(
        \mem[3][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][12]  ( .D(n94), .CP(clk), .RN(n1), .Q(
        \mem[3][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][11]  ( .D(n95), .CP(clk), .RN(n1), .Q(
        \mem[3][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][10]  ( .D(n96), .CP(clk), .RN(n1), .Q(
        \mem[3][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][9]  ( .D(n97), .CP(clk), .RN(n1), .Q(\mem[3][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][8]  ( .D(n98), .CP(clk), .RN(n1), .Q(\mem[3][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][7]  ( .D(n99), .CP(clk), .RN(n1), .Q(\mem[3][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][6]  ( .D(n100), .CP(clk), .RN(n1), .Q(
        \mem[3][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][5]  ( .D(n101), .CP(clk), .RN(n1), .Q(
        \mem[3][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][4]  ( .D(n102), .CP(clk), .RN(n1), .Q(
        \mem[3][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][3]  ( .D(n103), .CP(clk), .RN(n1), .Q(
        \mem[3][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][2]  ( .D(n104), .CP(clk), .RN(n2), .Q(
        \mem[3][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][1]  ( .D(n105), .CP(clk), .RN(n2), .Q(
        \mem[3][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][0]  ( .D(n106), .CP(clk), .RN(n2), .Q(
        \mem[3][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][15]  ( .D(n107), .CP(clk), .RN(n2), .Q(
        \mem[2][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][14]  ( .D(n108), .CP(clk), .RN(n2), .Q(
        \mem[2][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][13]  ( .D(n109), .CP(clk), .RN(n2), .Q(
        \mem[2][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][12]  ( .D(n110), .CP(clk), .RN(n2), .Q(
        \mem[2][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][11]  ( .D(n111), .CP(clk), .RN(n2), .Q(
        \mem[2][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][10]  ( .D(n112), .CP(clk), .RN(n2), .Q(
        \mem[2][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][9]  ( .D(n113), .CP(clk), .RN(n2), .Q(
        \mem[2][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][8]  ( .D(n114), .CP(clk), .RN(n2), .Q(
        \mem[2][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][7]  ( .D(n115), .CP(clk), .RN(n2), .Q(
        \mem[2][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][6]  ( .D(n116), .CP(clk), .RN(n2), .Q(
        \mem[2][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][5]  ( .D(n117), .CP(clk), .RN(n3), .Q(
        \mem[2][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][4]  ( .D(n118), .CP(clk), .RN(n3), .Q(
        \mem[2][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][3]  ( .D(n119), .CP(clk), .RN(n3), .Q(
        \mem[2][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][2]  ( .D(n120), .CP(clk), .RN(n3), .Q(
        \mem[2][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][1]  ( .D(n121), .CP(clk), .RN(n3), .Q(
        \mem[2][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][0]  ( .D(n122), .CP(clk), .RN(n3), .Q(
        \mem[2][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][15]  ( .D(n123), .CP(clk), .RN(n3), .Q(
        \mem[1][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][14]  ( .D(n124), .CP(clk), .RN(n3), .Q(
        \mem[1][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][13]  ( .D(n125), .CP(clk), .RN(n3), .Q(
        \mem[1][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][12]  ( .D(n126), .CP(clk), .RN(n3), .Q(
        \mem[1][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][11]  ( .D(n127), .CP(clk), .RN(n3), .Q(
        \mem[1][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][10]  ( .D(n128), .CP(clk), .RN(n3), .Q(
        \mem[1][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][9]  ( .D(n129), .CP(clk), .RN(n3), .Q(
        \mem[1][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][8]  ( .D(n130), .CP(clk), .RN(n4), .Q(
        \mem[1][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][7]  ( .D(n131), .CP(clk), .RN(n4), .Q(
        \mem[1][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][6]  ( .D(n132), .CP(clk), .RN(n4), .Q(
        \mem[1][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][5]  ( .D(n133), .CP(clk), .RN(n4), .Q(
        \mem[1][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][4]  ( .D(n134), .CP(clk), .RN(n4), .Q(
        \mem[1][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][3]  ( .D(n135), .CP(clk), .RN(n4), .Q(
        \mem[1][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][2]  ( .D(n136), .CP(clk), .RN(n4), .Q(
        \mem[1][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][1]  ( .D(n137), .CP(clk), .RN(n4), .Q(
        \mem[1][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][0]  ( .D(n138), .CP(clk), .RN(n4), .Q(
        \mem[1][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][15]  ( .D(n139), .CP(clk), .RN(n4), .Q(
        \mem[0][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][14]  ( .D(n140), .CP(clk), .RN(n4), .Q(
        \mem[0][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][13]  ( .D(n141), .CP(clk), .RN(n4), .Q(
        \mem[0][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][12]  ( .D(n142), .CP(clk), .RN(n4), .Q(
        \mem[0][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][11]  ( .D(n143), .CP(clk), .RN(n5), .Q(
        \mem[0][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][10]  ( .D(n144), .CP(clk), .RN(n5), .Q(
        \mem[0][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][9]  ( .D(n145), .CP(clk), .RN(n5), .Q(
        \mem[0][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][8]  ( .D(n146), .CP(clk), .RN(n5), .Q(
        \mem[0][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][7]  ( .D(n147), .CP(clk), .RN(n5), .Q(
        \mem[0][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][6]  ( .D(n148), .CP(clk), .RN(n5), .Q(
        \mem[0][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][5]  ( .D(n149), .CP(clk), .RN(n5), .Q(
        \mem[0][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][4]  ( .D(n150), .CP(clk), .RN(n5), .Q(
        \mem[0][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][3]  ( .D(n151), .CP(clk), .RN(n5), .Q(
        \mem[0][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][2]  ( .D(n152), .CP(clk), .RN(n5), .Q(
        \mem[0][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][1]  ( .D(n153), .CP(clk), .RN(n5), .Q(
        \mem[0][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][0]  ( .D(n154), .CP(clk), .RN(n5), .Q(
        \mem[0][0] ) );
  HS65_LS_DFPRQX9 \rd_data_reg[15]  ( .D(N17), .CP(clk), .RN(n5), .Q(
        rd_data[15]) );
  HS65_LS_DFPRQX9 \rd_data_reg[14]  ( .D(N18), .CP(clk), .RN(n6), .Q(
        rd_data[14]) );
  HS65_LS_DFPRQX9 \rd_data_reg[13]  ( .D(N19), .CP(clk), .RN(n6), .Q(
        rd_data[13]) );
  HS65_LS_DFPRQX9 \rd_data_reg[12]  ( .D(N20), .CP(clk), .RN(n6), .Q(
        rd_data[12]) );
  HS65_LS_DFPRQX9 \rd_data_reg[11]  ( .D(N21), .CP(clk), .RN(n6), .Q(
        rd_data[11]) );
  HS65_LS_DFPRQX9 \rd_data_reg[10]  ( .D(N22), .CP(clk), .RN(n6), .Q(
        rd_data[10]) );
  HS65_LS_DFPRQX9 \rd_data_reg[9]  ( .D(N23), .CP(clk), .RN(n6), .Q(rd_data[9]) );
  HS65_LS_DFPRQX9 \rd_data_reg[8]  ( .D(N24), .CP(clk), .RN(n6), .Q(rd_data[8]) );
  HS65_LS_DFPRQX9 \rd_data_reg[7]  ( .D(N25), .CP(clk), .RN(n6), .Q(rd_data[7]) );
  HS65_LS_DFPRQX9 \rd_data_reg[6]  ( .D(N26), .CP(clk), .RN(n6), .Q(rd_data[6]) );
  HS65_LS_DFPRQX9 \rd_data_reg[5]  ( .D(N27), .CP(clk), .RN(n6), .Q(rd_data[5]) );
  HS65_LS_DFPRQX9 \rd_data_reg[4]  ( .D(N28), .CP(clk), .RN(n6), .Q(rd_data[4]) );
  HS65_LS_DFPRQX9 \rd_data_reg[3]  ( .D(N29), .CP(clk), .RN(n6), .Q(rd_data[3]) );
  HS65_LS_DFPRQX9 \rd_data_reg[2]  ( .D(N30), .CP(clk), .RN(n6), .Q(rd_data[2]) );
  HS65_LS_DFPRQX9 \rd_data_reg[1]  ( .D(N31), .CP(clk), .RN(n7), .Q(rd_data[1]) );
  HS65_LS_DFPRQX9 \rd_data_reg[0]  ( .D(N32), .CP(clk), .RN(n7), .Q(rd_data[0]) );
  HS65_LS_BFX9 U3 ( .A(n81), .Z(n4) );
  HS65_LS_BFX9 U4 ( .A(n81), .Z(n3) );
  HS65_LS_BFX9 U5 ( .A(n81), .Z(n2) );
  HS65_LS_BFX9 U6 ( .A(n83), .Z(n81) );
  HS65_LS_BFX9 U7 ( .A(n8), .Z(n6) );
  HS65_LS_BFX9 U8 ( .A(n8), .Z(n5) );
  HS65_LS_BFX9 U9 ( .A(n82), .Z(n1) );
  HS65_LS_BFX9 U10 ( .A(n83), .Z(n82) );
  HS65_LS_BFX9 U11 ( .A(n8), .Z(n7) );
  HS65_LS_BFX9 U12 ( .A(n83), .Z(n8) );
  HS65_LS_IVX9 U13 ( .A(reset), .Z(n83) );
  HS65_LS_IVX9 U14 ( .A(n161), .Z(n86) );
  HS65_LS_IVX9 U15 ( .A(n162), .Z(n87) );
  HS65_LS_NAND3X5 U16 ( .A(wr_ena), .B(n88), .C(wr_addr[0]), .Z(n161) );
  HS65_LS_IVX9 U17 ( .A(wr_addr[0]), .Z(n89) );
  HS65_LS_NAND3X5 U18 ( .A(n89), .B(n88), .C(wr_ena), .Z(n162) );
  HS65_LS_IVX9 U19 ( .A(n160), .Z(n85) );
  HS65_LS_IVX9 U20 ( .A(n159), .Z(n84) );
  HS65_LS_NAND3X5 U21 ( .A(wr_ena), .B(n89), .C(wr_addr[1]), .Z(n160) );
  HS65_LS_NOR2X6 U22 ( .A(n90), .B(rd_addr[1]), .Z(n157) );
  HS65_LS_NOR2X6 U23 ( .A(rd_addr[0]), .B(rd_addr[1]), .Z(n158) );
  HS65_LS_IVX9 U24 ( .A(wr_addr[1]), .Z(n88) );
  HS65_LS_NAND3X5 U25 ( .A(wr_addr[0]), .B(wr_ena), .C(wr_addr[1]), .Z(n159)
         );
  HS65_LS_AND2X4 U26 ( .A(rd_addr[1]), .B(n90), .Z(n156) );
  HS65_LS_IVX9 U27 ( .A(rd_addr[0]), .Z(n90) );
  HS65_LS_AND2X4 U28 ( .A(rd_addr[1]), .B(rd_addr[0]), .Z(n155) );
  HS65_LS_MX41X7 U29 ( .D0(n158), .S0(\mem[0][0] ), .D1(n157), .S1(\mem[1][0] ), .D2(n156), .S2(\mem[2][0] ), .D3(n155), .S3(\mem[3][0] ), .Z(N32) );
  HS65_LS_MX41X7 U30 ( .D0(n158), .S0(\mem[0][1] ), .D1(n157), .S1(\mem[1][1] ), .D2(n156), .S2(\mem[2][1] ), .D3(n155), .S3(\mem[3][1] ), .Z(N31) );
  HS65_LS_MX41X7 U31 ( .D0(n158), .S0(\mem[0][2] ), .D1(n157), .S1(\mem[1][2] ), .D2(n156), .S2(\mem[2][2] ), .D3(n155), .S3(\mem[3][2] ), .Z(N30) );
  HS65_LS_MX41X7 U32 ( .D0(n158), .S0(\mem[0][3] ), .D1(n157), .S1(\mem[1][3] ), .D2(n156), .S2(\mem[2][3] ), .D3(n155), .S3(\mem[3][3] ), .Z(N29) );
  HS65_LS_MX41X7 U33 ( .D0(n158), .S0(\mem[0][4] ), .D1(n157), .S1(\mem[1][4] ), .D2(n156), .S2(\mem[2][4] ), .D3(n155), .S3(\mem[3][4] ), .Z(N28) );
  HS65_LS_MX41X7 U34 ( .D0(n158), .S0(\mem[0][5] ), .D1(n157), .S1(\mem[1][5] ), .D2(n156), .S2(\mem[2][5] ), .D3(n155), .S3(\mem[3][5] ), .Z(N27) );
  HS65_LS_MX41X7 U35 ( .D0(n158), .S0(\mem[0][6] ), .D1(n157), .S1(\mem[1][6] ), .D2(n156), .S2(\mem[2][6] ), .D3(n155), .S3(\mem[3][6] ), .Z(N26) );
  HS65_LS_MX41X7 U36 ( .D0(n158), .S0(\mem[0][7] ), .D1(n157), .S1(\mem[1][7] ), .D2(n156), .S2(\mem[2][7] ), .D3(n155), .S3(\mem[3][7] ), .Z(N25) );
  HS65_LS_MX41X7 U37 ( .D0(n158), .S0(\mem[0][8] ), .D1(n157), .S1(\mem[1][8] ), .D2(n156), .S2(\mem[2][8] ), .D3(n155), .S3(\mem[3][8] ), .Z(N24) );
  HS65_LS_MX41X7 U38 ( .D0(n158), .S0(\mem[0][9] ), .D1(n157), .S1(\mem[1][9] ), .D2(n156), .S2(\mem[2][9] ), .D3(n155), .S3(\mem[3][9] ), .Z(N23) );
  HS65_LS_MX41X7 U39 ( .D0(n158), .S0(\mem[0][10] ), .D1(n157), .S1(
        \mem[1][10] ), .D2(n156), .S2(\mem[2][10] ), .D3(n155), .S3(
        \mem[3][10] ), .Z(N22) );
  HS65_LS_MX41X7 U40 ( .D0(n158), .S0(\mem[0][11] ), .D1(n157), .S1(
        \mem[1][11] ), .D2(n156), .S2(\mem[2][11] ), .D3(n155), .S3(
        \mem[3][11] ), .Z(N21) );
  HS65_LS_MX41X7 U41 ( .D0(n158), .S0(\mem[0][12] ), .D1(n157), .S1(
        \mem[1][12] ), .D2(n156), .S2(\mem[2][12] ), .D3(n155), .S3(
        \mem[3][12] ), .Z(N20) );
  HS65_LS_MX41X7 U42 ( .D0(n158), .S0(\mem[0][13] ), .D1(n157), .S1(
        \mem[1][13] ), .D2(n156), .S2(\mem[2][13] ), .D3(n155), .S3(
        \mem[3][13] ), .Z(N19) );
  HS65_LS_MX41X7 U43 ( .D0(n158), .S0(\mem[0][14] ), .D1(n157), .S1(
        \mem[1][14] ), .D2(n156), .S2(\mem[2][14] ), .D3(n155), .S3(
        \mem[3][14] ), .Z(N18) );
  HS65_LS_MX41X7 U44 ( .D0(n158), .S0(\mem[0][15] ), .D1(n157), .S1(
        \mem[1][15] ), .D2(n156), .S2(\mem[2][15] ), .D3(n155), .S3(
        \mem[3][15] ), .Z(N17) );
  HS65_LS_AO22X9 U45 ( .A(wr_data[0]), .B(n86), .C(n161), .D(\mem[1][0] ), .Z(
        n138) );
  HS65_LS_AO22X9 U46 ( .A(wr_data[1]), .B(n86), .C(n161), .D(\mem[1][1] ), .Z(
        n137) );
  HS65_LS_AO22X9 U47 ( .A(wr_data[2]), .B(n86), .C(n161), .D(\mem[1][2] ), .Z(
        n136) );
  HS65_LS_AO22X9 U48 ( .A(wr_data[3]), .B(n86), .C(n161), .D(\mem[1][3] ), .Z(
        n135) );
  HS65_LS_AO22X9 U49 ( .A(wr_data[4]), .B(n86), .C(n161), .D(\mem[1][4] ), .Z(
        n134) );
  HS65_LS_AO22X9 U50 ( .A(wr_data[5]), .B(n86), .C(n161), .D(\mem[1][5] ), .Z(
        n133) );
  HS65_LS_AO22X9 U51 ( .A(wr_data[6]), .B(n86), .C(n161), .D(\mem[1][6] ), .Z(
        n132) );
  HS65_LS_AO22X9 U52 ( .A(wr_data[7]), .B(n86), .C(n161), .D(\mem[1][7] ), .Z(
        n131) );
  HS65_LS_AO22X9 U53 ( .A(wr_data[8]), .B(n86), .C(n161), .D(\mem[1][8] ), .Z(
        n130) );
  HS65_LS_AO22X9 U54 ( .A(wr_data[9]), .B(n86), .C(n161), .D(\mem[1][9] ), .Z(
        n129) );
  HS65_LS_AO22X9 U55 ( .A(wr_data[10]), .B(n86), .C(n161), .D(\mem[1][10] ), 
        .Z(n128) );
  HS65_LS_AO22X9 U56 ( .A(wr_data[11]), .B(n86), .C(n161), .D(\mem[1][11] ), 
        .Z(n127) );
  HS65_LS_AO22X9 U57 ( .A(wr_data[12]), .B(n86), .C(n161), .D(\mem[1][12] ), 
        .Z(n126) );
  HS65_LS_AO22X9 U58 ( .A(wr_data[13]), .B(n86), .C(n161), .D(\mem[1][13] ), 
        .Z(n125) );
  HS65_LS_AO22X9 U59 ( .A(wr_data[14]), .B(n86), .C(n161), .D(\mem[1][14] ), 
        .Z(n124) );
  HS65_LS_AO22X9 U60 ( .A(wr_data[15]), .B(n86), .C(n161), .D(\mem[1][15] ), 
        .Z(n123) );
  HS65_LS_AO22X9 U61 ( .A(wr_data[0]), .B(n85), .C(n160), .D(\mem[2][0] ), .Z(
        n122) );
  HS65_LS_AO22X9 U62 ( .A(wr_data[1]), .B(n85), .C(n160), .D(\mem[2][1] ), .Z(
        n121) );
  HS65_LS_AO22X9 U63 ( .A(wr_data[2]), .B(n85), .C(n160), .D(\mem[2][2] ), .Z(
        n120) );
  HS65_LS_AO22X9 U64 ( .A(wr_data[3]), .B(n85), .C(n160), .D(\mem[2][3] ), .Z(
        n119) );
  HS65_LS_AO22X9 U65 ( .A(wr_data[4]), .B(n85), .C(n160), .D(\mem[2][4] ), .Z(
        n118) );
  HS65_LS_AO22X9 U66 ( .A(wr_data[5]), .B(n85), .C(n160), .D(\mem[2][5] ), .Z(
        n117) );
  HS65_LS_AO22X9 U67 ( .A(wr_data[6]), .B(n85), .C(n160), .D(\mem[2][6] ), .Z(
        n116) );
  HS65_LS_AO22X9 U68 ( .A(wr_data[7]), .B(n85), .C(n160), .D(\mem[2][7] ), .Z(
        n115) );
  HS65_LS_AO22X9 U69 ( .A(wr_data[8]), .B(n85), .C(n160), .D(\mem[2][8] ), .Z(
        n114) );
  HS65_LS_AO22X9 U70 ( .A(wr_data[9]), .B(n85), .C(n160), .D(\mem[2][9] ), .Z(
        n113) );
  HS65_LS_AO22X9 U71 ( .A(wr_data[10]), .B(n85), .C(n160), .D(\mem[2][10] ), 
        .Z(n112) );
  HS65_LS_AO22X9 U72 ( .A(wr_data[11]), .B(n85), .C(n160), .D(\mem[2][11] ), 
        .Z(n111) );
  HS65_LS_AO22X9 U73 ( .A(wr_data[12]), .B(n85), .C(n160), .D(\mem[2][12] ), 
        .Z(n110) );
  HS65_LS_AO22X9 U74 ( .A(wr_data[13]), .B(n85), .C(n160), .D(\mem[2][13] ), 
        .Z(n109) );
  HS65_LS_AO22X9 U75 ( .A(wr_data[14]), .B(n85), .C(n160), .D(\mem[2][14] ), 
        .Z(n108) );
  HS65_LS_AO22X9 U76 ( .A(wr_data[15]), .B(n85), .C(n160), .D(\mem[2][15] ), 
        .Z(n107) );
  HS65_LS_AO22X9 U77 ( .A(n87), .B(wr_data[0]), .C(n162), .D(\mem[0][0] ), .Z(
        n154) );
  HS65_LS_AO22X9 U78 ( .A(n87), .B(wr_data[1]), .C(n162), .D(\mem[0][1] ), .Z(
        n153) );
  HS65_LS_AO22X9 U79 ( .A(n87), .B(wr_data[2]), .C(n162), .D(\mem[0][2] ), .Z(
        n152) );
  HS65_LS_AO22X9 U80 ( .A(n87), .B(wr_data[3]), .C(n162), .D(\mem[0][3] ), .Z(
        n151) );
  HS65_LS_AO22X9 U81 ( .A(n87), .B(wr_data[4]), .C(n162), .D(\mem[0][4] ), .Z(
        n150) );
  HS65_LS_AO22X9 U82 ( .A(n87), .B(wr_data[5]), .C(n162), .D(\mem[0][5] ), .Z(
        n149) );
  HS65_LS_AO22X9 U83 ( .A(n87), .B(wr_data[6]), .C(n162), .D(\mem[0][6] ), .Z(
        n148) );
  HS65_LS_AO22X9 U84 ( .A(n87), .B(wr_data[7]), .C(n162), .D(\mem[0][7] ), .Z(
        n147) );
  HS65_LS_AO22X9 U85 ( .A(n87), .B(wr_data[8]), .C(n162), .D(\mem[0][8] ), .Z(
        n146) );
  HS65_LS_AO22X9 U86 ( .A(n87), .B(wr_data[9]), .C(n162), .D(\mem[0][9] ), .Z(
        n145) );
  HS65_LS_AO22X9 U87 ( .A(n87), .B(wr_data[10]), .C(n162), .D(\mem[0][10] ), 
        .Z(n144) );
  HS65_LS_AO22X9 U88 ( .A(n87), .B(wr_data[11]), .C(n162), .D(\mem[0][11] ), 
        .Z(n143) );
  HS65_LS_AO22X9 U89 ( .A(n87), .B(wr_data[12]), .C(n162), .D(\mem[0][12] ), 
        .Z(n142) );
  HS65_LS_AO22X9 U90 ( .A(n87), .B(wr_data[13]), .C(n162), .D(\mem[0][13] ), 
        .Z(n141) );
  HS65_LS_AO22X9 U91 ( .A(n87), .B(wr_data[14]), .C(n162), .D(\mem[0][14] ), 
        .Z(n140) );
  HS65_LS_AO22X9 U92 ( .A(n87), .B(wr_data[15]), .C(n162), .D(\mem[0][15] ), 
        .Z(n139) );
  HS65_LS_AO22X9 U93 ( .A(wr_data[0]), .B(n84), .C(n159), .D(\mem[3][0] ), .Z(
        n106) );
  HS65_LS_AO22X9 U94 ( .A(wr_data[1]), .B(n84), .C(n159), .D(\mem[3][1] ), .Z(
        n105) );
  HS65_LS_AO22X9 U95 ( .A(wr_data[2]), .B(n84), .C(n159), .D(\mem[3][2] ), .Z(
        n104) );
  HS65_LS_AO22X9 U96 ( .A(wr_data[3]), .B(n84), .C(n159), .D(\mem[3][3] ), .Z(
        n103) );
  HS65_LS_AO22X9 U97 ( .A(wr_data[4]), .B(n84), .C(n159), .D(\mem[3][4] ), .Z(
        n102) );
  HS65_LS_AO22X9 U98 ( .A(wr_data[5]), .B(n84), .C(n159), .D(\mem[3][5] ), .Z(
        n101) );
  HS65_LS_AO22X9 U99 ( .A(wr_data[6]), .B(n84), .C(n159), .D(\mem[3][6] ), .Z(
        n100) );
  HS65_LS_AO22X9 U100 ( .A(wr_data[7]), .B(n84), .C(n159), .D(\mem[3][7] ), 
        .Z(n99) );
  HS65_LS_AO22X9 U101 ( .A(wr_data[8]), .B(n84), .C(n159), .D(\mem[3][8] ), 
        .Z(n98) );
  HS65_LS_AO22X9 U102 ( .A(wr_data[9]), .B(n84), .C(n159), .D(\mem[3][9] ), 
        .Z(n97) );
  HS65_LS_AO22X9 U103 ( .A(wr_data[10]), .B(n84), .C(n159), .D(\mem[3][10] ), 
        .Z(n96) );
  HS65_LS_AO22X9 U104 ( .A(wr_data[11]), .B(n84), .C(n159), .D(\mem[3][11] ), 
        .Z(n95) );
  HS65_LS_AO22X9 U105 ( .A(wr_data[12]), .B(n84), .C(n159), .D(\mem[3][12] ), 
        .Z(n94) );
  HS65_LS_AO22X9 U106 ( .A(wr_data[13]), .B(n84), .C(n159), .D(\mem[3][13] ), 
        .Z(n93) );
  HS65_LS_AO22X9 U107 ( .A(wr_data[14]), .B(n84), .C(n159), .D(\mem[3][14] ), 
        .Z(n92) );
  HS65_LS_AO22X9 U108 ( .A(wr_data[15]), .B(n84), .C(n159), .D(\mem[3][15] ), 
        .Z(n91) );
endmodule


module bram_DATA32_ADDR2_1 ( clk, reset, rd_addr, wr_addr, wr_data, wr_ena, 
        rd_data );
  input [1:0] rd_addr;
  input [1:0] wr_addr;
  input [31:0] wr_data;
  output [31:0] rd_data;
  input clk, reset, wr_ena;
  wire   \mem[3][31] , \mem[3][30] , \mem[3][29] , \mem[3][28] , \mem[3][27] ,
         \mem[3][26] , \mem[3][25] , \mem[3][24] , \mem[3][23] , \mem[3][22] ,
         \mem[3][21] , \mem[3][20] , \mem[3][19] , \mem[3][18] , \mem[3][17] ,
         \mem[3][16] , \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] ,
         \mem[3][11] , \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] ,
         \mem[3][6] , \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] ,
         \mem[3][1] , \mem[3][0] , \mem[2][31] , \mem[2][30] , \mem[2][29] ,
         \mem[2][28] , \mem[2][27] , \mem[2][26] , \mem[2][25] , \mem[2][24] ,
         \mem[2][23] , \mem[2][22] , \mem[2][21] , \mem[2][20] , \mem[2][19] ,
         \mem[2][18] , \mem[2][17] , \mem[2][16] , \mem[2][15] , \mem[2][14] ,
         \mem[2][13] , \mem[2][12] , \mem[2][11] , \mem[2][10] , \mem[2][9] ,
         \mem[2][8] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][31] ,
         \mem[1][30] , \mem[1][29] , \mem[1][28] , \mem[1][27] , \mem[1][26] ,
         \mem[1][25] , \mem[1][24] , \mem[1][23] , \mem[1][22] , \mem[1][21] ,
         \mem[1][20] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][31] , \mem[0][30] , \mem[0][29] , \mem[0][28] ,
         \mem[0][27] , \mem[0][26] , \mem[0][25] , \mem[0][24] , \mem[0][23] ,
         \mem[0][22] , \mem[0][21] , \mem[0][20] , \mem[0][19] , \mem[0][18] ,
         \mem[0][17] , \mem[0][16] , \mem[0][15] , \mem[0][14] , \mem[0][13] ,
         \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] , \mem[0][8] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N17, N18, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36,
         N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327;

  HS65_LS_DFPRQX9 \mem_reg[3][31]  ( .D(n193), .CP(clk), .RN(n171), .Q(
        \mem[3][31] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][30]  ( .D(n194), .CP(clk), .RN(n171), .Q(
        \mem[3][30] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][29]  ( .D(n195), .CP(clk), .RN(n171), .Q(
        \mem[3][29] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][28]  ( .D(n196), .CP(clk), .RN(n171), .Q(
        \mem[3][28] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][27]  ( .D(n197), .CP(clk), .RN(n171), .Q(
        \mem[3][27] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][26]  ( .D(n198), .CP(clk), .RN(n171), .Q(
        \mem[3][26] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][25]  ( .D(n199), .CP(clk), .RN(n171), .Q(
        \mem[3][25] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][24]  ( .D(n200), .CP(clk), .RN(n171), .Q(
        \mem[3][24] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][23]  ( .D(n201), .CP(clk), .RN(n171), .Q(
        \mem[3][23] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][22]  ( .D(n202), .CP(clk), .RN(n171), .Q(
        \mem[3][22] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][21]  ( .D(n203), .CP(clk), .RN(n171), .Q(
        \mem[3][21] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][20]  ( .D(n204), .CP(clk), .RN(n171), .Q(
        \mem[3][20] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][19]  ( .D(n205), .CP(clk), .RN(n171), .Q(
        \mem[3][19] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][18]  ( .D(n206), .CP(clk), .RN(n172), .Q(
        \mem[3][18] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][17]  ( .D(n207), .CP(clk), .RN(n172), .Q(
        \mem[3][17] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][16]  ( .D(n208), .CP(clk), .RN(n172), .Q(
        \mem[3][16] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][15]  ( .D(n209), .CP(clk), .RN(n172), .Q(
        \mem[3][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][14]  ( .D(n210), .CP(clk), .RN(n172), .Q(
        \mem[3][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][13]  ( .D(n211), .CP(clk), .RN(n172), .Q(
        \mem[3][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][12]  ( .D(n212), .CP(clk), .RN(n172), .Q(
        \mem[3][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][11]  ( .D(n213), .CP(clk), .RN(n172), .Q(
        \mem[3][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][10]  ( .D(n214), .CP(clk), .RN(n172), .Q(
        \mem[3][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][9]  ( .D(n215), .CP(clk), .RN(n172), .Q(
        \mem[3][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][8]  ( .D(n216), .CP(clk), .RN(n172), .Q(
        \mem[3][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][7]  ( .D(n217), .CP(clk), .RN(n172), .Q(
        \mem[3][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][6]  ( .D(n218), .CP(clk), .RN(n172), .Q(
        \mem[3][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][5]  ( .D(n219), .CP(clk), .RN(n173), .Q(
        \mem[3][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][4]  ( .D(n220), .CP(clk), .RN(n173), .Q(
        \mem[3][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][3]  ( .D(n221), .CP(clk), .RN(n173), .Q(
        \mem[3][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][2]  ( .D(n222), .CP(clk), .RN(n173), .Q(
        \mem[3][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][1]  ( .D(n223), .CP(clk), .RN(n173), .Q(
        \mem[3][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][0]  ( .D(n224), .CP(clk), .RN(n173), .Q(
        \mem[3][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][31]  ( .D(n225), .CP(clk), .RN(n173), .Q(
        \mem[2][31] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][30]  ( .D(n226), .CP(clk), .RN(n173), .Q(
        \mem[2][30] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][29]  ( .D(n227), .CP(clk), .RN(n173), .Q(
        \mem[2][29] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][28]  ( .D(n228), .CP(clk), .RN(n173), .Q(
        \mem[2][28] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][27]  ( .D(n229), .CP(clk), .RN(n173), .Q(
        \mem[2][27] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][26]  ( .D(n230), .CP(clk), .RN(n173), .Q(
        \mem[2][26] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][25]  ( .D(n231), .CP(clk), .RN(n173), .Q(
        \mem[2][25] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][24]  ( .D(n232), .CP(clk), .RN(n174), .Q(
        \mem[2][24] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][23]  ( .D(n233), .CP(clk), .RN(n174), .Q(
        \mem[2][23] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][22]  ( .D(n234), .CP(clk), .RN(n174), .Q(
        \mem[2][22] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][21]  ( .D(n235), .CP(clk), .RN(n174), .Q(
        \mem[2][21] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][20]  ( .D(n236), .CP(clk), .RN(n174), .Q(
        \mem[2][20] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][19]  ( .D(n237), .CP(clk), .RN(n174), .Q(
        \mem[2][19] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][18]  ( .D(n238), .CP(clk), .RN(n174), .Q(
        \mem[2][18] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][17]  ( .D(n239), .CP(clk), .RN(n174), .Q(
        \mem[2][17] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][16]  ( .D(n240), .CP(clk), .RN(n174), .Q(
        \mem[2][16] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][15]  ( .D(n241), .CP(clk), .RN(n174), .Q(
        \mem[2][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][14]  ( .D(n242), .CP(clk), .RN(n174), .Q(
        \mem[2][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][13]  ( .D(n243), .CP(clk), .RN(n174), .Q(
        \mem[2][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][12]  ( .D(n244), .CP(clk), .RN(n174), .Q(
        \mem[2][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][11]  ( .D(n245), .CP(clk), .RN(n175), .Q(
        \mem[2][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][10]  ( .D(n246), .CP(clk), .RN(n175), .Q(
        \mem[2][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][9]  ( .D(n247), .CP(clk), .RN(n175), .Q(
        \mem[2][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][8]  ( .D(n248), .CP(clk), .RN(n175), .Q(
        \mem[2][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][7]  ( .D(n249), .CP(clk), .RN(n175), .Q(
        \mem[2][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][6]  ( .D(n250), .CP(clk), .RN(n175), .Q(
        \mem[2][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][5]  ( .D(n251), .CP(clk), .RN(n175), .Q(
        \mem[2][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][4]  ( .D(n252), .CP(clk), .RN(n175), .Q(
        \mem[2][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][3]  ( .D(n253), .CP(clk), .RN(n175), .Q(
        \mem[2][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][2]  ( .D(n254), .CP(clk), .RN(n175), .Q(
        \mem[2][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][1]  ( .D(n255), .CP(clk), .RN(n175), .Q(
        \mem[2][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][0]  ( .D(n256), .CP(clk), .RN(n175), .Q(
        \mem[2][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][31]  ( .D(n257), .CP(clk), .RN(n175), .Q(
        \mem[1][31] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][30]  ( .D(n258), .CP(clk), .RN(n176), .Q(
        \mem[1][30] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][29]  ( .D(n259), .CP(clk), .RN(n176), .Q(
        \mem[1][29] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][28]  ( .D(n260), .CP(clk), .RN(n176), .Q(
        \mem[1][28] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][27]  ( .D(n261), .CP(clk), .RN(n176), .Q(
        \mem[1][27] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][26]  ( .D(n262), .CP(clk), .RN(n176), .Q(
        \mem[1][26] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][25]  ( .D(n263), .CP(clk), .RN(n176), .Q(
        \mem[1][25] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][24]  ( .D(n264), .CP(clk), .RN(n176), .Q(
        \mem[1][24] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][23]  ( .D(n265), .CP(clk), .RN(n176), .Q(
        \mem[1][23] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][22]  ( .D(n266), .CP(clk), .RN(n176), .Q(
        \mem[1][22] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][21]  ( .D(n267), .CP(clk), .RN(n176), .Q(
        \mem[1][21] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][20]  ( .D(n268), .CP(clk), .RN(n176), .Q(
        \mem[1][20] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][19]  ( .D(n269), .CP(clk), .RN(n176), .Q(
        \mem[1][19] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][18]  ( .D(n270), .CP(clk), .RN(n176), .Q(
        \mem[1][18] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][17]  ( .D(n271), .CP(clk), .RN(n177), .Q(
        \mem[1][17] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][16]  ( .D(n272), .CP(clk), .RN(n177), .Q(
        \mem[1][16] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][15]  ( .D(n273), .CP(clk), .RN(n177), .Q(
        \mem[1][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][14]  ( .D(n274), .CP(clk), .RN(n177), .Q(
        \mem[1][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][13]  ( .D(n275), .CP(clk), .RN(n177), .Q(
        \mem[1][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][12]  ( .D(n276), .CP(clk), .RN(n177), .Q(
        \mem[1][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][11]  ( .D(n277), .CP(clk), .RN(n177), .Q(
        \mem[1][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][10]  ( .D(n278), .CP(clk), .RN(n177), .Q(
        \mem[1][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][9]  ( .D(n279), .CP(clk), .RN(n177), .Q(
        \mem[1][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][8]  ( .D(n280), .CP(clk), .RN(n177), .Q(
        \mem[1][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][7]  ( .D(n281), .CP(clk), .RN(n177), .Q(
        \mem[1][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][6]  ( .D(n282), .CP(clk), .RN(n177), .Q(
        \mem[1][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][5]  ( .D(n283), .CP(clk), .RN(n177), .Q(
        \mem[1][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][4]  ( .D(n284), .CP(clk), .RN(n178), .Q(
        \mem[1][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][3]  ( .D(n285), .CP(clk), .RN(n178), .Q(
        \mem[1][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][2]  ( .D(n286), .CP(clk), .RN(n178), .Q(
        \mem[1][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][1]  ( .D(n287), .CP(clk), .RN(n178), .Q(
        \mem[1][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][0]  ( .D(n288), .CP(clk), .RN(n178), .Q(
        \mem[1][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][31]  ( .D(n289), .CP(clk), .RN(n178), .Q(
        \mem[0][31] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][30]  ( .D(n290), .CP(clk), .RN(n178), .Q(
        \mem[0][30] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][29]  ( .D(n291), .CP(clk), .RN(n178), .Q(
        \mem[0][29] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][28]  ( .D(n292), .CP(clk), .RN(n178), .Q(
        \mem[0][28] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][27]  ( .D(n293), .CP(clk), .RN(n178), .Q(
        \mem[0][27] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][26]  ( .D(n294), .CP(clk), .RN(n178), .Q(
        \mem[0][26] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][25]  ( .D(n295), .CP(clk), .RN(n178), .Q(
        \mem[0][25] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][24]  ( .D(n296), .CP(clk), .RN(n178), .Q(
        \mem[0][24] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][23]  ( .D(n297), .CP(clk), .RN(n179), .Q(
        \mem[0][23] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][22]  ( .D(n298), .CP(clk), .RN(n179), .Q(
        \mem[0][22] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][21]  ( .D(n299), .CP(clk), .RN(n179), .Q(
        \mem[0][21] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][20]  ( .D(n300), .CP(clk), .RN(n179), .Q(
        \mem[0][20] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][19]  ( .D(n301), .CP(clk), .RN(n179), .Q(
        \mem[0][19] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][18]  ( .D(n302), .CP(clk), .RN(n179), .Q(
        \mem[0][18] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][17]  ( .D(n303), .CP(clk), .RN(n179), .Q(
        \mem[0][17] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][16]  ( .D(n304), .CP(clk), .RN(n179), .Q(
        \mem[0][16] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][15]  ( .D(n305), .CP(clk), .RN(n179), .Q(
        \mem[0][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][14]  ( .D(n306), .CP(clk), .RN(n179), .Q(
        \mem[0][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][13]  ( .D(n307), .CP(clk), .RN(n179), .Q(
        \mem[0][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][12]  ( .D(n308), .CP(clk), .RN(n179), .Q(
        \mem[0][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][11]  ( .D(n309), .CP(clk), .RN(n179), .Q(
        \mem[0][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][10]  ( .D(n310), .CP(clk), .RN(n180), .Q(
        \mem[0][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][9]  ( .D(n311), .CP(clk), .RN(n180), .Q(
        \mem[0][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][8]  ( .D(n312), .CP(clk), .RN(n180), .Q(
        \mem[0][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][7]  ( .D(n313), .CP(clk), .RN(n180), .Q(
        \mem[0][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][6]  ( .D(n314), .CP(clk), .RN(n180), .Q(
        \mem[0][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][5]  ( .D(n315), .CP(clk), .RN(n180), .Q(
        \mem[0][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][4]  ( .D(n316), .CP(clk), .RN(n180), .Q(
        \mem[0][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][3]  ( .D(n317), .CP(clk), .RN(n180), .Q(
        \mem[0][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][2]  ( .D(n318), .CP(clk), .RN(n180), .Q(
        \mem[0][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][1]  ( .D(n319), .CP(clk), .RN(n180), .Q(
        \mem[0][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][0]  ( .D(n320), .CP(clk), .RN(n180), .Q(
        \mem[0][0] ) );
  HS65_LS_DFPRQX9 \rd_data_reg[31]  ( .D(N17), .CP(clk), .RN(n180), .Q(
        rd_data[31]) );
  HS65_LS_DFPRQX9 \rd_data_reg[30]  ( .D(N18), .CP(clk), .RN(n180), .Q(
        rd_data[30]) );
  HS65_LS_DFPRQX9 \rd_data_reg[29]  ( .D(N19), .CP(clk), .RN(n181), .Q(
        rd_data[29]) );
  HS65_LS_DFPRQX9 \rd_data_reg[28]  ( .D(N20), .CP(clk), .RN(n181), .Q(
        rd_data[28]) );
  HS65_LS_DFPRQX9 \rd_data_reg[27]  ( .D(N21), .CP(clk), .RN(n181), .Q(
        rd_data[27]) );
  HS65_LS_DFPRQX9 \rd_data_reg[26]  ( .D(N22), .CP(clk), .RN(n181), .Q(
        rd_data[26]) );
  HS65_LS_DFPRQX9 \rd_data_reg[25]  ( .D(N23), .CP(clk), .RN(n181), .Q(
        rd_data[25]) );
  HS65_LS_DFPRQX9 \rd_data_reg[24]  ( .D(N24), .CP(clk), .RN(n181), .Q(
        rd_data[24]) );
  HS65_LS_DFPRQX9 \rd_data_reg[23]  ( .D(N25), .CP(clk), .RN(n181), .Q(
        rd_data[23]) );
  HS65_LS_DFPRQX9 \rd_data_reg[22]  ( .D(N26), .CP(clk), .RN(n181), .Q(
        rd_data[22]) );
  HS65_LS_DFPRQX9 \rd_data_reg[21]  ( .D(N27), .CP(clk), .RN(n181), .Q(
        rd_data[21]) );
  HS65_LS_DFPRQX9 \rd_data_reg[20]  ( .D(N28), .CP(clk), .RN(n181), .Q(
        rd_data[20]) );
  HS65_LS_DFPRQX9 \rd_data_reg[19]  ( .D(N29), .CP(clk), .RN(n181), .Q(
        rd_data[19]) );
  HS65_LS_DFPRQX9 \rd_data_reg[18]  ( .D(N30), .CP(clk), .RN(n181), .Q(
        rd_data[18]) );
  HS65_LS_DFPRQX9 \rd_data_reg[17]  ( .D(N31), .CP(clk), .RN(n181), .Q(
        rd_data[17]) );
  HS65_LS_DFPRQX9 \rd_data_reg[16]  ( .D(N32), .CP(clk), .RN(n182), .Q(
        rd_data[16]) );
  HS65_LS_DFPRQX9 \rd_data_reg[15]  ( .D(N33), .CP(clk), .RN(n182), .Q(
        rd_data[15]) );
  HS65_LS_DFPRQX9 \rd_data_reg[14]  ( .D(N34), .CP(clk), .RN(n182), .Q(
        rd_data[14]) );
  HS65_LS_DFPRQX9 \rd_data_reg[13]  ( .D(N35), .CP(clk), .RN(n182), .Q(
        rd_data[13]) );
  HS65_LS_DFPRQX9 \rd_data_reg[12]  ( .D(N36), .CP(clk), .RN(n182), .Q(
        rd_data[12]) );
  HS65_LS_DFPRQX9 \rd_data_reg[11]  ( .D(N37), .CP(clk), .RN(n182), .Q(
        rd_data[11]) );
  HS65_LS_DFPRQX9 \rd_data_reg[10]  ( .D(N38), .CP(clk), .RN(n182), .Q(
        rd_data[10]) );
  HS65_LS_DFPRQX9 \rd_data_reg[9]  ( .D(N39), .CP(clk), .RN(n182), .Q(
        rd_data[9]) );
  HS65_LS_DFPRQX9 \rd_data_reg[8]  ( .D(N40), .CP(clk), .RN(n182), .Q(
        rd_data[8]) );
  HS65_LS_DFPRQX9 \rd_data_reg[7]  ( .D(N41), .CP(clk), .RN(n182), .Q(
        rd_data[7]) );
  HS65_LS_DFPRQX9 \rd_data_reg[6]  ( .D(N42), .CP(clk), .RN(n182), .Q(
        rd_data[6]) );
  HS65_LS_DFPRQX9 \rd_data_reg[5]  ( .D(N43), .CP(clk), .RN(n182), .Q(
        rd_data[5]) );
  HS65_LS_DFPRQX9 \rd_data_reg[4]  ( .D(N44), .CP(clk), .RN(n182), .Q(
        rd_data[4]) );
  HS65_LS_DFPRQX9 \rd_data_reg[3]  ( .D(N45), .CP(clk), .RN(n183), .Q(
        rd_data[3]) );
  HS65_LS_DFPRQX9 \rd_data_reg[2]  ( .D(N46), .CP(clk), .RN(n183), .Q(
        rd_data[2]) );
  HS65_LS_DFPRQX9 \rd_data_reg[1]  ( .D(N47), .CP(clk), .RN(n183), .Q(
        rd_data[1]) );
  HS65_LS_DFPRQX9 \rd_data_reg[0]  ( .D(N48), .CP(clk), .RN(n183), .Q(
        rd_data[0]) );
  HS65_LS_AND3X9 U3 ( .A(n191), .B(n190), .C(wr_ena), .Z(n1) );
  HS65_LS_BFX9 U4 ( .A(n165), .Z(n162) );
  HS65_LS_BFX9 U5 ( .A(n1), .Z(n168) );
  HS65_LS_BFX9 U6 ( .A(n155), .Z(n152) );
  HS65_LS_BFX9 U7 ( .A(n160), .Z(n157) );
  HS65_LS_AND2X4 U8 ( .A(rd_addr[1]), .B(rd_addr[0]), .Z(n321) );
  HS65_LS_AND2X4 U9 ( .A(rd_addr[1]), .B(n192), .Z(n322) );
  HS65_LS_BFX9 U10 ( .A(n185), .Z(n180) );
  HS65_LS_BFX9 U11 ( .A(n185), .Z(n179) );
  HS65_LS_BFX9 U12 ( .A(n185), .Z(n178) );
  HS65_LS_BFX9 U13 ( .A(n186), .Z(n177) );
  HS65_LS_BFX9 U14 ( .A(n186), .Z(n176) );
  HS65_LS_BFX9 U15 ( .A(n186), .Z(n175) );
  HS65_LS_BFX9 U16 ( .A(n187), .Z(n174) );
  HS65_LS_BFX9 U17 ( .A(n187), .Z(n173) );
  HS65_LS_BFX9 U18 ( .A(n187), .Z(n172) );
  HS65_LS_BFX9 U19 ( .A(n188), .Z(n185) );
  HS65_LS_BFX9 U20 ( .A(n188), .Z(n186) );
  HS65_LS_BFX9 U21 ( .A(n189), .Z(n187) );
  HS65_LS_BFX9 U22 ( .A(n184), .Z(n182) );
  HS65_LS_BFX9 U23 ( .A(n184), .Z(n181) );
  HS65_LS_BFX9 U24 ( .A(n188), .Z(n171) );
  HS65_LS_BFX9 U25 ( .A(n189), .Z(n188) );
  HS65_LS_BFX9 U26 ( .A(n184), .Z(n183) );
  HS65_LS_BFX9 U27 ( .A(n189), .Z(n184) );
  HS65_LS_IVX9 U28 ( .A(reset), .Z(n189) );
  HS65_LS_IVX9 U29 ( .A(n168), .Z(n167) );
  HS65_LS_IVX9 U30 ( .A(n168), .Z(n166) );
  HS65_LS_IVX9 U31 ( .A(n162), .Z(n161) );
  HS65_LS_BFX9 U32 ( .A(n1), .Z(n169) );
  HS65_LS_BFX9 U33 ( .A(n165), .Z(n163) );
  HS65_LS_BFX9 U34 ( .A(n1), .Z(n170) );
  HS65_LS_BFX9 U35 ( .A(n162), .Z(n164) );
  HS65_LS_IVX9 U36 ( .A(n157), .Z(n156) );
  HS65_LS_IVX9 U37 ( .A(n152), .Z(n151) );
  HS65_LS_BFX9 U38 ( .A(n160), .Z(n158) );
  HS65_LS_BFX9 U39 ( .A(n155), .Z(n153) );
  HS65_LS_BFX9 U40 ( .A(n157), .Z(n159) );
  HS65_LS_BFX9 U41 ( .A(n152), .Z(n154) );
  HS65_LS_IVX9 U42 ( .A(n327), .Z(n165) );
  HS65_LS_IVX9 U43 ( .A(wr_addr[0]), .Z(n191) );
  HS65_LS_NAND3X5 U44 ( .A(wr_ena), .B(n190), .C(wr_addr[0]), .Z(n327) );
  HS65_LS_BFX9 U45 ( .A(n322), .Z(n6) );
  HS65_LS_BFX9 U46 ( .A(n322), .Z(n5) );
  HS65_LS_BFX9 U47 ( .A(n321), .Z(n3) );
  HS65_LS_BFX9 U48 ( .A(n321), .Z(n2) );
  HS65_LS_BFX9 U49 ( .A(n8), .Z(n145) );
  HS65_LS_BFX9 U50 ( .A(n8), .Z(n9) );
  HS65_LS_BFX9 U51 ( .A(n147), .Z(n149) );
  HS65_LS_BFX9 U52 ( .A(n147), .Z(n148) );
  HS65_LS_BFX9 U53 ( .A(n321), .Z(n4) );
  HS65_LS_BFX9 U54 ( .A(n322), .Z(n7) );
  HS65_LS_BFX9 U55 ( .A(n8), .Z(n146) );
  HS65_LS_BFX9 U56 ( .A(n147), .Z(n150) );
  HS65_LS_IVX9 U57 ( .A(n326), .Z(n160) );
  HS65_LS_IVX9 U58 ( .A(n325), .Z(n155) );
  HS65_LS_BFX9 U59 ( .A(n324), .Z(n147) );
  HS65_LS_NOR2X6 U60 ( .A(rd_addr[0]), .B(rd_addr[1]), .Z(n324) );
  HS65_LS_BFX9 U61 ( .A(n323), .Z(n8) );
  HS65_LS_NOR2X6 U62 ( .A(n192), .B(rd_addr[1]), .Z(n323) );
  HS65_LS_IVX9 U63 ( .A(wr_addr[1]), .Z(n190) );
  HS65_LS_NAND3X5 U64 ( .A(wr_addr[0]), .B(wr_ena), .C(wr_addr[1]), .Z(n325)
         );
  HS65_LS_NAND3X5 U65 ( .A(wr_ena), .B(n191), .C(wr_addr[1]), .Z(n326) );
  HS65_LS_IVX9 U66 ( .A(rd_addr[0]), .Z(n192) );
  HS65_LS_MX41X7 U67 ( .D0(n150), .S0(\mem[0][0] ), .D1(n146), .S1(\mem[1][0] ), .D2(n7), .S2(\mem[2][0] ), .D3(n4), .S3(\mem[3][0] ), .Z(N48) );
  HS65_LS_MX41X7 U68 ( .D0(n150), .S0(\mem[0][1] ), .D1(n146), .S1(\mem[1][1] ), .D2(n7), .S2(\mem[2][1] ), .D3(n4), .S3(\mem[3][1] ), .Z(N47) );
  HS65_LS_MX41X7 U69 ( .D0(n150), .S0(\mem[0][2] ), .D1(n146), .S1(\mem[1][2] ), .D2(n7), .S2(\mem[2][2] ), .D3(n4), .S3(\mem[3][2] ), .Z(N46) );
  HS65_LS_MX41X7 U70 ( .D0(n150), .S0(\mem[0][3] ), .D1(n146), .S1(\mem[1][3] ), .D2(n7), .S2(\mem[2][3] ), .D3(n4), .S3(\mem[3][3] ), .Z(N45) );
  HS65_LS_MX41X7 U71 ( .D0(n150), .S0(\mem[0][4] ), .D1(n146), .S1(\mem[1][4] ), .D2(n7), .S2(\mem[2][4] ), .D3(n4), .S3(\mem[3][4] ), .Z(N44) );
  HS65_LS_MX41X7 U72 ( .D0(n150), .S0(\mem[0][5] ), .D1(n146), .S1(\mem[1][5] ), .D2(n7), .S2(\mem[2][5] ), .D3(n4), .S3(\mem[3][5] ), .Z(N43) );
  HS65_LS_MX41X7 U73 ( .D0(n150), .S0(\mem[0][6] ), .D1(n146), .S1(\mem[1][6] ), .D2(n6), .S2(\mem[2][6] ), .D3(n4), .S3(\mem[3][6] ), .Z(N42) );
  HS65_LS_MX41X7 U74 ( .D0(n150), .S0(\mem[0][7] ), .D1(n146), .S1(\mem[1][7] ), .D2(n6), .S2(\mem[2][7] ), .D3(n4), .S3(\mem[3][7] ), .Z(N41) );
  HS65_LS_MX41X7 U75 ( .D0(n149), .S0(\mem[0][8] ), .D1(n145), .S1(\mem[1][8] ), .D2(n6), .S2(\mem[2][8] ), .D3(n3), .S3(\mem[3][8] ), .Z(N40) );
  HS65_LS_MX41X7 U76 ( .D0(n149), .S0(\mem[0][9] ), .D1(n145), .S1(\mem[1][9] ), .D2(n6), .S2(\mem[2][9] ), .D3(n3), .S3(\mem[3][9] ), .Z(N39) );
  HS65_LS_MX41X7 U77 ( .D0(n149), .S0(\mem[0][10] ), .D1(n145), .S1(
        \mem[1][10] ), .D2(n6), .S2(\mem[2][10] ), .D3(n3), .S3(\mem[3][10] ), 
        .Z(N38) );
  HS65_LS_MX41X7 U78 ( .D0(n149), .S0(\mem[0][11] ), .D1(n145), .S1(
        \mem[1][11] ), .D2(n6), .S2(\mem[2][11] ), .D3(n3), .S3(\mem[3][11] ), 
        .Z(N37) );
  HS65_LS_MX41X7 U79 ( .D0(n149), .S0(\mem[0][12] ), .D1(n145), .S1(
        \mem[1][12] ), .D2(n6), .S2(\mem[2][12] ), .D3(n3), .S3(\mem[3][12] ), 
        .Z(N36) );
  HS65_LS_MX41X7 U80 ( .D0(n149), .S0(\mem[0][13] ), .D1(n145), .S1(
        \mem[1][13] ), .D2(n6), .S2(\mem[2][13] ), .D3(n3), .S3(\mem[3][13] ), 
        .Z(N35) );
  HS65_LS_MX41X7 U81 ( .D0(n149), .S0(\mem[0][14] ), .D1(n145), .S1(
        \mem[1][14] ), .D2(n6), .S2(\mem[2][14] ), .D3(n3), .S3(\mem[3][14] ), 
        .Z(N34) );
  HS65_LS_MX41X7 U82 ( .D0(n149), .S0(\mem[0][15] ), .D1(n145), .S1(
        \mem[1][15] ), .D2(n6), .S2(\mem[2][15] ), .D3(n3), .S3(\mem[3][15] ), 
        .Z(N33) );
  HS65_LS_MX41X7 U83 ( .D0(n149), .S0(\mem[0][16] ), .D1(n145), .S1(
        \mem[1][16] ), .D2(n6), .S2(\mem[2][16] ), .D3(n3), .S3(\mem[3][16] ), 
        .Z(N32) );
  HS65_LS_MX41X7 U84 ( .D0(n149), .S0(\mem[0][17] ), .D1(n145), .S1(
        \mem[1][17] ), .D2(n6), .S2(\mem[2][17] ), .D3(n3), .S3(\mem[3][17] ), 
        .Z(N31) );
  HS65_LS_MX41X7 U85 ( .D0(n149), .S0(\mem[0][18] ), .D1(n145), .S1(
        \mem[1][18] ), .D2(n6), .S2(\mem[2][18] ), .D3(n3), .S3(\mem[3][18] ), 
        .Z(N30) );
  HS65_LS_MX41X7 U86 ( .D0(n149), .S0(\mem[0][19] ), .D1(n145), .S1(
        \mem[1][19] ), .D2(n5), .S2(\mem[2][19] ), .D3(n3), .S3(\mem[3][19] ), 
        .Z(N29) );
  HS65_LS_MX41X7 U87 ( .D0(n148), .S0(\mem[0][20] ), .D1(n9), .S1(\mem[1][20] ), .D2(n5), .S2(\mem[2][20] ), .D3(n2), .S3(\mem[3][20] ), .Z(N28) );
  HS65_LS_MX41X7 U88 ( .D0(n148), .S0(\mem[0][21] ), .D1(n9), .S1(\mem[1][21] ), .D2(n5), .S2(\mem[2][21] ), .D3(n2), .S3(\mem[3][21] ), .Z(N27) );
  HS65_LS_MX41X7 U89 ( .D0(n148), .S0(\mem[0][22] ), .D1(n9), .S1(\mem[1][22] ), .D2(n5), .S2(\mem[2][22] ), .D3(n2), .S3(\mem[3][22] ), .Z(N26) );
  HS65_LS_MX41X7 U90 ( .D0(n148), .S0(\mem[0][23] ), .D1(n9), .S1(\mem[1][23] ), .D2(n5), .S2(\mem[2][23] ), .D3(n2), .S3(\mem[3][23] ), .Z(N25) );
  HS65_LS_MX41X7 U91 ( .D0(n148), .S0(\mem[0][24] ), .D1(n9), .S1(\mem[1][24] ), .D2(n5), .S2(\mem[2][24] ), .D3(n2), .S3(\mem[3][24] ), .Z(N24) );
  HS65_LS_MX41X7 U92 ( .D0(n148), .S0(\mem[0][25] ), .D1(n9), .S1(\mem[1][25] ), .D2(n5), .S2(\mem[2][25] ), .D3(n2), .S3(\mem[3][25] ), .Z(N23) );
  HS65_LS_MX41X7 U93 ( .D0(n148), .S0(\mem[0][26] ), .D1(n9), .S1(\mem[1][26] ), .D2(n5), .S2(\mem[2][26] ), .D3(n2), .S3(\mem[3][26] ), .Z(N22) );
  HS65_LS_MX41X7 U94 ( .D0(n148), .S0(\mem[0][27] ), .D1(n9), .S1(\mem[1][27] ), .D2(n5), .S2(\mem[2][27] ), .D3(n2), .S3(\mem[3][27] ), .Z(N21) );
  HS65_LS_MX41X7 U95 ( .D0(n148), .S0(\mem[0][28] ), .D1(n9), .S1(\mem[1][28] ), .D2(n5), .S2(\mem[2][28] ), .D3(n2), .S3(\mem[3][28] ), .Z(N20) );
  HS65_LS_MX41X7 U96 ( .D0(n148), .S0(\mem[0][29] ), .D1(n9), .S1(\mem[1][29] ), .D2(n5), .S2(\mem[2][29] ), .D3(n2), .S3(\mem[3][29] ), .Z(N19) );
  HS65_LS_MX41X7 U97 ( .D0(n148), .S0(\mem[0][30] ), .D1(n9), .S1(\mem[1][30] ), .D2(n5), .S2(\mem[2][30] ), .D3(n2), .S3(\mem[3][30] ), .Z(N18) );
  HS65_LS_MX41X7 U98 ( .D0(n148), .S0(\mem[0][31] ), .D1(n9), .S1(\mem[1][31] ), .D2(n5), .S2(\mem[2][31] ), .D3(n2), .S3(\mem[3][31] ), .Z(N17) );
  HS65_LS_AO22X9 U99 ( .A(wr_data[0]), .B(n154), .C(n151), .D(\mem[3][0] ), 
        .Z(n224) );
  HS65_LS_AO22X9 U100 ( .A(wr_data[1]), .B(n154), .C(n151), .D(\mem[3][1] ), 
        .Z(n223) );
  HS65_LS_AO22X9 U101 ( .A(wr_data[2]), .B(n154), .C(n151), .D(\mem[3][2] ), 
        .Z(n222) );
  HS65_LS_AO22X9 U102 ( .A(wr_data[3]), .B(n154), .C(n151), .D(\mem[3][3] ), 
        .Z(n221) );
  HS65_LS_AO22X9 U103 ( .A(wr_data[4]), .B(n154), .C(n151), .D(\mem[3][4] ), 
        .Z(n220) );
  HS65_LS_AO22X9 U104 ( .A(wr_data[5]), .B(n154), .C(n151), .D(\mem[3][5] ), 
        .Z(n219) );
  HS65_LS_AO22X9 U105 ( .A(wr_data[6]), .B(n154), .C(n151), .D(\mem[3][6] ), 
        .Z(n218) );
  HS65_LS_AO22X9 U106 ( .A(wr_data[7]), .B(n154), .C(n151), .D(\mem[3][7] ), 
        .Z(n217) );
  HS65_LS_AO22X9 U107 ( .A(wr_data[8]), .B(n154), .C(n151), .D(\mem[3][8] ), 
        .Z(n216) );
  HS65_LS_AO22X9 U108 ( .A(wr_data[9]), .B(n154), .C(n151), .D(\mem[3][9] ), 
        .Z(n215) );
  HS65_LS_AO22X9 U109 ( .A(wr_data[10]), .B(n154), .C(n151), .D(\mem[3][10] ), 
        .Z(n214) );
  HS65_LS_AO22X9 U110 ( .A(wr_data[11]), .B(n153), .C(n151), .D(\mem[3][11] ), 
        .Z(n213) );
  HS65_LS_AO22X9 U111 ( .A(wr_data[12]), .B(n153), .C(n151), .D(\mem[3][12] ), 
        .Z(n212) );
  HS65_LS_AO22X9 U112 ( .A(wr_data[13]), .B(n153), .C(n151), .D(\mem[3][13] ), 
        .Z(n211) );
  HS65_LS_AO22X9 U113 ( .A(wr_data[14]), .B(n153), .C(n151), .D(\mem[3][14] ), 
        .Z(n210) );
  HS65_LS_AO22X9 U114 ( .A(wr_data[15]), .B(n153), .C(n151), .D(\mem[3][15] ), 
        .Z(n209) );
  HS65_LS_AO22X9 U115 ( .A(wr_data[16]), .B(n153), .C(n151), .D(\mem[3][16] ), 
        .Z(n208) );
  HS65_LS_AO22X9 U116 ( .A(wr_data[17]), .B(n153), .C(n151), .D(\mem[3][17] ), 
        .Z(n207) );
  HS65_LS_AO22X9 U117 ( .A(wr_data[18]), .B(n153), .C(n151), .D(\mem[3][18] ), 
        .Z(n206) );
  HS65_LS_AO22X9 U118 ( .A(wr_data[19]), .B(n153), .C(n151), .D(\mem[3][19] ), 
        .Z(n205) );
  HS65_LS_AO22X9 U119 ( .A(wr_data[20]), .B(n153), .C(n325), .D(\mem[3][20] ), 
        .Z(n204) );
  HS65_LS_AO22X9 U120 ( .A(wr_data[21]), .B(n153), .C(n325), .D(\mem[3][21] ), 
        .Z(n203) );
  HS65_LS_AO22X9 U121 ( .A(wr_data[22]), .B(n153), .C(n325), .D(\mem[3][22] ), 
        .Z(n202) );
  HS65_LS_AO22X9 U122 ( .A(wr_data[23]), .B(n153), .C(n325), .D(\mem[3][23] ), 
        .Z(n201) );
  HS65_LS_AO22X9 U123 ( .A(wr_data[24]), .B(n153), .C(n325), .D(\mem[3][24] ), 
        .Z(n200) );
  HS65_LS_AO22X9 U124 ( .A(wr_data[25]), .B(n153), .C(n325), .D(\mem[3][25] ), 
        .Z(n199) );
  HS65_LS_AO22X9 U125 ( .A(wr_data[26]), .B(n153), .C(n325), .D(\mem[3][26] ), 
        .Z(n198) );
  HS65_LS_AO22X9 U126 ( .A(wr_data[27]), .B(n153), .C(n325), .D(\mem[3][27] ), 
        .Z(n197) );
  HS65_LS_AO22X9 U127 ( .A(wr_data[28]), .B(n153), .C(n325), .D(\mem[3][28] ), 
        .Z(n196) );
  HS65_LS_AO22X9 U128 ( .A(wr_data[29]), .B(n153), .C(n325), .D(\mem[3][29] ), 
        .Z(n195) );
  HS65_LS_AO22X9 U129 ( .A(wr_data[30]), .B(n153), .C(n325), .D(\mem[3][30] ), 
        .Z(n194) );
  HS65_LS_AO22X9 U130 ( .A(wr_data[31]), .B(n152), .C(n325), .D(\mem[3][31] ), 
        .Z(n193) );
  HS65_LS_AO22X9 U131 ( .A(wr_data[0]), .B(n164), .C(n161), .D(\mem[1][0] ), 
        .Z(n288) );
  HS65_LS_AO22X9 U132 ( .A(wr_data[1]), .B(n164), .C(n161), .D(\mem[1][1] ), 
        .Z(n287) );
  HS65_LS_AO22X9 U133 ( .A(wr_data[2]), .B(n164), .C(n161), .D(\mem[1][2] ), 
        .Z(n286) );
  HS65_LS_AO22X9 U134 ( .A(wr_data[3]), .B(n164), .C(n161), .D(\mem[1][3] ), 
        .Z(n285) );
  HS65_LS_AO22X9 U135 ( .A(wr_data[4]), .B(n164), .C(n161), .D(\mem[1][4] ), 
        .Z(n284) );
  HS65_LS_AO22X9 U136 ( .A(wr_data[5]), .B(n164), .C(n161), .D(\mem[1][5] ), 
        .Z(n283) );
  HS65_LS_AO22X9 U137 ( .A(wr_data[6]), .B(n164), .C(n161), .D(\mem[1][6] ), 
        .Z(n282) );
  HS65_LS_AO22X9 U138 ( .A(wr_data[7]), .B(n164), .C(n161), .D(\mem[1][7] ), 
        .Z(n281) );
  HS65_LS_AO22X9 U139 ( .A(wr_data[8]), .B(n164), .C(n161), .D(\mem[1][8] ), 
        .Z(n280) );
  HS65_LS_AO22X9 U140 ( .A(wr_data[9]), .B(n164), .C(n161), .D(\mem[1][9] ), 
        .Z(n279) );
  HS65_LS_AO22X9 U141 ( .A(wr_data[10]), .B(n164), .C(n161), .D(\mem[1][10] ), 
        .Z(n278) );
  HS65_LS_AO22X9 U142 ( .A(wr_data[11]), .B(n163), .C(n161), .D(\mem[1][11] ), 
        .Z(n277) );
  HS65_LS_AO22X9 U143 ( .A(wr_data[12]), .B(n163), .C(n161), .D(\mem[1][12] ), 
        .Z(n276) );
  HS65_LS_AO22X9 U144 ( .A(wr_data[13]), .B(n163), .C(n161), .D(\mem[1][13] ), 
        .Z(n275) );
  HS65_LS_AO22X9 U145 ( .A(wr_data[14]), .B(n163), .C(n161), .D(\mem[1][14] ), 
        .Z(n274) );
  HS65_LS_AO22X9 U146 ( .A(wr_data[15]), .B(n163), .C(n161), .D(\mem[1][15] ), 
        .Z(n273) );
  HS65_LS_AO22X9 U147 ( .A(wr_data[16]), .B(n163), .C(n161), .D(\mem[1][16] ), 
        .Z(n272) );
  HS65_LS_AO22X9 U148 ( .A(wr_data[17]), .B(n163), .C(n161), .D(\mem[1][17] ), 
        .Z(n271) );
  HS65_LS_AO22X9 U149 ( .A(wr_data[18]), .B(n163), .C(n161), .D(\mem[1][18] ), 
        .Z(n270) );
  HS65_LS_AO22X9 U150 ( .A(wr_data[19]), .B(n163), .C(n161), .D(\mem[1][19] ), 
        .Z(n269) );
  HS65_LS_AO22X9 U151 ( .A(wr_data[20]), .B(n163), .C(n327), .D(\mem[1][20] ), 
        .Z(n268) );
  HS65_LS_AO22X9 U152 ( .A(wr_data[21]), .B(n163), .C(n327), .D(\mem[1][21] ), 
        .Z(n267) );
  HS65_LS_AO22X9 U153 ( .A(wr_data[22]), .B(n163), .C(n327), .D(\mem[1][22] ), 
        .Z(n266) );
  HS65_LS_AO22X9 U154 ( .A(wr_data[23]), .B(n163), .C(n327), .D(\mem[1][23] ), 
        .Z(n265) );
  HS65_LS_AO22X9 U155 ( .A(wr_data[24]), .B(n163), .C(n327), .D(\mem[1][24] ), 
        .Z(n264) );
  HS65_LS_AO22X9 U156 ( .A(wr_data[25]), .B(n163), .C(n327), .D(\mem[1][25] ), 
        .Z(n263) );
  HS65_LS_AO22X9 U157 ( .A(wr_data[26]), .B(n163), .C(n327), .D(\mem[1][26] ), 
        .Z(n262) );
  HS65_LS_AO22X9 U158 ( .A(wr_data[27]), .B(n163), .C(n327), .D(\mem[1][27] ), 
        .Z(n261) );
  HS65_LS_AO22X9 U159 ( .A(wr_data[28]), .B(n163), .C(n327), .D(\mem[1][28] ), 
        .Z(n260) );
  HS65_LS_AO22X9 U160 ( .A(wr_data[29]), .B(n163), .C(n327), .D(\mem[1][29] ), 
        .Z(n259) );
  HS65_LS_AO22X9 U161 ( .A(wr_data[30]), .B(n163), .C(n327), .D(\mem[1][30] ), 
        .Z(n258) );
  HS65_LS_AO22X9 U162 ( .A(wr_data[31]), .B(n162), .C(n327), .D(\mem[1][31] ), 
        .Z(n257) );
  HS65_LS_AO22X9 U163 ( .A(n170), .B(wr_data[0]), .C(n167), .D(\mem[0][0] ), 
        .Z(n320) );
  HS65_LS_AO22X9 U164 ( .A(n170), .B(wr_data[1]), .C(n166), .D(\mem[0][1] ), 
        .Z(n319) );
  HS65_LS_AO22X9 U165 ( .A(n170), .B(wr_data[2]), .C(n167), .D(\mem[0][2] ), 
        .Z(n318) );
  HS65_LS_AO22X9 U166 ( .A(n170), .B(wr_data[3]), .C(n166), .D(\mem[0][3] ), 
        .Z(n317) );
  HS65_LS_AO22X9 U167 ( .A(n170), .B(wr_data[4]), .C(n167), .D(\mem[0][4] ), 
        .Z(n316) );
  HS65_LS_AO22X9 U168 ( .A(n170), .B(wr_data[5]), .C(n166), .D(\mem[0][5] ), 
        .Z(n315) );
  HS65_LS_AO22X9 U169 ( .A(n170), .B(wr_data[6]), .C(n167), .D(\mem[0][6] ), 
        .Z(n314) );
  HS65_LS_AO22X9 U170 ( .A(n170), .B(wr_data[7]), .C(n167), .D(\mem[0][7] ), 
        .Z(n313) );
  HS65_LS_AO22X9 U171 ( .A(n170), .B(wr_data[8]), .C(n167), .D(\mem[0][8] ), 
        .Z(n312) );
  HS65_LS_AO22X9 U172 ( .A(n170), .B(wr_data[9]), .C(n167), .D(\mem[0][9] ), 
        .Z(n311) );
  HS65_LS_AO22X9 U173 ( .A(n170), .B(wr_data[10]), .C(n167), .D(\mem[0][10] ), 
        .Z(n310) );
  HS65_LS_AO22X9 U174 ( .A(n169), .B(wr_data[11]), .C(n167), .D(\mem[0][11] ), 
        .Z(n309) );
  HS65_LS_AO22X9 U175 ( .A(n169), .B(wr_data[12]), .C(n167), .D(\mem[0][12] ), 
        .Z(n308) );
  HS65_LS_AO22X9 U176 ( .A(n169), .B(wr_data[13]), .C(n167), .D(\mem[0][13] ), 
        .Z(n307) );
  HS65_LS_AO22X9 U177 ( .A(n169), .B(wr_data[14]), .C(n167), .D(\mem[0][14] ), 
        .Z(n306) );
  HS65_LS_AO22X9 U178 ( .A(n169), .B(wr_data[15]), .C(n167), .D(\mem[0][15] ), 
        .Z(n305) );
  HS65_LS_AO22X9 U179 ( .A(n169), .B(wr_data[16]), .C(n167), .D(\mem[0][16] ), 
        .Z(n304) );
  HS65_LS_AO22X9 U180 ( .A(n169), .B(wr_data[17]), .C(n167), .D(\mem[0][17] ), 
        .Z(n303) );
  HS65_LS_AO22X9 U181 ( .A(n169), .B(wr_data[18]), .C(n167), .D(\mem[0][18] ), 
        .Z(n302) );
  HS65_LS_AO22X9 U182 ( .A(n169), .B(wr_data[19]), .C(n166), .D(\mem[0][19] ), 
        .Z(n301) );
  HS65_LS_AO22X9 U183 ( .A(n169), .B(wr_data[20]), .C(n166), .D(\mem[0][20] ), 
        .Z(n300) );
  HS65_LS_AO22X9 U184 ( .A(n169), .B(wr_data[21]), .C(n166), .D(\mem[0][21] ), 
        .Z(n299) );
  HS65_LS_AO22X9 U185 ( .A(n169), .B(wr_data[22]), .C(n166), .D(\mem[0][22] ), 
        .Z(n298) );
  HS65_LS_AO22X9 U186 ( .A(n169), .B(wr_data[23]), .C(n166), .D(\mem[0][23] ), 
        .Z(n297) );
  HS65_LS_AO22X9 U187 ( .A(n169), .B(wr_data[24]), .C(n166), .D(\mem[0][24] ), 
        .Z(n296) );
  HS65_LS_AO22X9 U188 ( .A(n169), .B(wr_data[25]), .C(n166), .D(\mem[0][25] ), 
        .Z(n295) );
  HS65_LS_AO22X9 U189 ( .A(n169), .B(wr_data[26]), .C(n166), .D(\mem[0][26] ), 
        .Z(n294) );
  HS65_LS_AO22X9 U190 ( .A(n169), .B(wr_data[27]), .C(n166), .D(\mem[0][27] ), 
        .Z(n293) );
  HS65_LS_AO22X9 U191 ( .A(n169), .B(wr_data[28]), .C(n166), .D(\mem[0][28] ), 
        .Z(n292) );
  HS65_LS_AO22X9 U192 ( .A(n169), .B(wr_data[29]), .C(n166), .D(\mem[0][29] ), 
        .Z(n291) );
  HS65_LS_AO22X9 U193 ( .A(n169), .B(wr_data[30]), .C(n166), .D(\mem[0][30] ), 
        .Z(n290) );
  HS65_LS_AO22X9 U194 ( .A(n168), .B(wr_data[31]), .C(n166), .D(\mem[0][31] ), 
        .Z(n289) );
  HS65_LS_AO22X9 U195 ( .A(wr_data[0]), .B(n159), .C(n156), .D(\mem[2][0] ), 
        .Z(n256) );
  HS65_LS_AO22X9 U196 ( .A(wr_data[1]), .B(n159), .C(n156), .D(\mem[2][1] ), 
        .Z(n255) );
  HS65_LS_AO22X9 U197 ( .A(wr_data[2]), .B(n159), .C(n156), .D(\mem[2][2] ), 
        .Z(n254) );
  HS65_LS_AO22X9 U198 ( .A(wr_data[3]), .B(n159), .C(n156), .D(\mem[2][3] ), 
        .Z(n253) );
  HS65_LS_AO22X9 U199 ( .A(wr_data[4]), .B(n159), .C(n156), .D(\mem[2][4] ), 
        .Z(n252) );
  HS65_LS_AO22X9 U200 ( .A(wr_data[5]), .B(n159), .C(n156), .D(\mem[2][5] ), 
        .Z(n251) );
  HS65_LS_AO22X9 U201 ( .A(wr_data[6]), .B(n159), .C(n156), .D(\mem[2][6] ), 
        .Z(n250) );
  HS65_LS_AO22X9 U202 ( .A(wr_data[7]), .B(n159), .C(n156), .D(\mem[2][7] ), 
        .Z(n249) );
  HS65_LS_AO22X9 U203 ( .A(wr_data[8]), .B(n159), .C(n156), .D(\mem[2][8] ), 
        .Z(n248) );
  HS65_LS_AO22X9 U204 ( .A(wr_data[9]), .B(n159), .C(n156), .D(\mem[2][9] ), 
        .Z(n247) );
  HS65_LS_AO22X9 U205 ( .A(wr_data[10]), .B(n159), .C(n156), .D(\mem[2][10] ), 
        .Z(n246) );
  HS65_LS_AO22X9 U206 ( .A(wr_data[11]), .B(n158), .C(n156), .D(\mem[2][11] ), 
        .Z(n245) );
  HS65_LS_AO22X9 U207 ( .A(wr_data[12]), .B(n158), .C(n156), .D(\mem[2][12] ), 
        .Z(n244) );
  HS65_LS_AO22X9 U208 ( .A(wr_data[13]), .B(n158), .C(n156), .D(\mem[2][13] ), 
        .Z(n243) );
  HS65_LS_AO22X9 U209 ( .A(wr_data[14]), .B(n158), .C(n156), .D(\mem[2][14] ), 
        .Z(n242) );
  HS65_LS_AO22X9 U210 ( .A(wr_data[15]), .B(n158), .C(n156), .D(\mem[2][15] ), 
        .Z(n241) );
  HS65_LS_AO22X9 U211 ( .A(wr_data[16]), .B(n158), .C(n156), .D(\mem[2][16] ), 
        .Z(n240) );
  HS65_LS_AO22X9 U212 ( .A(wr_data[17]), .B(n158), .C(n156), .D(\mem[2][17] ), 
        .Z(n239) );
  HS65_LS_AO22X9 U213 ( .A(wr_data[18]), .B(n158), .C(n156), .D(\mem[2][18] ), 
        .Z(n238) );
  HS65_LS_AO22X9 U214 ( .A(wr_data[19]), .B(n158), .C(n156), .D(\mem[2][19] ), 
        .Z(n237) );
  HS65_LS_AO22X9 U215 ( .A(wr_data[20]), .B(n158), .C(n326), .D(\mem[2][20] ), 
        .Z(n236) );
  HS65_LS_AO22X9 U216 ( .A(wr_data[21]), .B(n158), .C(n326), .D(\mem[2][21] ), 
        .Z(n235) );
  HS65_LS_AO22X9 U217 ( .A(wr_data[22]), .B(n158), .C(n326), .D(\mem[2][22] ), 
        .Z(n234) );
  HS65_LS_AO22X9 U218 ( .A(wr_data[23]), .B(n158), .C(n326), .D(\mem[2][23] ), 
        .Z(n233) );
  HS65_LS_AO22X9 U219 ( .A(wr_data[24]), .B(n158), .C(n326), .D(\mem[2][24] ), 
        .Z(n232) );
  HS65_LS_AO22X9 U220 ( .A(wr_data[25]), .B(n158), .C(n326), .D(\mem[2][25] ), 
        .Z(n231) );
  HS65_LS_AO22X9 U221 ( .A(wr_data[26]), .B(n158), .C(n326), .D(\mem[2][26] ), 
        .Z(n230) );
  HS65_LS_AO22X9 U222 ( .A(wr_data[27]), .B(n158), .C(n326), .D(\mem[2][27] ), 
        .Z(n229) );
  HS65_LS_AO22X9 U223 ( .A(wr_data[28]), .B(n158), .C(n326), .D(\mem[2][28] ), 
        .Z(n228) );
  HS65_LS_AO22X9 U224 ( .A(wr_data[29]), .B(n158), .C(n326), .D(\mem[2][29] ), 
        .Z(n227) );
  HS65_LS_AO22X9 U225 ( .A(wr_data[30]), .B(n158), .C(n326), .D(\mem[2][30] ), 
        .Z(n226) );
  HS65_LS_AO22X9 U226 ( .A(wr_data[31]), .B(n157), .C(n326), .D(\mem[2][31] ), 
        .Z(n225) );
endmodule


module bram_DATA16_ADDR2_1 ( clk, reset, rd_addr, wr_addr, wr_data, wr_ena, 
        rd_data );
  input [1:0] rd_addr;
  input [1:0] wr_addr;
  input [15:0] wr_data;
  output [15:0] rd_data;
  input clk, reset, wr_ena;
  wire   \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] ,
         \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][15] , \mem[1][14] , \mem[1][13] ,
         \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] , \mem[1][8] ,
         \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] ,
         \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][15] , \mem[0][14] ,
         \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] ,
         \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] ,
         \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, n1,
         n2, n3, n4, n5, n6, n7, n8, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162;

  HS65_LS_DFPRQX9 \mem_reg[3][15]  ( .D(n91), .CP(clk), .RN(n1), .Q(
        \mem[3][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][14]  ( .D(n92), .CP(clk), .RN(n1), .Q(
        \mem[3][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][13]  ( .D(n93), .CP(clk), .RN(n1), .Q(
        \mem[3][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][12]  ( .D(n94), .CP(clk), .RN(n1), .Q(
        \mem[3][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][11]  ( .D(n95), .CP(clk), .RN(n1), .Q(
        \mem[3][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][10]  ( .D(n96), .CP(clk), .RN(n1), .Q(
        \mem[3][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][9]  ( .D(n97), .CP(clk), .RN(n1), .Q(\mem[3][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][8]  ( .D(n98), .CP(clk), .RN(n1), .Q(\mem[3][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][7]  ( .D(n99), .CP(clk), .RN(n1), .Q(\mem[3][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][6]  ( .D(n100), .CP(clk), .RN(n1), .Q(
        \mem[3][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][5]  ( .D(n101), .CP(clk), .RN(n1), .Q(
        \mem[3][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][4]  ( .D(n102), .CP(clk), .RN(n1), .Q(
        \mem[3][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][3]  ( .D(n103), .CP(clk), .RN(n1), .Q(
        \mem[3][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][2]  ( .D(n104), .CP(clk), .RN(n2), .Q(
        \mem[3][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][1]  ( .D(n105), .CP(clk), .RN(n2), .Q(
        \mem[3][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[3][0]  ( .D(n106), .CP(clk), .RN(n2), .Q(
        \mem[3][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][15]  ( .D(n107), .CP(clk), .RN(n2), .Q(
        \mem[2][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][14]  ( .D(n108), .CP(clk), .RN(n2), .Q(
        \mem[2][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][13]  ( .D(n109), .CP(clk), .RN(n2), .Q(
        \mem[2][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][12]  ( .D(n110), .CP(clk), .RN(n2), .Q(
        \mem[2][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][11]  ( .D(n111), .CP(clk), .RN(n2), .Q(
        \mem[2][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][10]  ( .D(n112), .CP(clk), .RN(n2), .Q(
        \mem[2][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][9]  ( .D(n113), .CP(clk), .RN(n2), .Q(
        \mem[2][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][8]  ( .D(n114), .CP(clk), .RN(n2), .Q(
        \mem[2][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][7]  ( .D(n115), .CP(clk), .RN(n2), .Q(
        \mem[2][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][6]  ( .D(n116), .CP(clk), .RN(n2), .Q(
        \mem[2][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][5]  ( .D(n117), .CP(clk), .RN(n3), .Q(
        \mem[2][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][4]  ( .D(n118), .CP(clk), .RN(n3), .Q(
        \mem[2][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][3]  ( .D(n119), .CP(clk), .RN(n3), .Q(
        \mem[2][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][2]  ( .D(n120), .CP(clk), .RN(n3), .Q(
        \mem[2][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][1]  ( .D(n121), .CP(clk), .RN(n3), .Q(
        \mem[2][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[2][0]  ( .D(n122), .CP(clk), .RN(n3), .Q(
        \mem[2][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][15]  ( .D(n123), .CP(clk), .RN(n3), .Q(
        \mem[1][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][14]  ( .D(n124), .CP(clk), .RN(n3), .Q(
        \mem[1][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][13]  ( .D(n125), .CP(clk), .RN(n3), .Q(
        \mem[1][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][12]  ( .D(n126), .CP(clk), .RN(n3), .Q(
        \mem[1][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][11]  ( .D(n127), .CP(clk), .RN(n3), .Q(
        \mem[1][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][10]  ( .D(n128), .CP(clk), .RN(n3), .Q(
        \mem[1][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][9]  ( .D(n129), .CP(clk), .RN(n3), .Q(
        \mem[1][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][8]  ( .D(n130), .CP(clk), .RN(n4), .Q(
        \mem[1][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][7]  ( .D(n131), .CP(clk), .RN(n4), .Q(
        \mem[1][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][6]  ( .D(n132), .CP(clk), .RN(n4), .Q(
        \mem[1][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][5]  ( .D(n133), .CP(clk), .RN(n4), .Q(
        \mem[1][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][4]  ( .D(n134), .CP(clk), .RN(n4), .Q(
        \mem[1][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][3]  ( .D(n135), .CP(clk), .RN(n4), .Q(
        \mem[1][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][2]  ( .D(n136), .CP(clk), .RN(n4), .Q(
        \mem[1][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][1]  ( .D(n137), .CP(clk), .RN(n4), .Q(
        \mem[1][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][0]  ( .D(n138), .CP(clk), .RN(n4), .Q(
        \mem[1][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][15]  ( .D(n139), .CP(clk), .RN(n4), .Q(
        \mem[0][15] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][14]  ( .D(n140), .CP(clk), .RN(n4), .Q(
        \mem[0][14] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][13]  ( .D(n141), .CP(clk), .RN(n4), .Q(
        \mem[0][13] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][12]  ( .D(n142), .CP(clk), .RN(n4), .Q(
        \mem[0][12] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][11]  ( .D(n143), .CP(clk), .RN(n5), .Q(
        \mem[0][11] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][10]  ( .D(n144), .CP(clk), .RN(n5), .Q(
        \mem[0][10] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][9]  ( .D(n145), .CP(clk), .RN(n5), .Q(
        \mem[0][9] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][8]  ( .D(n146), .CP(clk), .RN(n5), .Q(
        \mem[0][8] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][7]  ( .D(n147), .CP(clk), .RN(n5), .Q(
        \mem[0][7] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][6]  ( .D(n148), .CP(clk), .RN(n5), .Q(
        \mem[0][6] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][5]  ( .D(n149), .CP(clk), .RN(n5), .Q(
        \mem[0][5] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][4]  ( .D(n150), .CP(clk), .RN(n5), .Q(
        \mem[0][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][3]  ( .D(n151), .CP(clk), .RN(n5), .Q(
        \mem[0][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][2]  ( .D(n152), .CP(clk), .RN(n5), .Q(
        \mem[0][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][1]  ( .D(n153), .CP(clk), .RN(n5), .Q(
        \mem[0][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][0]  ( .D(n154), .CP(clk), .RN(n5), .Q(
        \mem[0][0] ) );
  HS65_LS_DFPRQX9 \rd_data_reg[15]  ( .D(N17), .CP(clk), .RN(n5), .Q(
        rd_data[15]) );
  HS65_LS_DFPRQX9 \rd_data_reg[14]  ( .D(N18), .CP(clk), .RN(n6), .Q(
        rd_data[14]) );
  HS65_LS_DFPRQX9 \rd_data_reg[13]  ( .D(N19), .CP(clk), .RN(n6), .Q(
        rd_data[13]) );
  HS65_LS_DFPRQX9 \rd_data_reg[12]  ( .D(N20), .CP(clk), .RN(n6), .Q(
        rd_data[12]) );
  HS65_LS_DFPRQX9 \rd_data_reg[11]  ( .D(N21), .CP(clk), .RN(n6), .Q(
        rd_data[11]) );
  HS65_LS_DFPRQX9 \rd_data_reg[10]  ( .D(N22), .CP(clk), .RN(n6), .Q(
        rd_data[10]) );
  HS65_LS_DFPRQX9 \rd_data_reg[9]  ( .D(N23), .CP(clk), .RN(n6), .Q(rd_data[9]) );
  HS65_LS_DFPRQX9 \rd_data_reg[8]  ( .D(N24), .CP(clk), .RN(n6), .Q(rd_data[8]) );
  HS65_LS_DFPRQX9 \rd_data_reg[7]  ( .D(N25), .CP(clk), .RN(n6), .Q(rd_data[7]) );
  HS65_LS_DFPRQX9 \rd_data_reg[6]  ( .D(N26), .CP(clk), .RN(n6), .Q(rd_data[6]) );
  HS65_LS_DFPRQX9 \rd_data_reg[5]  ( .D(N27), .CP(clk), .RN(n6), .Q(rd_data[5]) );
  HS65_LS_DFPRQX9 \rd_data_reg[4]  ( .D(N28), .CP(clk), .RN(n6), .Q(rd_data[4]) );
  HS65_LS_DFPRQX9 \rd_data_reg[3]  ( .D(N29), .CP(clk), .RN(n6), .Q(rd_data[3]) );
  HS65_LS_DFPRQX9 \rd_data_reg[2]  ( .D(N30), .CP(clk), .RN(n6), .Q(rd_data[2]) );
  HS65_LS_DFPRQX9 \rd_data_reg[1]  ( .D(N31), .CP(clk), .RN(n7), .Q(rd_data[1]) );
  HS65_LS_DFPRQX9 \rd_data_reg[0]  ( .D(N32), .CP(clk), .RN(n7), .Q(rd_data[0]) );
  HS65_LS_BFX9 U3 ( .A(n81), .Z(n4) );
  HS65_LS_BFX9 U4 ( .A(n81), .Z(n3) );
  HS65_LS_BFX9 U5 ( .A(n81), .Z(n2) );
  HS65_LS_BFX9 U6 ( .A(n83), .Z(n81) );
  HS65_LS_BFX9 U7 ( .A(n8), .Z(n6) );
  HS65_LS_BFX9 U8 ( .A(n8), .Z(n5) );
  HS65_LS_BFX9 U9 ( .A(n82), .Z(n1) );
  HS65_LS_BFX9 U10 ( .A(n83), .Z(n82) );
  HS65_LS_BFX9 U11 ( .A(n8), .Z(n7) );
  HS65_LS_BFX9 U12 ( .A(n83), .Z(n8) );
  HS65_LS_IVX9 U13 ( .A(reset), .Z(n83) );
  HS65_LS_IVX9 U14 ( .A(n161), .Z(n85) );
  HS65_LS_IVX9 U15 ( .A(n162), .Z(n84) );
  HS65_LS_NAND3X5 U16 ( .A(wr_ena), .B(n86), .C(wr_addr[0]), .Z(n161) );
  HS65_LS_IVX9 U17 ( .A(wr_addr[0]), .Z(n89) );
  HS65_LS_NAND3X5 U18 ( .A(n89), .B(n86), .C(wr_ena), .Z(n162) );
  HS65_LS_IVX9 U19 ( .A(n160), .Z(n88) );
  HS65_LS_IVX9 U20 ( .A(n159), .Z(n87) );
  HS65_LS_NAND3X5 U21 ( .A(wr_ena), .B(n89), .C(wr_addr[1]), .Z(n160) );
  HS65_LS_NOR2X6 U22 ( .A(n90), .B(rd_addr[1]), .Z(n157) );
  HS65_LS_NOR2X6 U23 ( .A(rd_addr[0]), .B(rd_addr[1]), .Z(n158) );
  HS65_LS_IVX9 U24 ( .A(wr_addr[1]), .Z(n86) );
  HS65_LS_NAND3X5 U25 ( .A(wr_addr[0]), .B(wr_ena), .C(wr_addr[1]), .Z(n159)
         );
  HS65_LS_AND2X4 U26 ( .A(rd_addr[1]), .B(n90), .Z(n156) );
  HS65_LS_IVX9 U27 ( .A(rd_addr[0]), .Z(n90) );
  HS65_LS_AND2X4 U28 ( .A(rd_addr[1]), .B(rd_addr[0]), .Z(n155) );
  HS65_LS_MX41X7 U29 ( .D0(n158), .S0(\mem[0][0] ), .D1(n157), .S1(\mem[1][0] ), .D2(n156), .S2(\mem[2][0] ), .D3(n155), .S3(\mem[3][0] ), .Z(N32) );
  HS65_LS_MX41X7 U30 ( .D0(n158), .S0(\mem[0][1] ), .D1(n157), .S1(\mem[1][1] ), .D2(n156), .S2(\mem[2][1] ), .D3(n155), .S3(\mem[3][1] ), .Z(N31) );
  HS65_LS_MX41X7 U31 ( .D0(n158), .S0(\mem[0][2] ), .D1(n157), .S1(\mem[1][2] ), .D2(n156), .S2(\mem[2][2] ), .D3(n155), .S3(\mem[3][2] ), .Z(N30) );
  HS65_LS_MX41X7 U32 ( .D0(n158), .S0(\mem[0][3] ), .D1(n157), .S1(\mem[1][3] ), .D2(n156), .S2(\mem[2][3] ), .D3(n155), .S3(\mem[3][3] ), .Z(N29) );
  HS65_LS_MX41X7 U33 ( .D0(n158), .S0(\mem[0][4] ), .D1(n157), .S1(\mem[1][4] ), .D2(n156), .S2(\mem[2][4] ), .D3(n155), .S3(\mem[3][4] ), .Z(N28) );
  HS65_LS_MX41X7 U34 ( .D0(n158), .S0(\mem[0][5] ), .D1(n157), .S1(\mem[1][5] ), .D2(n156), .S2(\mem[2][5] ), .D3(n155), .S3(\mem[3][5] ), .Z(N27) );
  HS65_LS_MX41X7 U35 ( .D0(n158), .S0(\mem[0][6] ), .D1(n157), .S1(\mem[1][6] ), .D2(n156), .S2(\mem[2][6] ), .D3(n155), .S3(\mem[3][6] ), .Z(N26) );
  HS65_LS_MX41X7 U36 ( .D0(n158), .S0(\mem[0][7] ), .D1(n157), .S1(\mem[1][7] ), .D2(n156), .S2(\mem[2][7] ), .D3(n155), .S3(\mem[3][7] ), .Z(N25) );
  HS65_LS_MX41X7 U37 ( .D0(n158), .S0(\mem[0][8] ), .D1(n157), .S1(\mem[1][8] ), .D2(n156), .S2(\mem[2][8] ), .D3(n155), .S3(\mem[3][8] ), .Z(N24) );
  HS65_LS_MX41X7 U38 ( .D0(n158), .S0(\mem[0][9] ), .D1(n157), .S1(\mem[1][9] ), .D2(n156), .S2(\mem[2][9] ), .D3(n155), .S3(\mem[3][9] ), .Z(N23) );
  HS65_LS_MX41X7 U39 ( .D0(n158), .S0(\mem[0][10] ), .D1(n157), .S1(
        \mem[1][10] ), .D2(n156), .S2(\mem[2][10] ), .D3(n155), .S3(
        \mem[3][10] ), .Z(N22) );
  HS65_LS_MX41X7 U40 ( .D0(n158), .S0(\mem[0][11] ), .D1(n157), .S1(
        \mem[1][11] ), .D2(n156), .S2(\mem[2][11] ), .D3(n155), .S3(
        \mem[3][11] ), .Z(N21) );
  HS65_LS_MX41X7 U41 ( .D0(n158), .S0(\mem[0][12] ), .D1(n157), .S1(
        \mem[1][12] ), .D2(n156), .S2(\mem[2][12] ), .D3(n155), .S3(
        \mem[3][12] ), .Z(N20) );
  HS65_LS_MX41X7 U42 ( .D0(n158), .S0(\mem[0][13] ), .D1(n157), .S1(
        \mem[1][13] ), .D2(n156), .S2(\mem[2][13] ), .D3(n155), .S3(
        \mem[3][13] ), .Z(N19) );
  HS65_LS_MX41X7 U43 ( .D0(n158), .S0(\mem[0][14] ), .D1(n157), .S1(
        \mem[1][14] ), .D2(n156), .S2(\mem[2][14] ), .D3(n155), .S3(
        \mem[3][14] ), .Z(N18) );
  HS65_LS_MX41X7 U44 ( .D0(n158), .S0(\mem[0][15] ), .D1(n157), .S1(
        \mem[1][15] ), .D2(n156), .S2(\mem[2][15] ), .D3(n155), .S3(
        \mem[3][15] ), .Z(N17) );
  HS65_LS_AO22X9 U45 ( .A(wr_data[0]), .B(n85), .C(n161), .D(\mem[1][0] ), .Z(
        n138) );
  HS65_LS_AO22X9 U46 ( .A(wr_data[1]), .B(n85), .C(n161), .D(\mem[1][1] ), .Z(
        n137) );
  HS65_LS_AO22X9 U47 ( .A(wr_data[2]), .B(n85), .C(n161), .D(\mem[1][2] ), .Z(
        n136) );
  HS65_LS_AO22X9 U48 ( .A(wr_data[3]), .B(n85), .C(n161), .D(\mem[1][3] ), .Z(
        n135) );
  HS65_LS_AO22X9 U49 ( .A(wr_data[4]), .B(n85), .C(n161), .D(\mem[1][4] ), .Z(
        n134) );
  HS65_LS_AO22X9 U50 ( .A(wr_data[5]), .B(n85), .C(n161), .D(\mem[1][5] ), .Z(
        n133) );
  HS65_LS_AO22X9 U51 ( .A(wr_data[6]), .B(n85), .C(n161), .D(\mem[1][6] ), .Z(
        n132) );
  HS65_LS_AO22X9 U52 ( .A(wr_data[7]), .B(n85), .C(n161), .D(\mem[1][7] ), .Z(
        n131) );
  HS65_LS_AO22X9 U53 ( .A(wr_data[8]), .B(n85), .C(n161), .D(\mem[1][8] ), .Z(
        n130) );
  HS65_LS_AO22X9 U54 ( .A(wr_data[9]), .B(n85), .C(n161), .D(\mem[1][9] ), .Z(
        n129) );
  HS65_LS_AO22X9 U55 ( .A(wr_data[10]), .B(n85), .C(n161), .D(\mem[1][10] ), 
        .Z(n128) );
  HS65_LS_AO22X9 U56 ( .A(wr_data[11]), .B(n85), .C(n161), .D(\mem[1][11] ), 
        .Z(n127) );
  HS65_LS_AO22X9 U57 ( .A(wr_data[12]), .B(n85), .C(n161), .D(\mem[1][12] ), 
        .Z(n126) );
  HS65_LS_AO22X9 U58 ( .A(wr_data[13]), .B(n85), .C(n161), .D(\mem[1][13] ), 
        .Z(n125) );
  HS65_LS_AO22X9 U59 ( .A(wr_data[14]), .B(n85), .C(n161), .D(\mem[1][14] ), 
        .Z(n124) );
  HS65_LS_AO22X9 U60 ( .A(wr_data[15]), .B(n85), .C(n161), .D(\mem[1][15] ), 
        .Z(n123) );
  HS65_LS_AO22X9 U61 ( .A(wr_data[0]), .B(n88), .C(n160), .D(\mem[2][0] ), .Z(
        n122) );
  HS65_LS_AO22X9 U62 ( .A(wr_data[1]), .B(n88), .C(n160), .D(\mem[2][1] ), .Z(
        n121) );
  HS65_LS_AO22X9 U63 ( .A(wr_data[2]), .B(n88), .C(n160), .D(\mem[2][2] ), .Z(
        n120) );
  HS65_LS_AO22X9 U64 ( .A(wr_data[3]), .B(n88), .C(n160), .D(\mem[2][3] ), .Z(
        n119) );
  HS65_LS_AO22X9 U65 ( .A(wr_data[4]), .B(n88), .C(n160), .D(\mem[2][4] ), .Z(
        n118) );
  HS65_LS_AO22X9 U66 ( .A(wr_data[5]), .B(n88), .C(n160), .D(\mem[2][5] ), .Z(
        n117) );
  HS65_LS_AO22X9 U67 ( .A(wr_data[6]), .B(n88), .C(n160), .D(\mem[2][6] ), .Z(
        n116) );
  HS65_LS_AO22X9 U68 ( .A(wr_data[7]), .B(n88), .C(n160), .D(\mem[2][7] ), .Z(
        n115) );
  HS65_LS_AO22X9 U69 ( .A(wr_data[8]), .B(n88), .C(n160), .D(\mem[2][8] ), .Z(
        n114) );
  HS65_LS_AO22X9 U70 ( .A(wr_data[9]), .B(n88), .C(n160), .D(\mem[2][9] ), .Z(
        n113) );
  HS65_LS_AO22X9 U71 ( .A(wr_data[10]), .B(n88), .C(n160), .D(\mem[2][10] ), 
        .Z(n112) );
  HS65_LS_AO22X9 U72 ( .A(wr_data[11]), .B(n88), .C(n160), .D(\mem[2][11] ), 
        .Z(n111) );
  HS65_LS_AO22X9 U73 ( .A(wr_data[12]), .B(n88), .C(n160), .D(\mem[2][12] ), 
        .Z(n110) );
  HS65_LS_AO22X9 U74 ( .A(wr_data[13]), .B(n88), .C(n160), .D(\mem[2][13] ), 
        .Z(n109) );
  HS65_LS_AO22X9 U75 ( .A(wr_data[14]), .B(n88), .C(n160), .D(\mem[2][14] ), 
        .Z(n108) );
  HS65_LS_AO22X9 U76 ( .A(wr_data[15]), .B(n88), .C(n160), .D(\mem[2][15] ), 
        .Z(n107) );
  HS65_LS_AO22X9 U77 ( .A(n84), .B(wr_data[0]), .C(n162), .D(\mem[0][0] ), .Z(
        n154) );
  HS65_LS_AO22X9 U78 ( .A(n84), .B(wr_data[1]), .C(n162), .D(\mem[0][1] ), .Z(
        n153) );
  HS65_LS_AO22X9 U79 ( .A(n84), .B(wr_data[2]), .C(n162), .D(\mem[0][2] ), .Z(
        n152) );
  HS65_LS_AO22X9 U80 ( .A(n84), .B(wr_data[3]), .C(n162), .D(\mem[0][3] ), .Z(
        n151) );
  HS65_LS_AO22X9 U81 ( .A(n84), .B(wr_data[4]), .C(n162), .D(\mem[0][4] ), .Z(
        n150) );
  HS65_LS_AO22X9 U82 ( .A(n84), .B(wr_data[5]), .C(n162), .D(\mem[0][5] ), .Z(
        n149) );
  HS65_LS_AO22X9 U83 ( .A(n84), .B(wr_data[6]), .C(n162), .D(\mem[0][6] ), .Z(
        n148) );
  HS65_LS_AO22X9 U84 ( .A(n84), .B(wr_data[7]), .C(n162), .D(\mem[0][7] ), .Z(
        n147) );
  HS65_LS_AO22X9 U85 ( .A(n84), .B(wr_data[8]), .C(n162), .D(\mem[0][8] ), .Z(
        n146) );
  HS65_LS_AO22X9 U86 ( .A(n84), .B(wr_data[9]), .C(n162), .D(\mem[0][9] ), .Z(
        n145) );
  HS65_LS_AO22X9 U87 ( .A(n84), .B(wr_data[10]), .C(n162), .D(\mem[0][10] ), 
        .Z(n144) );
  HS65_LS_AO22X9 U88 ( .A(n84), .B(wr_data[11]), .C(n162), .D(\mem[0][11] ), 
        .Z(n143) );
  HS65_LS_AO22X9 U89 ( .A(n84), .B(wr_data[12]), .C(n162), .D(\mem[0][12] ), 
        .Z(n142) );
  HS65_LS_AO22X9 U90 ( .A(n84), .B(wr_data[13]), .C(n162), .D(\mem[0][13] ), 
        .Z(n141) );
  HS65_LS_AO22X9 U91 ( .A(n84), .B(wr_data[14]), .C(n162), .D(\mem[0][14] ), 
        .Z(n140) );
  HS65_LS_AO22X9 U92 ( .A(n84), .B(wr_data[15]), .C(n162), .D(\mem[0][15] ), 
        .Z(n139) );
  HS65_LS_AO22X9 U93 ( .A(wr_data[0]), .B(n87), .C(n159), .D(\mem[3][0] ), .Z(
        n106) );
  HS65_LS_AO22X9 U94 ( .A(wr_data[1]), .B(n87), .C(n159), .D(\mem[3][1] ), .Z(
        n105) );
  HS65_LS_AO22X9 U95 ( .A(wr_data[2]), .B(n87), .C(n159), .D(\mem[3][2] ), .Z(
        n104) );
  HS65_LS_AO22X9 U96 ( .A(wr_data[3]), .B(n87), .C(n159), .D(\mem[3][3] ), .Z(
        n103) );
  HS65_LS_AO22X9 U97 ( .A(wr_data[4]), .B(n87), .C(n159), .D(\mem[3][4] ), .Z(
        n102) );
  HS65_LS_AO22X9 U98 ( .A(wr_data[5]), .B(n87), .C(n159), .D(\mem[3][5] ), .Z(
        n101) );
  HS65_LS_AO22X9 U99 ( .A(wr_data[6]), .B(n87), .C(n159), .D(\mem[3][6] ), .Z(
        n100) );
  HS65_LS_AO22X9 U100 ( .A(wr_data[7]), .B(n87), .C(n159), .D(\mem[3][7] ), 
        .Z(n99) );
  HS65_LS_AO22X9 U101 ( .A(wr_data[8]), .B(n87), .C(n159), .D(\mem[3][8] ), 
        .Z(n98) );
  HS65_LS_AO22X9 U102 ( .A(wr_data[9]), .B(n87), .C(n159), .D(\mem[3][9] ), 
        .Z(n97) );
  HS65_LS_AO22X9 U103 ( .A(wr_data[10]), .B(n87), .C(n159), .D(\mem[3][10] ), 
        .Z(n96) );
  HS65_LS_AO22X9 U104 ( .A(wr_data[11]), .B(n87), .C(n159), .D(\mem[3][11] ), 
        .Z(n95) );
  HS65_LS_AO22X9 U105 ( .A(wr_data[12]), .B(n87), .C(n159), .D(\mem[3][12] ), 
        .Z(n94) );
  HS65_LS_AO22X9 U106 ( .A(wr_data[13]), .B(n87), .C(n159), .D(\mem[3][13] ), 
        .Z(n93) );
  HS65_LS_AO22X9 U107 ( .A(wr_data[14]), .B(n87), .C(n159), .D(\mem[3][14] ), 
        .Z(n92) );
  HS65_LS_AO22X9 U108 ( .A(wr_data[15]), .B(n87), .C(n159), .D(\mem[3][15] ), 
        .Z(n91) );
endmodule


module dma_sdp_DATA64_ADDR2_1 ( clk, reset, ren, wen, waddr, wdata, raddr, 
        rdata );
  input [2:0] ren;
  input [2:0] wen;
  input [1:0] waddr;
  input [63:0] wdata;
  input [1:0] raddr;
  output [63:0] rdata;
  input clk, reset;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n41, n42, n43, n44, n45, n46, n47, n48;
  wire   [2:0] sel_out;
  wire   [15:0] rdata0;
  wire   [31:0] rdata1;
  wire   [15:0] rdata2;

  HS65_LS_DFPRQX9 \sel_out_reg[2]  ( .D(ren[2]), .CP(clk), .RN(n5), .Q(
        sel_out[2]) );
  HS65_LS_DFPRQX9 \sel_out_reg[1]  ( .D(ren[1]), .CP(clk), .RN(n5), .Q(
        sel_out[1]) );
  HS65_LS_DFPRQX9 \sel_out_reg[0]  ( .D(ren[0]), .CP(clk), .RN(n5), .Q(
        sel_out[0]) );
  bram_DATA16_ADDR2_2 dma0 ( .clk(clk), .reset(reset), .rd_addr(raddr), 
        .wr_addr(waddr), .wr_data(wdata[63:48]), .wr_ena(wen[2]), .rd_data(
        rdata0) );
  bram_DATA32_ADDR2_1 dma1 ( .clk(clk), .reset(reset), .rd_addr(raddr), 
        .wr_addr(waddr), .wr_data(wdata[47:16]), .wr_ena(wen[1]), .rd_data(
        rdata1) );
  bram_DATA16_ADDR2_1 dma2 ( .clk(clk), .reset(reset), .rd_addr(raddr), 
        .wr_addr(waddr), .wr_data(wdata[15:0]), .wr_ena(wen[0]), .rd_data(
        rdata2) );
  HS65_LS_NAND3X5 U3 ( .A(sel_out[2]), .B(sel_out[1]), .C(sel_out[0]), .Z(n46)
         );
  HS65_LS_IVX9 U4 ( .A(reset), .Z(n5) );
  HS65_LS_NOR2X6 U5 ( .A(n2), .B(n13), .Z(rdata[40]) );
  HS65_LS_NOR2X6 U6 ( .A(n2), .B(n12), .Z(rdata[41]) );
  HS65_LS_NOR2X6 U7 ( .A(n2), .B(n11), .Z(rdata[42]) );
  HS65_LS_NOR2X6 U8 ( .A(n2), .B(n10), .Z(rdata[43]) );
  HS65_LS_NOR2X6 U9 ( .A(n2), .B(n9), .Z(rdata[44]) );
  HS65_LS_NOR2X6 U10 ( .A(n2), .B(n8), .Z(rdata[45]) );
  HS65_LS_NOR2X6 U11 ( .A(n2), .B(n14), .Z(rdata[39]) );
  HS65_LS_BFX9 U12 ( .A(n46), .Z(n2) );
  HS65_LS_NOR2X6 U13 ( .A(n2), .B(n15), .Z(rdata[38]) );
  HS65_LS_NOR2X6 U14 ( .A(n3), .B(n19), .Z(rdata[34]) );
  HS65_LS_NOR2X6 U15 ( .A(n2), .B(n18), .Z(rdata[35]) );
  HS65_LS_NOR2X6 U16 ( .A(n3), .B(n17), .Z(rdata[36]) );
  HS65_LS_NOR2X6 U17 ( .A(n2), .B(n16), .Z(rdata[37]) );
  HS65_LS_NOR2X6 U18 ( .A(n3), .B(n20), .Z(rdata[33]) );
  HS65_LS_BFX9 U19 ( .A(n46), .Z(n3) );
  HS65_LS_BFX9 U20 ( .A(n46), .Z(n1) );
  HS65_LS_BFX9 U21 ( .A(n46), .Z(n4) );
  HS65_LS_IVX9 U22 ( .A(n45), .Z(n42) );
  HS65_LS_NOR2X6 U23 ( .A(n2), .B(n7), .Z(rdata[46]) );
  HS65_LS_NOR2X6 U24 ( .A(n2), .B(n6), .Z(rdata[47]) );
  HS65_LS_NAND3X5 U25 ( .A(n44), .B(n43), .C(sel_out[1]), .Z(n45) );
  HS65_LS_IVX9 U26 ( .A(sel_out[0]), .Z(n44) );
  HS65_LS_IVX9 U27 ( .A(sel_out[2]), .Z(n43) );
  HS65_LS_OAI22X6 U28 ( .A(n45), .B(n19), .C(n1), .D(n35), .Z(rdata[18]) );
  HS65_LS_IVX9 U29 ( .A(rdata1[2]), .Z(n35) );
  HS65_LS_OAI22X6 U30 ( .A(n45), .B(n18), .C(n1), .D(n34), .Z(rdata[19]) );
  HS65_LS_IVX9 U31 ( .A(rdata1[3]), .Z(n34) );
  HS65_LS_OAI22X6 U32 ( .A(n45), .B(n17), .C(n1), .D(n33), .Z(rdata[20]) );
  HS65_LS_IVX9 U33 ( .A(rdata1[4]), .Z(n33) );
  HS65_LS_OAI22X6 U34 ( .A(n45), .B(n16), .C(n1), .D(n32), .Z(rdata[21]) );
  HS65_LS_IVX9 U35 ( .A(rdata1[5]), .Z(n32) );
  HS65_LS_OAI22X6 U36 ( .A(n45), .B(n15), .C(n31), .D(n3), .Z(rdata[22]) );
  HS65_LS_IVX9 U37 ( .A(rdata1[6]), .Z(n31) );
  HS65_LS_OAI22X6 U38 ( .A(n45), .B(n14), .C(n30), .D(n3), .Z(rdata[23]) );
  HS65_LS_IVX9 U39 ( .A(rdata1[7]), .Z(n30) );
  HS65_LS_OAI22X6 U40 ( .A(n45), .B(n13), .C(n29), .D(n3), .Z(rdata[24]) );
  HS65_LS_IVX9 U41 ( .A(rdata1[8]), .Z(n29) );
  HS65_LS_OAI22X6 U42 ( .A(n45), .B(n12), .C(n28), .D(n3), .Z(rdata[25]) );
  HS65_LS_IVX9 U43 ( .A(rdata1[9]), .Z(n28) );
  HS65_LS_OAI22X6 U44 ( .A(n45), .B(n11), .C(n1), .D(n27), .Z(rdata[26]) );
  HS65_LS_IVX9 U45 ( .A(rdata1[10]), .Z(n27) );
  HS65_LS_OAI22X6 U46 ( .A(n45), .B(n10), .C(n1), .D(n26), .Z(rdata[27]) );
  HS65_LS_IVX9 U47 ( .A(rdata1[11]), .Z(n26) );
  HS65_LS_OAI22X6 U48 ( .A(n45), .B(n20), .C(n1), .D(n36), .Z(rdata[17]) );
  HS65_LS_IVX9 U49 ( .A(rdata1[1]), .Z(n36) );
  HS65_LS_NOR2X6 U50 ( .A(n3), .B(n21), .Z(rdata[32]) );
  HS65_LS_NOR2AX3 U51 ( .A(rdata0[15]), .B(n3), .Z(rdata[63]) );
  HS65_LS_IVX9 U52 ( .A(rdata1[18]), .Z(n19) );
  HS65_LS_IVX9 U53 ( .A(rdata1[19]), .Z(n18) );
  HS65_LS_IVX9 U54 ( .A(rdata1[17]), .Z(n20) );
  HS65_LS_NOR2AX3 U55 ( .A(rdata0[3]), .B(n3), .Z(rdata[51]) );
  HS65_LS_NOR2AX3 U56 ( .A(rdata0[4]), .B(n4), .Z(rdata[52]) );
  HS65_LS_NOR2AX3 U57 ( .A(rdata0[7]), .B(n4), .Z(rdata[55]) );
  HS65_LS_NOR2AX3 U58 ( .A(rdata0[8]), .B(n4), .Z(rdata[56]) );
  HS65_LS_NOR2AX3 U59 ( .A(rdata0[10]), .B(n4), .Z(rdata[58]) );
  HS65_LS_NOR2AX3 U60 ( .A(rdata0[1]), .B(n3), .Z(rdata[49]) );
  HS65_LS_NOR2AX3 U61 ( .A(rdata0[2]), .B(n3), .Z(rdata[50]) );
  HS65_LS_NOR2AX3 U62 ( .A(rdata0[5]), .B(n4), .Z(rdata[53]) );
  HS65_LS_NOR2AX3 U63 ( .A(rdata0[6]), .B(n4), .Z(rdata[54]) );
  HS65_LS_NOR2AX3 U64 ( .A(rdata0[9]), .B(n4), .Z(rdata[57]) );
  HS65_LS_NOR2AX3 U65 ( .A(rdata0[11]), .B(n4), .Z(rdata[59]) );
  HS65_LS_NOR2AX3 U66 ( .A(rdata0[14]), .B(n4), .Z(rdata[62]) );
  HS65_LS_OAI31X5 U67 ( .A(n44), .B(sel_out[2]), .C(sel_out[1]), .D(n2), .Z(
        n47) );
  HS65_LS_NOR3X4 U68 ( .A(sel_out[0]), .B(sel_out[1]), .C(n43), .Z(n48) );
  HS65_LS_OAI22X6 U69 ( .A(n45), .B(n9), .C(n1), .D(n25), .Z(rdata[28]) );
  HS65_LS_IVX9 U70 ( .A(rdata1[12]), .Z(n25) );
  HS65_LS_OAI22X6 U71 ( .A(n45), .B(n8), .C(n1), .D(n24), .Z(rdata[29]) );
  HS65_LS_IVX9 U72 ( .A(rdata1[13]), .Z(n24) );
  HS65_LS_OAI22X6 U73 ( .A(n45), .B(n7), .C(n1), .D(n23), .Z(rdata[30]) );
  HS65_LS_IVX9 U74 ( .A(rdata1[14]), .Z(n23) );
  HS65_LS_OAI22X6 U75 ( .A(n45), .B(n6), .C(n1), .D(n22), .Z(rdata[31]) );
  HS65_LS_IVX9 U76 ( .A(rdata1[15]), .Z(n22) );
  HS65_LS_OAI22X6 U77 ( .A(n45), .B(n21), .C(n1), .D(n41), .Z(rdata[16]) );
  HS65_LS_IVX9 U78 ( .A(rdata1[0]), .Z(n41) );
  HS65_LS_NOR2AX3 U79 ( .A(rdata0[0]), .B(n3), .Z(rdata[48]) );
  HS65_LS_IVX9 U80 ( .A(rdata1[20]), .Z(n17) );
  HS65_LS_IVX9 U81 ( .A(rdata1[21]), .Z(n16) );
  HS65_LS_IVX9 U82 ( .A(rdata1[22]), .Z(n15) );
  HS65_LS_IVX9 U83 ( .A(rdata1[23]), .Z(n14) );
  HS65_LS_IVX9 U84 ( .A(rdata1[24]), .Z(n13) );
  HS65_LS_IVX9 U85 ( .A(rdata1[25]), .Z(n12) );
  HS65_LS_IVX9 U86 ( .A(rdata1[26]), .Z(n11) );
  HS65_LS_IVX9 U87 ( .A(rdata1[27]), .Z(n10) );
  HS65_LS_IVX9 U88 ( .A(rdata1[28]), .Z(n9) );
  HS65_LS_IVX9 U89 ( .A(rdata1[29]), .Z(n8) );
  HS65_LS_IVX9 U90 ( .A(rdata1[30]), .Z(n7) );
  HS65_LS_IVX9 U91 ( .A(rdata1[31]), .Z(n6) );
  HS65_LS_IVX9 U92 ( .A(rdata1[16]), .Z(n21) );
  HS65_LS_AO222X4 U93 ( .A(rdata0[0]), .B(n48), .C(rdata1[0]), .D(n42), .E(
        rdata2[0]), .F(n47), .Z(rdata[0]) );
  HS65_LS_AO222X4 U94 ( .A(rdata0[1]), .B(n48), .C(rdata1[1]), .D(n42), .E(
        rdata2[1]), .F(n47), .Z(rdata[1]) );
  HS65_LS_AO222X4 U95 ( .A(rdata0[2]), .B(n48), .C(rdata1[2]), .D(n42), .E(
        rdata2[2]), .F(n47), .Z(rdata[2]) );
  HS65_LS_AO222X4 U96 ( .A(rdata0[3]), .B(n48), .C(rdata1[3]), .D(n42), .E(
        rdata2[3]), .F(n47), .Z(rdata[3]) );
  HS65_LS_AO222X4 U97 ( .A(rdata0[4]), .B(n48), .C(rdata1[4]), .D(n42), .E(
        rdata2[4]), .F(n47), .Z(rdata[4]) );
  HS65_LS_AO222X4 U98 ( .A(rdata0[5]), .B(n48), .C(rdata1[5]), .D(n42), .E(
        rdata2[5]), .F(n47), .Z(rdata[5]) );
  HS65_LS_AO222X4 U99 ( .A(rdata0[6]), .B(n48), .C(rdata1[6]), .D(n42), .E(
        rdata2[6]), .F(n47), .Z(rdata[6]) );
  HS65_LS_AO222X4 U100 ( .A(rdata0[7]), .B(n48), .C(rdata1[7]), .D(n42), .E(
        rdata2[7]), .F(n47), .Z(rdata[7]) );
  HS65_LS_AO222X4 U101 ( .A(rdata0[8]), .B(n48), .C(rdata1[8]), .D(n42), .E(
        rdata2[8]), .F(n47), .Z(rdata[8]) );
  HS65_LS_AO222X4 U102 ( .A(rdata0[9]), .B(n48), .C(rdata1[9]), .D(n42), .E(
        rdata2[9]), .F(n47), .Z(rdata[9]) );
  HS65_LS_AO222X4 U103 ( .A(rdata0[10]), .B(n48), .C(rdata1[10]), .D(n42), .E(
        rdata2[10]), .F(n47), .Z(rdata[10]) );
  HS65_LS_AO222X4 U104 ( .A(rdata0[11]), .B(n48), .C(rdata1[11]), .D(n42), .E(
        rdata2[11]), .F(n47), .Z(rdata[11]) );
  HS65_LS_AO222X4 U105 ( .A(rdata0[12]), .B(n48), .C(rdata1[12]), .D(n42), .E(
        rdata2[12]), .F(n47), .Z(rdata[12]) );
  HS65_LS_AO222X4 U106 ( .A(rdata0[13]), .B(n48), .C(rdata1[13]), .D(n42), .E(
        rdata2[13]), .F(n47), .Z(rdata[13]) );
  HS65_LS_AO222X4 U107 ( .A(rdata0[14]), .B(n48), .C(rdata1[14]), .D(n42), .E(
        rdata2[14]), .F(n47), .Z(rdata[14]) );
  HS65_LS_AO222X4 U108 ( .A(rdata0[15]), .B(n48), .C(rdata1[15]), .D(n42), .E(
        rdata2[15]), .F(n47), .Z(rdata[15]) );
  HS65_LS_NOR2AX3 U109 ( .A(rdata0[12]), .B(n4), .Z(rdata[60]) );
  HS65_LS_NOR2AX3 U110 ( .A(rdata0[13]), .B(n4), .Z(rdata[61]) );
endmodule


module bram_DATA5_ADDR3_1 ( clk, reset, rd_addr, wr_addr, wr_data, wr_ena, 
        rd_data );
  input [2:0] rd_addr;
  input [2:0] wr_addr;
  input [4:0] wr_data;
  output [4:0] rd_data;
  input clk, reset, wr_ena;
  wire   \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N34,
         N35, N36, N37, N38, n1, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218;

  HS65_LS_DFPRQX9 \mem_reg[5][4]  ( .D(n131), .CP(clk), .RN(n1), .Q(
        \mem[5][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[5][3]  ( .D(n132), .CP(clk), .RN(n1), .Q(
        \mem[5][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[5][2]  ( .D(n133), .CP(clk), .RN(n1), .Q(
        \mem[5][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[5][1]  ( .D(n134), .CP(clk), .RN(n1), .Q(
        \mem[5][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[5][0]  ( .D(n135), .CP(clk), .RN(n22), .Q(
        \mem[5][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[4][4]  ( .D(n136), .CP(clk), .RN(n22), .Q(
        \mem[4][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[4][3]  ( .D(n137), .CP(clk), .RN(n22), .Q(
        \mem[4][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[4][2]  ( .D(n138), .CP(clk), .RN(n22), .Q(
        \mem[4][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[4][1]  ( .D(n139), .CP(clk), .RN(n22), .Q(
        \mem[4][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[4][0]  ( .D(n140), .CP(clk), .RN(n22), .Q(
        \mem[4][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][4]  ( .D(n151), .CP(clk), .RN(n22), .Q(
        \mem[1][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][3]  ( .D(n152), .CP(clk), .RN(n22), .Q(
        \mem[1][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][2]  ( .D(n153), .CP(clk), .RN(n22), .Q(
        \mem[1][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][1]  ( .D(n154), .CP(clk), .RN(n22), .Q(
        \mem[1][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[1][0]  ( .D(n155), .CP(clk), .RN(n22), .Q(
        \mem[1][0] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][4]  ( .D(n156), .CP(clk), .RN(n22), .Q(
        \mem[0][4] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][3]  ( .D(n157), .CP(clk), .RN(n1), .Q(
        \mem[0][3] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][2]  ( .D(n158), .CP(clk), .RN(n1), .Q(
        \mem[0][2] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][1]  ( .D(n159), .CP(clk), .RN(n1), .Q(
        \mem[0][1] ) );
  HS65_LS_DFPRQX9 \mem_reg[0][0]  ( .D(n160), .CP(clk), .RN(n1), .Q(
        \mem[0][0] ) );
  HS65_LS_DFPRQX9 \rd_data_reg[4]  ( .D(N34), .CP(clk), .RN(n1), .Q(rd_data[4]) );
  HS65_LS_DFPRQX9 \rd_data_reg[3]  ( .D(N35), .CP(clk), .RN(n1), .Q(rd_data[3]) );
  HS65_LS_DFPRQX9 \rd_data_reg[2]  ( .D(N36), .CP(clk), .RN(n1), .Q(rd_data[2]) );
  HS65_LS_DFPRQX9 \rd_data_reg[1]  ( .D(N37), .CP(clk), .RN(n1), .Q(rd_data[1]) );
  HS65_LS_DFPRQX9 \rd_data_reg[0]  ( .D(N38), .CP(clk), .RN(n1), .Q(rd_data[0]) );
  HS65_LS_DFPRQNX9 \mem_reg[7][4]  ( .D(n121), .CP(clk), .RN(n23), .QN(n218)
         );
  HS65_LS_DFPRQNX9 \mem_reg[7][3]  ( .D(n122), .CP(clk), .RN(n22), .QN(n217)
         );
  HS65_LS_DFPRQNX9 \mem_reg[7][2]  ( .D(n123), .CP(clk), .RN(n24), .QN(n216)
         );
  HS65_LS_DFPRQNX9 \mem_reg[7][1]  ( .D(n124), .CP(clk), .RN(n24), .QN(n215)
         );
  HS65_LS_DFPRQNX9 \mem_reg[7][0]  ( .D(n125), .CP(clk), .RN(n24), .QN(n214)
         );
  HS65_LS_DFPRQNX9 \mem_reg[3][4]  ( .D(n141), .CP(clk), .RN(n23), .QN(n208)
         );
  HS65_LS_DFPRQNX9 \mem_reg[3][3]  ( .D(n142), .CP(clk), .RN(n23), .QN(n207)
         );
  HS65_LS_DFPRQNX9 \mem_reg[3][2]  ( .D(n143), .CP(clk), .RN(n23), .QN(n206)
         );
  HS65_LS_DFPRQNX9 \mem_reg[3][1]  ( .D(n144), .CP(clk), .RN(n23), .QN(n205)
         );
  HS65_LS_DFPRQNX9 \mem_reg[3][0]  ( .D(n145), .CP(clk), .RN(n23), .QN(n204)
         );
  HS65_LS_DFPRQNX9 \mem_reg[6][4]  ( .D(n126), .CP(clk), .RN(n24), .QN(n213)
         );
  HS65_LS_DFPRQNX9 \mem_reg[6][3]  ( .D(n127), .CP(clk), .RN(n24), .QN(n212)
         );
  HS65_LS_DFPRQNX9 \mem_reg[6][2]  ( .D(n128), .CP(clk), .RN(n23), .QN(n211)
         );
  HS65_LS_DFPRQNX9 \mem_reg[6][1]  ( .D(n129), .CP(clk), .RN(n23), .QN(n210)
         );
  HS65_LS_DFPRQNX9 \mem_reg[6][0]  ( .D(n130), .CP(clk), .RN(n23), .QN(n209)
         );
  HS65_LS_DFPRQNX9 \mem_reg[2][4]  ( .D(n146), .CP(clk), .RN(n23), .QN(n203)
         );
  HS65_LS_DFPRQNX9 \mem_reg[2][3]  ( .D(n147), .CP(clk), .RN(n23), .QN(n202)
         );
  HS65_LS_DFPRQNX9 \mem_reg[2][2]  ( .D(n148), .CP(clk), .RN(n23), .QN(n201)
         );
  HS65_LS_DFPRQNX9 \mem_reg[2][1]  ( .D(n149), .CP(clk), .RN(n23), .QN(n200)
         );
  HS65_LS_DFPRQNX9 \mem_reg[2][0]  ( .D(n150), .CP(clk), .RN(n23), .QN(n199)
         );
  HS65_LS_BFX9 U3 ( .A(n25), .Z(n1) );
  HS65_LS_BFX9 U4 ( .A(n25), .Z(n22) );
  HS65_LS_BFX9 U5 ( .A(n25), .Z(n23) );
  HS65_LS_BFX9 U6 ( .A(n25), .Z(n24) );
  HS65_LS_IVX9 U7 ( .A(reset), .Z(n25) );
  HS65_LS_IVX9 U8 ( .A(n198), .Z(n35) );
  HS65_LS_IVX9 U9 ( .A(n193), .Z(n31) );
  HS65_LS_IVX9 U10 ( .A(n194), .Z(n32) );
  HS65_LS_IVX9 U11 ( .A(n190), .Z(n29) );
  HS65_LS_IVX9 U12 ( .A(n189), .Z(n28) );
  HS65_LS_IVX9 U13 ( .A(n195), .Z(n33) );
  HS65_LS_NAND3X5 U14 ( .A(n37), .B(n36), .C(n197), .Z(n198) );
  HS65_LS_NAND3X5 U15 ( .A(n37), .B(n36), .C(n192), .Z(n193) );
  HS65_LS_IVX9 U16 ( .A(n191), .Z(n30) );
  HS65_LS_IVX9 U17 ( .A(n196), .Z(n34) );
  HS65_LS_NOR3X4 U18 ( .A(n26), .B(rd_addr[1]), .C(n27), .Z(n186) );
  HS65_LS_NOR3X4 U19 ( .A(rd_addr[1]), .B(rd_addr[2]), .C(n26), .Z(n181) );
  HS65_LS_NOR3X4 U20 ( .A(rd_addr[1]), .B(rd_addr[2]), .C(rd_addr[0]), .Z(n180) );
  HS65_LS_NOR3X4 U21 ( .A(rd_addr[0]), .B(rd_addr[1]), .C(n27), .Z(n185) );
  HS65_LS_NAND3X5 U22 ( .A(n26), .B(n27), .C(rd_addr[1]), .Z(n178) );
  HS65_LS_NAND3X5 U23 ( .A(rd_addr[0]), .B(n27), .C(rd_addr[1]), .Z(n177) );
  HS65_LS_NAND3X5 U24 ( .A(rd_addr[1]), .B(n26), .C(rd_addr[2]), .Z(n183) );
  HS65_LS_NAND3X5 U25 ( .A(rd_addr[1]), .B(rd_addr[0]), .C(rd_addr[2]), .Z(
        n182) );
  HS65_LS_OAI22X6 U26 ( .A(n199), .B(n178), .C(n204), .D(n177), .Z(n179) );
  HS65_LS_OAI22X6 U27 ( .A(n200), .B(n178), .C(n205), .D(n177), .Z(n173) );
  HS65_LS_OAI22X6 U28 ( .A(n201), .B(n178), .C(n206), .D(n177), .Z(n169) );
  HS65_LS_OAI22X6 U29 ( .A(n202), .B(n178), .C(n207), .D(n177), .Z(n165) );
  HS65_LS_OAI22X6 U30 ( .A(n203), .B(n178), .C(n208), .D(n177), .Z(n161) );
  HS65_LS_IVX9 U31 ( .A(rd_addr[0]), .Z(n26) );
  HS65_LS_IVX9 U32 ( .A(rd_addr[2]), .Z(n27) );
  HS65_LS_OAI22X6 U33 ( .A(n120), .B(n194), .C(n32), .D(n204), .Z(n145) );
  HS65_LS_OAI22X6 U34 ( .A(n119), .B(n194), .C(n32), .D(n205), .Z(n144) );
  HS65_LS_OAI22X6 U35 ( .A(n118), .B(n194), .C(n32), .D(n206), .Z(n143) );
  HS65_LS_OAI22X6 U36 ( .A(n117), .B(n194), .C(n32), .D(n207), .Z(n142) );
  HS65_LS_OAI22X6 U37 ( .A(n38), .B(n194), .C(n32), .D(n208), .Z(n141) );
  HS65_LS_OAI22X6 U38 ( .A(n120), .B(n190), .C(n29), .D(n209), .Z(n130) );
  HS65_LS_OAI22X6 U39 ( .A(n119), .B(n190), .C(n29), .D(n210), .Z(n129) );
  HS65_LS_OAI22X6 U40 ( .A(n118), .B(n190), .C(n29), .D(n211), .Z(n128) );
  HS65_LS_OAI22X6 U41 ( .A(n117), .B(n190), .C(n29), .D(n212), .Z(n127) );
  HS65_LS_OAI22X6 U42 ( .A(n38), .B(n190), .C(n29), .D(n213), .Z(n126) );
  HS65_LS_OAI22X6 U43 ( .A(n120), .B(n189), .C(n28), .D(n214), .Z(n125) );
  HS65_LS_OAI22X6 U44 ( .A(n119), .B(n189), .C(n28), .D(n215), .Z(n124) );
  HS65_LS_OAI22X6 U45 ( .A(n118), .B(n189), .C(n28), .D(n216), .Z(n123) );
  HS65_LS_OAI22X6 U46 ( .A(n117), .B(n189), .C(n28), .D(n217), .Z(n122) );
  HS65_LS_OAI22X6 U47 ( .A(n38), .B(n189), .C(n28), .D(n218), .Z(n121) );
  HS65_LS_OAI22X6 U48 ( .A(n120), .B(n195), .C(n33), .D(n199), .Z(n150) );
  HS65_LS_OAI22X6 U49 ( .A(n119), .B(n195), .C(n33), .D(n200), .Z(n149) );
  HS65_LS_OAI22X6 U50 ( .A(n118), .B(n195), .C(n33), .D(n201), .Z(n148) );
  HS65_LS_OAI22X6 U51 ( .A(n117), .B(n195), .C(n33), .D(n202), .Z(n147) );
  HS65_LS_OAI22X6 U52 ( .A(n38), .B(n195), .C(n33), .D(n203), .Z(n146) );
  HS65_LS_NAND2X7 U53 ( .A(n188), .B(n187), .Z(N38) );
  HS65_LS_AOI212X4 U54 ( .A(n186), .B(\mem[5][0] ), .C(n185), .D(\mem[4][0] ), 
        .E(n184), .Z(n187) );
  HS65_LS_AOI212X4 U55 ( .A(n181), .B(\mem[1][0] ), .C(n180), .D(\mem[0][0] ), 
        .E(n179), .Z(n188) );
  HS65_LS_OAI22X6 U56 ( .A(n209), .B(n183), .C(n214), .D(n182), .Z(n184) );
  HS65_LS_NAND2X7 U57 ( .A(n176), .B(n175), .Z(N37) );
  HS65_LS_AOI212X4 U58 ( .A(n186), .B(\mem[5][1] ), .C(n185), .D(\mem[4][1] ), 
        .E(n174), .Z(n175) );
  HS65_LS_AOI212X4 U59 ( .A(n181), .B(\mem[1][1] ), .C(n180), .D(\mem[0][1] ), 
        .E(n173), .Z(n176) );
  HS65_LS_OAI22X6 U60 ( .A(n210), .B(n183), .C(n215), .D(n182), .Z(n174) );
  HS65_LS_NAND2X7 U61 ( .A(n172), .B(n171), .Z(N36) );
  HS65_LS_AOI212X4 U62 ( .A(n186), .B(\mem[5][2] ), .C(n185), .D(\mem[4][2] ), 
        .E(n170), .Z(n171) );
  HS65_LS_AOI212X4 U63 ( .A(n181), .B(\mem[1][2] ), .C(n180), .D(\mem[0][2] ), 
        .E(n169), .Z(n172) );
  HS65_LS_OAI22X6 U64 ( .A(n211), .B(n183), .C(n216), .D(n182), .Z(n170) );
  HS65_LS_NAND2X7 U65 ( .A(n168), .B(n167), .Z(N35) );
  HS65_LS_AOI212X4 U66 ( .A(n186), .B(\mem[5][3] ), .C(n185), .D(\mem[4][3] ), 
        .E(n166), .Z(n167) );
  HS65_LS_AOI212X4 U67 ( .A(n181), .B(\mem[1][3] ), .C(n180), .D(\mem[0][3] ), 
        .E(n165), .Z(n168) );
  HS65_LS_OAI22X6 U68 ( .A(n212), .B(n183), .C(n217), .D(n182), .Z(n166) );
  HS65_LS_NAND2X7 U69 ( .A(n164), .B(n163), .Z(N34) );
  HS65_LS_AOI212X4 U70 ( .A(n186), .B(\mem[5][4] ), .C(n185), .D(\mem[4][4] ), 
        .E(n162), .Z(n163) );
  HS65_LS_AOI212X4 U71 ( .A(n181), .B(\mem[1][4] ), .C(n180), .D(\mem[0][4] ), 
        .E(n161), .Z(n164) );
  HS65_LS_OAI22X6 U72 ( .A(n213), .B(n183), .C(n218), .D(n182), .Z(n162) );
  HS65_LS_AO22X9 U73 ( .A(n35), .B(wr_data[0]), .C(n198), .D(\mem[0][0] ), .Z(
        n160) );
  HS65_LS_AO22X9 U74 ( .A(n35), .B(wr_data[1]), .C(n198), .D(\mem[0][1] ), .Z(
        n159) );
  HS65_LS_AO22X9 U75 ( .A(n35), .B(wr_data[2]), .C(n198), .D(\mem[0][2] ), .Z(
        n158) );
  HS65_LS_AO22X9 U76 ( .A(n35), .B(wr_data[3]), .C(n198), .D(\mem[0][3] ), .Z(
        n157) );
  HS65_LS_AO22X9 U77 ( .A(n35), .B(wr_data[4]), .C(n198), .D(\mem[0][4] ), .Z(
        n156) );
  HS65_LS_AO22X9 U78 ( .A(wr_data[0]), .B(n31), .C(n193), .D(\mem[4][0] ), .Z(
        n140) );
  HS65_LS_AO22X9 U79 ( .A(wr_data[1]), .B(n31), .C(n193), .D(\mem[4][1] ), .Z(
        n139) );
  HS65_LS_AO22X9 U80 ( .A(wr_data[2]), .B(n31), .C(n193), .D(\mem[4][2] ), .Z(
        n138) );
  HS65_LS_AO22X9 U81 ( .A(wr_data[3]), .B(n31), .C(n193), .D(\mem[4][3] ), .Z(
        n137) );
  HS65_LS_AO22X9 U82 ( .A(wr_data[4]), .B(n31), .C(n193), .D(\mem[4][4] ), .Z(
        n136) );
  HS65_LS_AO22X9 U83 ( .A(wr_data[0]), .B(n30), .C(n191), .D(\mem[5][0] ), .Z(
        n135) );
  HS65_LS_AO22X9 U84 ( .A(wr_data[1]), .B(n30), .C(n191), .D(\mem[5][1] ), .Z(
        n134) );
  HS65_LS_AO22X9 U85 ( .A(wr_data[2]), .B(n30), .C(n191), .D(\mem[5][2] ), .Z(
        n133) );
  HS65_LS_AO22X9 U86 ( .A(wr_data[3]), .B(n30), .C(n191), .D(\mem[5][3] ), .Z(
        n132) );
  HS65_LS_AO22X9 U87 ( .A(wr_data[4]), .B(n30), .C(n191), .D(\mem[5][4] ), .Z(
        n131) );
  HS65_LS_AO22X9 U88 ( .A(wr_data[0]), .B(n34), .C(n196), .D(\mem[1][0] ), .Z(
        n155) );
  HS65_LS_AO22X9 U89 ( .A(wr_data[1]), .B(n34), .C(n196), .D(\mem[1][1] ), .Z(
        n154) );
  HS65_LS_AO22X9 U90 ( .A(wr_data[2]), .B(n34), .C(n196), .D(\mem[1][2] ), .Z(
        n153) );
  HS65_LS_AO22X9 U91 ( .A(wr_data[3]), .B(n34), .C(n196), .D(\mem[1][3] ), .Z(
        n152) );
  HS65_LS_AO22X9 U92 ( .A(wr_data[4]), .B(n34), .C(n196), .D(\mem[1][4] ), .Z(
        n151) );
  HS65_LS_NAND3X5 U93 ( .A(wr_addr[0]), .B(n197), .C(wr_addr[1]), .Z(n194) );
  HS65_LS_NAND3X5 U94 ( .A(wr_addr[1]), .B(n37), .C(n192), .Z(n190) );
  HS65_LS_NAND3X5 U95 ( .A(wr_addr[1]), .B(wr_addr[0]), .C(n192), .Z(n189) );
  HS65_LS_NAND3X5 U96 ( .A(n197), .B(n37), .C(wr_addr[1]), .Z(n195) );
  HS65_LS_NOR2AX3 U97 ( .A(wr_ena), .B(wr_addr[2]), .Z(n197) );
  HS65_LS_NAND3X5 U98 ( .A(wr_addr[0]), .B(n36), .C(n192), .Z(n191) );
  HS65_LS_NAND3X5 U99 ( .A(n197), .B(n36), .C(wr_addr[0]), .Z(n196) );
  HS65_LS_IVX9 U100 ( .A(wr_addr[0]), .Z(n37) );
  HS65_LS_IVX9 U101 ( .A(wr_data[0]), .Z(n120) );
  HS65_LS_IVX9 U102 ( .A(wr_data[1]), .Z(n119) );
  HS65_LS_IVX9 U103 ( .A(wr_data[2]), .Z(n118) );
  HS65_LS_IVX9 U104 ( .A(wr_data[3]), .Z(n117) );
  HS65_LS_IVX9 U105 ( .A(wr_data[4]), .Z(n38) );
  HS65_LS_IVX9 U106 ( .A(wr_addr[1]), .Z(n36) );
  HS65_LS_AND2X4 U107 ( .A(wr_addr[2]), .B(wr_ena), .Z(n192) );
endmodule


module nAdapter_1 ( na_clk, na_reset, .proc_in({\proc_in[MCMD][1] , 
        \proc_in[MCMD][0] , \proc_in[MADDR][31] , \proc_in[MADDR][30] , 
        \proc_in[MADDR][29] , \proc_in[MADDR][28] , \proc_in[MADDR][27] , 
        \proc_in[MADDR][26] , \proc_in[MADDR][25] , \proc_in[MADDR][24] , 
        \proc_in[MADDR][23] , \proc_in[MADDR][22] , \proc_in[MADDR][21] , 
        \proc_in[MADDR][20] , \proc_in[MADDR][19] , \proc_in[MADDR][18] , 
        \proc_in[MADDR][17] , \proc_in[MADDR][16] , \proc_in[MADDR][15] , 
        \proc_in[MADDR][14] , \proc_in[MADDR][13] , \proc_in[MADDR][12] , 
        \proc_in[MADDR][11] , \proc_in[MADDR][10] , \proc_in[MADDR][9] , 
        \proc_in[MADDR][8] , \proc_in[MADDR][7] , \proc_in[MADDR][6] , 
        \proc_in[MADDR][5] , \proc_in[MADDR][4] , \proc_in[MADDR][3] , 
        \proc_in[MADDR][2] , \proc_in[MADDR][1] , \proc_in[MADDR][0] , 
        \proc_in[MDATA][31] , \proc_in[MDATA][30] , \proc_in[MDATA][29] , 
        \proc_in[MDATA][28] , \proc_in[MDATA][27] , \proc_in[MDATA][26] , 
        \proc_in[MDATA][25] , \proc_in[MDATA][24] , \proc_in[MDATA][23] , 
        \proc_in[MDATA][22] , \proc_in[MDATA][21] , \proc_in[MDATA][20] , 
        \proc_in[MDATA][19] , \proc_in[MDATA][18] , \proc_in[MDATA][17] , 
        \proc_in[MDATA][16] , \proc_in[MDATA][15] , \proc_in[MDATA][14] , 
        \proc_in[MDATA][13] , \proc_in[MDATA][12] , \proc_in[MDATA][11] , 
        \proc_in[MDATA][10] , \proc_in[MDATA][9] , \proc_in[MDATA][8] , 
        \proc_in[MDATA][7] , \proc_in[MDATA][6] , \proc_in[MDATA][5] , 
        \proc_in[MDATA][4] , \proc_in[MDATA][3] , \proc_in[MDATA][2] , 
        \proc_in[MDATA][1] , \proc_in[MDATA][0] }), .proc_out({
        \proc_out[SCMDACCEPT] , \proc_out[SRESP] , \proc_out[SDATA][31] , 
        \proc_out[SDATA][30] , \proc_out[SDATA][29] , \proc_out[SDATA][28] , 
        \proc_out[SDATA][27] , \proc_out[SDATA][26] , \proc_out[SDATA][25] , 
        \proc_out[SDATA][24] , \proc_out[SDATA][23] , \proc_out[SDATA][22] , 
        \proc_out[SDATA][21] , \proc_out[SDATA][20] , \proc_out[SDATA][19] , 
        \proc_out[SDATA][18] , \proc_out[SDATA][17] , \proc_out[SDATA][16] , 
        \proc_out[SDATA][15] , \proc_out[SDATA][14] , \proc_out[SDATA][13] , 
        \proc_out[SDATA][12] , \proc_out[SDATA][11] , \proc_out[SDATA][10] , 
        \proc_out[SDATA][9] , \proc_out[SDATA][8] , \proc_out[SDATA][7] , 
        \proc_out[SDATA][6] , \proc_out[SDATA][5] , \proc_out[SDATA][4] , 
        \proc_out[SDATA][3] , \proc_out[SDATA][2] , \proc_out[SDATA][1] , 
        \proc_out[SDATA][0] }), .spm_in({\spm_in[SCMDACCEPT] , \spm_in[SRESP] , 
        \spm_in[SDATA][63] , \spm_in[SDATA][62] , \spm_in[SDATA][61] , 
        \spm_in[SDATA][60] , \spm_in[SDATA][59] , \spm_in[SDATA][58] , 
        \spm_in[SDATA][57] , \spm_in[SDATA][56] , \spm_in[SDATA][55] , 
        \spm_in[SDATA][54] , \spm_in[SDATA][53] , \spm_in[SDATA][52] , 
        \spm_in[SDATA][51] , \spm_in[SDATA][50] , \spm_in[SDATA][49] , 
        \spm_in[SDATA][48] , \spm_in[SDATA][47] , \spm_in[SDATA][46] , 
        \spm_in[SDATA][45] , \spm_in[SDATA][44] , \spm_in[SDATA][43] , 
        \spm_in[SDATA][42] , \spm_in[SDATA][41] , \spm_in[SDATA][40] , 
        \spm_in[SDATA][39] , \spm_in[SDATA][38] , \spm_in[SDATA][37] , 
        \spm_in[SDATA][36] , \spm_in[SDATA][35] , \spm_in[SDATA][34] , 
        \spm_in[SDATA][33] , \spm_in[SDATA][32] , \spm_in[SDATA][31] , 
        \spm_in[SDATA][30] , \spm_in[SDATA][29] , \spm_in[SDATA][28] , 
        \spm_in[SDATA][27] , \spm_in[SDATA][26] , \spm_in[SDATA][25] , 
        \spm_in[SDATA][24] , \spm_in[SDATA][23] , \spm_in[SDATA][22] , 
        \spm_in[SDATA][21] , \spm_in[SDATA][20] , \spm_in[SDATA][19] , 
        \spm_in[SDATA][18] , \spm_in[SDATA][17] , \spm_in[SDATA][16] , 
        \spm_in[SDATA][15] , \spm_in[SDATA][14] , \spm_in[SDATA][13] , 
        \spm_in[SDATA][12] , \spm_in[SDATA][11] , \spm_in[SDATA][10] , 
        \spm_in[SDATA][9] , \spm_in[SDATA][8] , \spm_in[SDATA][7] , 
        \spm_in[SDATA][6] , \spm_in[SDATA][5] , \spm_in[SDATA][4] , 
        \spm_in[SDATA][3] , \spm_in[SDATA][2] , \spm_in[SDATA][1] , 
        \spm_in[SDATA][0] }), .spm_out({\spm_out[MCMD][1] , \spm_out[MCMD][0] , 
        \spm_out[MADDR][31] , \spm_out[MADDR][30] , \spm_out[MADDR][29] , 
        \spm_out[MADDR][28] , \spm_out[MADDR][27] , \spm_out[MADDR][26] , 
        \spm_out[MADDR][25] , \spm_out[MADDR][24] , \spm_out[MADDR][23] , 
        \spm_out[MADDR][22] , \spm_out[MADDR][21] , \spm_out[MADDR][20] , 
        \spm_out[MADDR][19] , \spm_out[MADDR][18] , \spm_out[MADDR][17] , 
        \spm_out[MADDR][16] , \spm_out[MADDR][15] , \spm_out[MADDR][14] , 
        \spm_out[MADDR][13] , \spm_out[MADDR][12] , \spm_out[MADDR][11] , 
        \spm_out[MADDR][10] , \spm_out[MADDR][9] , \spm_out[MADDR][8] , 
        \spm_out[MADDR][7] , \spm_out[MADDR][6] , \spm_out[MADDR][5] , 
        \spm_out[MADDR][4] , \spm_out[MADDR][3] , \spm_out[MADDR][2] , 
        \spm_out[MADDR][1] , \spm_out[MADDR][0] , \spm_out[MDATA][63] , 
        \spm_out[MDATA][62] , \spm_out[MDATA][61] , \spm_out[MDATA][60] , 
        \spm_out[MDATA][59] , \spm_out[MDATA][58] , \spm_out[MDATA][57] , 
        \spm_out[MDATA][56] , \spm_out[MDATA][55] , \spm_out[MDATA][54] , 
        \spm_out[MDATA][53] , \spm_out[MDATA][52] , \spm_out[MDATA][51] , 
        \spm_out[MDATA][50] , \spm_out[MDATA][49] , \spm_out[MDATA][48] , 
        \spm_out[MDATA][47] , \spm_out[MDATA][46] , \spm_out[MDATA][45] , 
        \spm_out[MDATA][44] , \spm_out[MDATA][43] , \spm_out[MDATA][42] , 
        \spm_out[MDATA][41] , \spm_out[MDATA][40] , \spm_out[MDATA][39] , 
        \spm_out[MDATA][38] , \spm_out[MDATA][37] , \spm_out[MDATA][36] , 
        \spm_out[MDATA][35] , \spm_out[MDATA][34] , \spm_out[MDATA][33] , 
        \spm_out[MDATA][32] , \spm_out[MDATA][31] , \spm_out[MDATA][30] , 
        \spm_out[MDATA][29] , \spm_out[MDATA][28] , \spm_out[MDATA][27] , 
        \spm_out[MDATA][26] , \spm_out[MDATA][25] , \spm_out[MDATA][24] , 
        \spm_out[MDATA][23] , \spm_out[MDATA][22] , \spm_out[MDATA][21] , 
        \spm_out[MDATA][20] , \spm_out[MDATA][19] , \spm_out[MDATA][18] , 
        \spm_out[MDATA][17] , \spm_out[MDATA][16] , \spm_out[MDATA][15] , 
        \spm_out[MDATA][14] , \spm_out[MDATA][13] , \spm_out[MDATA][12] , 
        \spm_out[MDATA][11] , \spm_out[MDATA][10] , \spm_out[MDATA][9] , 
        \spm_out[MDATA][8] , \spm_out[MDATA][7] , \spm_out[MDATA][6] , 
        \spm_out[MDATA][5] , \spm_out[MDATA][4] , \spm_out[MDATA][3] , 
        \spm_out[MDATA][2] , \spm_out[MDATA][1] , \spm_out[MDATA][0] }), 
        pkt_in, pkt_out );
  input [34:0] pkt_in;
  output [34:0] pkt_out;
  input na_clk, na_reset, \proc_in[MCMD][1] , \proc_in[MCMD][0] ,
         \proc_in[MADDR][31] , \proc_in[MADDR][30] , \proc_in[MADDR][29] ,
         \proc_in[MADDR][28] , \proc_in[MADDR][27] , \proc_in[MADDR][26] ,
         \proc_in[MADDR][25] , \proc_in[MADDR][24] , \proc_in[MADDR][23] ,
         \proc_in[MADDR][22] , \proc_in[MADDR][21] , \proc_in[MADDR][20] ,
         \proc_in[MADDR][19] , \proc_in[MADDR][18] , \proc_in[MADDR][17] ,
         \proc_in[MADDR][16] , \proc_in[MADDR][15] , \proc_in[MADDR][14] ,
         \proc_in[MADDR][13] , \proc_in[MADDR][12] , \proc_in[MADDR][11] ,
         \proc_in[MADDR][10] , \proc_in[MADDR][9] , \proc_in[MADDR][8] ,
         \proc_in[MADDR][7] , \proc_in[MADDR][6] , \proc_in[MADDR][5] ,
         \proc_in[MADDR][4] , \proc_in[MADDR][3] , \proc_in[MADDR][2] ,
         \proc_in[MADDR][1] , \proc_in[MADDR][0] , \proc_in[MDATA][31] ,
         \proc_in[MDATA][30] , \proc_in[MDATA][29] , \proc_in[MDATA][28] ,
         \proc_in[MDATA][27] , \proc_in[MDATA][26] , \proc_in[MDATA][25] ,
         \proc_in[MDATA][24] , \proc_in[MDATA][23] , \proc_in[MDATA][22] ,
         \proc_in[MDATA][21] , \proc_in[MDATA][20] , \proc_in[MDATA][19] ,
         \proc_in[MDATA][18] , \proc_in[MDATA][17] , \proc_in[MDATA][16] ,
         \proc_in[MDATA][15] , \proc_in[MDATA][14] , \proc_in[MDATA][13] ,
         \proc_in[MDATA][12] , \proc_in[MDATA][11] , \proc_in[MDATA][10] ,
         \proc_in[MDATA][9] , \proc_in[MDATA][8] , \proc_in[MDATA][7] ,
         \proc_in[MDATA][6] , \proc_in[MDATA][5] , \proc_in[MDATA][4] ,
         \proc_in[MDATA][3] , \proc_in[MDATA][2] , \proc_in[MDATA][1] ,
         \proc_in[MDATA][0] , \spm_in[SCMDACCEPT] , \spm_in[SRESP] ,
         \spm_in[SDATA][63] , \spm_in[SDATA][62] , \spm_in[SDATA][61] ,
         \spm_in[SDATA][60] , \spm_in[SDATA][59] , \spm_in[SDATA][58] ,
         \spm_in[SDATA][57] , \spm_in[SDATA][56] , \spm_in[SDATA][55] ,
         \spm_in[SDATA][54] , \spm_in[SDATA][53] , \spm_in[SDATA][52] ,
         \spm_in[SDATA][51] , \spm_in[SDATA][50] , \spm_in[SDATA][49] ,
         \spm_in[SDATA][48] , \spm_in[SDATA][47] , \spm_in[SDATA][46] ,
         \spm_in[SDATA][45] , \spm_in[SDATA][44] , \spm_in[SDATA][43] ,
         \spm_in[SDATA][42] , \spm_in[SDATA][41] , \spm_in[SDATA][40] ,
         \spm_in[SDATA][39] , \spm_in[SDATA][38] , \spm_in[SDATA][37] ,
         \spm_in[SDATA][36] , \spm_in[SDATA][35] , \spm_in[SDATA][34] ,
         \spm_in[SDATA][33] , \spm_in[SDATA][32] , \spm_in[SDATA][31] ,
         \spm_in[SDATA][30] , \spm_in[SDATA][29] , \spm_in[SDATA][28] ,
         \spm_in[SDATA][27] , \spm_in[SDATA][26] , \spm_in[SDATA][25] ,
         \spm_in[SDATA][24] , \spm_in[SDATA][23] , \spm_in[SDATA][22] ,
         \spm_in[SDATA][21] , \spm_in[SDATA][20] , \spm_in[SDATA][19] ,
         \spm_in[SDATA][18] , \spm_in[SDATA][17] , \spm_in[SDATA][16] ,
         \spm_in[SDATA][15] , \spm_in[SDATA][14] , \spm_in[SDATA][13] ,
         \spm_in[SDATA][12] , \spm_in[SDATA][11] , \spm_in[SDATA][10] ,
         \spm_in[SDATA][9] , \spm_in[SDATA][8] , \spm_in[SDATA][7] ,
         \spm_in[SDATA][6] , \spm_in[SDATA][5] , \spm_in[SDATA][4] ,
         \spm_in[SDATA][3] , \spm_in[SDATA][2] , \spm_in[SDATA][1] ,
         \spm_in[SDATA][0] ;
  output \proc_out[SCMDACCEPT] , \proc_out[SRESP] , \proc_out[SDATA][31] ,
         \proc_out[SDATA][30] , \proc_out[SDATA][29] , \proc_out[SDATA][28] ,
         \proc_out[SDATA][27] , \proc_out[SDATA][26] , \proc_out[SDATA][25] ,
         \proc_out[SDATA][24] , \proc_out[SDATA][23] , \proc_out[SDATA][22] ,
         \proc_out[SDATA][21] , \proc_out[SDATA][20] , \proc_out[SDATA][19] ,
         \proc_out[SDATA][18] , \proc_out[SDATA][17] , \proc_out[SDATA][16] ,
         \proc_out[SDATA][15] , \proc_out[SDATA][14] , \proc_out[SDATA][13] ,
         \proc_out[SDATA][12] , \proc_out[SDATA][11] , \proc_out[SDATA][10] ,
         \proc_out[SDATA][9] , \proc_out[SDATA][8] , \proc_out[SDATA][7] ,
         \proc_out[SDATA][6] , \proc_out[SDATA][5] , \proc_out[SDATA][4] ,
         \proc_out[SDATA][3] , \proc_out[SDATA][2] , \proc_out[SDATA][1] ,
         \proc_out[SDATA][0] , \spm_out[MCMD][1] , \spm_out[MCMD][0] ,
         \spm_out[MADDR][31] , \spm_out[MADDR][30] , \spm_out[MADDR][29] ,
         \spm_out[MADDR][28] , \spm_out[MADDR][27] , \spm_out[MADDR][26] ,
         \spm_out[MADDR][25] , \spm_out[MADDR][24] , \spm_out[MADDR][23] ,
         \spm_out[MADDR][22] , \spm_out[MADDR][21] , \spm_out[MADDR][20] ,
         \spm_out[MADDR][19] , \spm_out[MADDR][18] , \spm_out[MADDR][17] ,
         \spm_out[MADDR][16] , \spm_out[MADDR][15] , \spm_out[MADDR][14] ,
         \spm_out[MADDR][13] , \spm_out[MADDR][12] , \spm_out[MADDR][11] ,
         \spm_out[MADDR][10] , \spm_out[MADDR][9] , \spm_out[MADDR][8] ,
         \spm_out[MADDR][7] , \spm_out[MADDR][6] , \spm_out[MADDR][5] ,
         \spm_out[MADDR][4] , \spm_out[MADDR][3] , \spm_out[MADDR][2] ,
         \spm_out[MADDR][1] , \spm_out[MADDR][0] , \spm_out[MDATA][63] ,
         \spm_out[MDATA][62] , \spm_out[MDATA][61] , \spm_out[MDATA][60] ,
         \spm_out[MDATA][59] , \spm_out[MDATA][58] , \spm_out[MDATA][57] ,
         \spm_out[MDATA][56] , \spm_out[MDATA][55] , \spm_out[MDATA][54] ,
         \spm_out[MDATA][53] , \spm_out[MDATA][52] , \spm_out[MDATA][51] ,
         \spm_out[MDATA][50] , \spm_out[MDATA][49] , \spm_out[MDATA][48] ,
         \spm_out[MDATA][47] , \spm_out[MDATA][46] , \spm_out[MDATA][45] ,
         \spm_out[MDATA][44] , \spm_out[MDATA][43] , \spm_out[MDATA][42] ,
         \spm_out[MDATA][41] , \spm_out[MDATA][40] , \spm_out[MDATA][39] ,
         \spm_out[MDATA][38] , \spm_out[MDATA][37] , \spm_out[MDATA][36] ,
         \spm_out[MDATA][35] , \spm_out[MDATA][34] , \spm_out[MDATA][33] ,
         \spm_out[MDATA][32] , \spm_out[MDATA][31] , \spm_out[MDATA][30] ,
         \spm_out[MDATA][29] , \spm_out[MDATA][28] , \spm_out[MDATA][27] ,
         \spm_out[MDATA][26] , \spm_out[MDATA][25] , \spm_out[MDATA][24] ,
         \spm_out[MDATA][23] , \spm_out[MDATA][22] , \spm_out[MDATA][21] ,
         \spm_out[MDATA][20] , \spm_out[MDATA][19] , \spm_out[MDATA][18] ,
         \spm_out[MDATA][17] , \spm_out[MDATA][16] , \spm_out[MDATA][15] ,
         \spm_out[MDATA][14] , \spm_out[MDATA][13] , \spm_out[MDATA][12] ,
         \spm_out[MDATA][11] , \spm_out[MDATA][10] , \spm_out[MDATA][9] ,
         \spm_out[MDATA][8] , \spm_out[MDATA][7] , \spm_out[MDATA][6] ,
         \spm_out[MDATA][5] , \spm_out[MDATA][4] , \spm_out[MDATA][3] ,
         \spm_out[MDATA][2] , \spm_out[MDATA][1] , \spm_out[MDATA][0] ;
  wire   \spm_out[MCMD][0] , \phase_prev[0] , \phase_next[1] , vld_pkt,
         \add_545/A[8] , \add_545/A[9] , \add_545/A[10] , \add_545/A[11] ,
         \add_545/A[12] , \add_545/A[13] , \add_545/A[14] , \add_545/A[15] ,
         \sub_544/A[1] , \sub_544/A[2] , \sub_544/A[3] , \sub_544/A[4] ,
         \sub_544/A[5] , \sub_544/A[6] , \sub_544/A[7] , \sub_544/A[8] ,
         \sub_544/A[9] , \sub_544/A[10] , \sub_544/A[11] , \sub_544/A[12] , n1,
         n2, n3, n4, n5, n6, n15, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n34, n35, n37, n39, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n62, n64, n72, n73, n74, n75, n77, n78, n79, n80, n84, n87,
         n88, n89, n90, n91, n93, n94, n95, n101, n102, n103, n104, n105, n106,
         n108, n109, n111, n112, n113, n114, n116, n117, n118, n120, n122,
         n124, n125, n127, n128, n129, n130, n132, n133, n134, n136, n137,
         n138, n139, n140, n142, n144, n149, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n310, n311,
         n312, n313, n314, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878;
  wire   [2:0] slt_index;
  wire   [2:0] dma_ren;
  wire   [2:0] dma_wen;
  wire   [1:0] dma_waddr;
  wire   [63:0] dma_wdata;
  wire   [1:0] dma_raddr;
  wire   [63:0] dma_rdata;
  wire   [4:0] slt_entry;
  wire   [1:0] state_cnt;
  wire   [4:0] config_reg;
  wire   [70:64] flit_buf;
  wire   [34:0] phitIn;
  wire   [31:0] mux_out;
  wire   [31:0] dOut_l;
  wire   [34:32] phit_togo;
  wire   [34:0] phitOut0;
  wire   [34:0] phitOut1;
  wire   [34:0] phitOut2;
  wire   [13:0] dma_cnt_new;
  wire   [15:0] dma_rp_new;
  wire   [15:0] dma_wp_new;
  wire   [6:0] address;
  wire   [31:0] dIn_h;
  assign \spm_out[MADDR][15]  = 1'b0;
  assign \spm_out[MADDR][16]  = 1'b0;
  assign \spm_out[MADDR][17]  = 1'b0;
  assign \spm_out[MADDR][18]  = 1'b0;
  assign \spm_out[MADDR][19]  = 1'b0;
  assign \spm_out[MADDR][20]  = 1'b0;
  assign \spm_out[MADDR][21]  = 1'b0;
  assign \spm_out[MADDR][22]  = 1'b0;
  assign \spm_out[MADDR][23]  = 1'b0;
  assign \spm_out[MADDR][24]  = 1'b0;
  assign \spm_out[MADDR][25]  = 1'b0;
  assign \spm_out[MADDR][26]  = 1'b0;
  assign \spm_out[MADDR][27]  = 1'b0;
  assign \spm_out[MADDR][28]  = 1'b0;
  assign \spm_out[MADDR][29]  = 1'b0;
  assign \spm_out[MADDR][30]  = 1'b0;
  assign \spm_out[MADDR][31]  = 1'b0;
  assign \spm_out[MCMD][1]  = \spm_out[MCMD][0] ;

  HS65_LS_DFPRQX9 \phase_next_reg[1]  ( .D(n676), .CP(na_clk), .RN(n348), .Q(
        \phase_next[1] ) );
  HS65_LS_DFPRQX9 \dOut_l_reg[31]  ( .D(n686), .CP(na_clk), .RN(n352), .Q(
        dOut_l[31]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[30]  ( .D(n687), .CP(na_clk), .RN(n350), .Q(
        dOut_l[30]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[29]  ( .D(n688), .CP(na_clk), .RN(n348), .Q(
        dOut_l[29]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[28]  ( .D(n689), .CP(na_clk), .RN(n346), .Q(
        dOut_l[28]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[27]  ( .D(n690), .CP(na_clk), .RN(n351), .Q(
        dOut_l[27]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[26]  ( .D(n691), .CP(na_clk), .RN(n349), .Q(
        dOut_l[26]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[25]  ( .D(n692), .CP(na_clk), .RN(n354), .Q(
        dOut_l[25]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[24]  ( .D(n693), .CP(na_clk), .RN(n353), .Q(
        dOut_l[24]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[23]  ( .D(n694), .CP(na_clk), .RN(n341), .Q(
        dOut_l[23]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[22]  ( .D(n695), .CP(na_clk), .RN(n347), .Q(
        dOut_l[22]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[21]  ( .D(n696), .CP(na_clk), .RN(n346), .Q(
        dOut_l[21]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[20]  ( .D(n697), .CP(na_clk), .RN(n344), .Q(
        dOut_l[20]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[19]  ( .D(n698), .CP(na_clk), .RN(n343), .Q(
        dOut_l[19]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[18]  ( .D(n699), .CP(na_clk), .RN(n342), .Q(
        dOut_l[18]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[17]  ( .D(n700), .CP(na_clk), .RN(n344), .Q(
        dOut_l[17]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[16]  ( .D(n701), .CP(na_clk), .RN(n343), .Q(
        dOut_l[16]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[15]  ( .D(n702), .CP(na_clk), .RN(n342), .Q(
        dOut_l[15]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[14]  ( .D(n703), .CP(na_clk), .RN(n345), .Q(
        dOut_l[14]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[13]  ( .D(n704), .CP(na_clk), .RN(n355), .Q(
        dOut_l[13]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[12]  ( .D(n705), .CP(na_clk), .RN(n351), .Q(
        dOut_l[12]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[11]  ( .D(n706), .CP(na_clk), .RN(n349), .Q(
        dOut_l[11]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[10]  ( .D(n707), .CP(na_clk), .RN(n354), .Q(
        dOut_l[10]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[9]  ( .D(n708), .CP(na_clk), .RN(n353), .Q(
        dOut_l[9]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[8]  ( .D(n709), .CP(na_clk), .RN(n341), .Q(
        dOut_l[8]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[7]  ( .D(n710), .CP(na_clk), .RN(n347), .Q(
        dOut_l[7]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[6]  ( .D(n711), .CP(na_clk), .RN(n346), .Q(
        dOut_l[6]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[5]  ( .D(n712), .CP(na_clk), .RN(n344), .Q(
        dOut_l[5]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[4]  ( .D(n713), .CP(na_clk), .RN(n343), .Q(
        dOut_l[4]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[3]  ( .D(n714), .CP(na_clk), .RN(n342), .Q(
        dOut_l[3]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[2]  ( .D(n715), .CP(na_clk), .RN(n345), .Q(
        dOut_l[2]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[1]  ( .D(n716), .CP(na_clk), .RN(n355), .Q(
        dOut_l[1]) );
  HS65_LS_DFPRQX9 \dOut_l_reg[0]  ( .D(n717), .CP(na_clk), .RN(n348), .Q(
        dOut_l[0]) );
  HS65_LS_DFPRQX9 \phitIn_reg[34]  ( .D(pkt_in[34]), .CP(na_clk), .RN(n342), 
        .Q(phitIn[34]) );
  HS65_LS_DFPRQX9 \phitIn_reg[33]  ( .D(pkt_in[33]), .CP(na_clk), .RN(n343), 
        .Q(phitIn[33]) );
  HS65_LS_DFPRQX9 vld_pkt_reg ( .D(n679), .CP(na_clk), .RN(n344), .Q(vld_pkt)
         );
  HS65_LS_DFPRQX9 \phitIn_reg[32]  ( .D(pkt_in[32]), .CP(na_clk), .RN(n346), 
        .Q(phitIn[32]) );
  HS65_LS_DFPRQX9 \phitIn_reg[31]  ( .D(pkt_in[31]), .CP(na_clk), .RN(n347), 
        .Q(phitIn[31]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[31]  ( .D(n718), .CP(na_clk), .RN(n341), .Q(
        dIn_h[31]) );
  HS65_LS_DFPRQX9 \phitIn_reg[30]  ( .D(pkt_in[30]), .CP(na_clk), .RN(n353), 
        .Q(phitIn[30]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[30]  ( .D(n719), .CP(na_clk), .RN(n354), .Q(
        dIn_h[30]) );
  HS65_LS_DFPRQX9 \phitIn_reg[29]  ( .D(pkt_in[29]), .CP(na_clk), .RN(n349), 
        .Q(phitIn[29]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[29]  ( .D(n720), .CP(na_clk), .RN(n351), .Q(
        dIn_h[29]) );
  HS65_LS_DFPRQX9 \phitIn_reg[28]  ( .D(pkt_in[28]), .CP(na_clk), .RN(n350), 
        .Q(phitIn[28]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[28]  ( .D(n721), .CP(na_clk), .RN(n352), .Q(
        dIn_h[28]) );
  HS65_LS_DFPRQX9 \phitIn_reg[27]  ( .D(pkt_in[27]), .CP(na_clk), .RN(n350), 
        .Q(phitIn[27]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[27]  ( .D(n722), .CP(na_clk), .RN(n350), .Q(
        dIn_h[27]) );
  HS65_LS_DFPRQX9 \phitIn_reg[26]  ( .D(pkt_in[26]), .CP(na_clk), .RN(n350), 
        .Q(phitIn[26]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[26]  ( .D(n723), .CP(na_clk), .RN(n350), .Q(
        dIn_h[26]) );
  HS65_LS_DFPRQX9 \phitIn_reg[25]  ( .D(pkt_in[25]), .CP(na_clk), .RN(n350), 
        .Q(phitIn[25]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[25]  ( .D(n724), .CP(na_clk), .RN(n350), .Q(
        dIn_h[25]) );
  HS65_LS_DFPRQX9 \phitIn_reg[24]  ( .D(pkt_in[24]), .CP(na_clk), .RN(n350), 
        .Q(phitIn[24]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[24]  ( .D(n725), .CP(na_clk), .RN(n350), .Q(
        dIn_h[24]) );
  HS65_LS_DFPRQX9 \phitIn_reg[23]  ( .D(pkt_in[23]), .CP(na_clk), .RN(n350), 
        .Q(phitIn[23]) );
  HS65_LS_DFPRQX9 \address_reg[6]  ( .D(n726), .CP(na_clk), .RN(n350), .Q(
        address[6]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[23]  ( .D(n727), .CP(na_clk), .RN(n350), .Q(
        dIn_h[23]) );
  HS65_LS_DFPRQX9 \phitIn_reg[22]  ( .D(pkt_in[22]), .CP(na_clk), .RN(n350), 
        .Q(phitIn[22]) );
  HS65_LS_DFPRQX9 \address_reg[5]  ( .D(n728), .CP(na_clk), .RN(n350), .Q(
        address[5]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[22]  ( .D(n729), .CP(na_clk), .RN(n350), .Q(
        dIn_h[22]) );
  HS65_LS_DFPRQX9 \phitIn_reg[21]  ( .D(pkt_in[21]), .CP(na_clk), .RN(n350), 
        .Q(phitIn[21]) );
  HS65_LS_DFPRQX9 \address_reg[4]  ( .D(n730), .CP(na_clk), .RN(n351), .Q(
        address[4]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[21]  ( .D(n731), .CP(na_clk), .RN(n351), .Q(
        dIn_h[21]) );
  HS65_LS_DFPRQX9 \phitIn_reg[20]  ( .D(pkt_in[20]), .CP(na_clk), .RN(n351), 
        .Q(phitIn[20]) );
  HS65_LS_DFPRQX9 \address_reg[3]  ( .D(n732), .CP(na_clk), .RN(n351), .Q(
        address[3]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[20]  ( .D(n733), .CP(na_clk), .RN(n351), .Q(
        dIn_h[20]) );
  HS65_LS_DFPRQX9 \phitIn_reg[19]  ( .D(pkt_in[19]), .CP(na_clk), .RN(n351), 
        .Q(phitIn[19]) );
  HS65_LS_DFPRQX9 \address_reg[2]  ( .D(n734), .CP(na_clk), .RN(n351), .Q(
        address[2]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[19]  ( .D(n735), .CP(na_clk), .RN(n351), .Q(
        dIn_h[19]) );
  HS65_LS_DFPRQX9 \phitIn_reg[18]  ( .D(pkt_in[18]), .CP(na_clk), .RN(n351), 
        .Q(phitIn[18]) );
  HS65_LS_DFPRQX9 \address_reg[1]  ( .D(n736), .CP(na_clk), .RN(n351), .Q(
        address[1]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[18]  ( .D(n737), .CP(na_clk), .RN(n351), .Q(
        dIn_h[18]) );
  HS65_LS_DFPRQX9 \phitIn_reg[17]  ( .D(pkt_in[17]), .CP(na_clk), .RN(n351), 
        .Q(phitIn[17]) );
  HS65_LS_DFPRQX9 \address_reg[0]  ( .D(n738), .CP(na_clk), .RN(n351), .Q(
        address[0]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[17]  ( .D(n739), .CP(na_clk), .RN(n351), .Q(
        dIn_h[17]) );
  HS65_LS_DFPRQX9 \phitIn_reg[16]  ( .D(pkt_in[16]), .CP(na_clk), .RN(n352), 
        .Q(phitIn[16]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[16]  ( .D(n740), .CP(na_clk), .RN(n352), .Q(
        dIn_h[16]) );
  HS65_LS_DFPRQX9 \phitIn_reg[15]  ( .D(pkt_in[15]), .CP(na_clk), .RN(n352), 
        .Q(phitIn[15]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[15]  ( .D(n741), .CP(na_clk), .RN(n352), .Q(
        dIn_h[15]) );
  HS65_LS_DFPRQX9 \phitIn_reg[14]  ( .D(pkt_in[14]), .CP(na_clk), .RN(n352), 
        .Q(phitIn[14]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[14]  ( .D(n742), .CP(na_clk), .RN(n352), .Q(
        dIn_h[14]) );
  HS65_LS_DFPRQX9 \phitIn_reg[13]  ( .D(pkt_in[13]), .CP(na_clk), .RN(n352), 
        .Q(phitIn[13]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[13]  ( .D(n743), .CP(na_clk), .RN(n352), .Q(
        dIn_h[13]) );
  HS65_LS_DFPRQX9 \phitIn_reg[12]  ( .D(pkt_in[12]), .CP(na_clk), .RN(n352), 
        .Q(phitIn[12]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[12]  ( .D(n744), .CP(na_clk), .RN(n352), .Q(
        dIn_h[12]) );
  HS65_LS_DFPRQX9 \phitIn_reg[11]  ( .D(pkt_in[11]), .CP(na_clk), .RN(n352), 
        .Q(phitIn[11]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[11]  ( .D(n745), .CP(na_clk), .RN(n352), .Q(
        dIn_h[11]) );
  HS65_LS_DFPRQX9 \phitIn_reg[10]  ( .D(pkt_in[10]), .CP(na_clk), .RN(n352), 
        .Q(phitIn[10]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[10]  ( .D(n746), .CP(na_clk), .RN(n352), .Q(
        dIn_h[10]) );
  HS65_LS_DFPRQX9 \phitIn_reg[9]  ( .D(pkt_in[9]), .CP(na_clk), .RN(n352), .Q(
        phitIn[9]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[9]  ( .D(n747), .CP(na_clk), .RN(n353), .Q(
        dIn_h[9]) );
  HS65_LS_DFPRQX9 \phitIn_reg[8]  ( .D(pkt_in[8]), .CP(na_clk), .RN(n353), .Q(
        phitIn[8]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[8]  ( .D(n748), .CP(na_clk), .RN(n353), .Q(
        dIn_h[8]) );
  HS65_LS_DFPRQX9 \phitIn_reg[7]  ( .D(pkt_in[7]), .CP(na_clk), .RN(n353), .Q(
        phitIn[7]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[7]  ( .D(n749), .CP(na_clk), .RN(n353), .Q(
        dIn_h[7]) );
  HS65_LS_DFPRQX9 \phitIn_reg[6]  ( .D(pkt_in[6]), .CP(na_clk), .RN(n353), .Q(
        phitIn[6]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[6]  ( .D(n750), .CP(na_clk), .RN(n353), .Q(
        dIn_h[6]) );
  HS65_LS_DFPRQX9 \phitIn_reg[5]  ( .D(pkt_in[5]), .CP(na_clk), .RN(n353), .Q(
        phitIn[5]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[5]  ( .D(n751), .CP(na_clk), .RN(n353), .Q(
        dIn_h[5]) );
  HS65_LS_DFPRQX9 \phitIn_reg[4]  ( .D(pkt_in[4]), .CP(na_clk), .RN(n353), .Q(
        phitIn[4]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[4]  ( .D(n752), .CP(na_clk), .RN(n353), .Q(
        dIn_h[4]) );
  HS65_LS_DFPRQX9 \phitIn_reg[3]  ( .D(pkt_in[3]), .CP(na_clk), .RN(n353), .Q(
        phitIn[3]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[3]  ( .D(n753), .CP(na_clk), .RN(n353), .Q(
        dIn_h[3]) );
  HS65_LS_DFPRQX9 \phitIn_reg[2]  ( .D(pkt_in[2]), .CP(na_clk), .RN(n353), .Q(
        phitIn[2]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[2]  ( .D(n754), .CP(na_clk), .RN(n353), .Q(
        dIn_h[2]) );
  HS65_LS_DFPRQX9 \phitIn_reg[1]  ( .D(pkt_in[1]), .CP(na_clk), .RN(n354), .Q(
        phitIn[1]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[1]  ( .D(n755), .CP(na_clk), .RN(n354), .Q(
        dIn_h[1]) );
  HS65_LS_DFPRQX9 \phitIn_reg[0]  ( .D(pkt_in[0]), .CP(na_clk), .RN(n354), .Q(
        phitIn[0]) );
  HS65_LS_DFPRQX9 \dIn_h_reg[0]  ( .D(n756), .CP(na_clk), .RN(n354), .Q(
        dIn_h[0]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[34]  ( .D(phit_togo[34]), .CP(na_clk), .RN(
        n354), .Q(phitOut0[34]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[33]  ( .D(n333), .CP(na_clk), .RN(n354), .Q(
        phitOut0[33]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[32]  ( .D(phit_togo[32]), .CP(na_clk), .RN(
        n354), .Q(phitOut0[32]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[31]  ( .D(mux_out[31]), .CP(na_clk), .RN(n354), 
        .Q(phitOut0[31]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[30]  ( .D(mux_out[30]), .CP(na_clk), .RN(n354), 
        .Q(phitOut0[30]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[29]  ( .D(mux_out[29]), .CP(na_clk), .RN(n354), 
        .Q(phitOut0[29]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[28]  ( .D(mux_out[28]), .CP(na_clk), .RN(n354), 
        .Q(phitOut0[28]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[27]  ( .D(mux_out[27]), .CP(na_clk), .RN(n354), 
        .Q(phitOut0[27]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[26]  ( .D(mux_out[26]), .CP(na_clk), .RN(n354), 
        .Q(phitOut0[26]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[25]  ( .D(mux_out[25]), .CP(na_clk), .RN(n354), 
        .Q(phitOut0[25]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[24]  ( .D(mux_out[24]), .CP(na_clk), .RN(n354), 
        .Q(phitOut0[24]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[23]  ( .D(mux_out[23]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[23]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[22]  ( .D(mux_out[22]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[22]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[21]  ( .D(mux_out[21]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[21]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[20]  ( .D(mux_out[20]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[20]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[19]  ( .D(mux_out[19]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[19]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[18]  ( .D(mux_out[18]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[18]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[17]  ( .D(mux_out[17]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[17]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[16]  ( .D(mux_out[16]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[16]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[15]  ( .D(mux_out[15]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[15]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[14]  ( .D(mux_out[14]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[14]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[13]  ( .D(mux_out[13]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[13]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[12]  ( .D(mux_out[12]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[12]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[11]  ( .D(mux_out[11]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[11]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[10]  ( .D(mux_out[10]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[10]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[9]  ( .D(mux_out[9]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[9]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[8]  ( .D(mux_out[8]), .CP(na_clk), .RN(n355), 
        .Q(phitOut0[8]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[7]  ( .D(mux_out[7]), .CP(na_clk), .RN(n348), 
        .Q(phitOut0[7]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[6]  ( .D(mux_out[6]), .CP(na_clk), .RN(n345), 
        .Q(phitOut0[6]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[5]  ( .D(mux_out[5]), .CP(na_clk), .RN(n342), 
        .Q(phitOut0[5]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[4]  ( .D(mux_out[4]), .CP(na_clk), .RN(n343), 
        .Q(phitOut0[4]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[3]  ( .D(mux_out[3]), .CP(na_clk), .RN(n344), 
        .Q(phitOut0[3]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[2]  ( .D(mux_out[2]), .CP(na_clk), .RN(n346), 
        .Q(phitOut0[2]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[1]  ( .D(mux_out[1]), .CP(na_clk), .RN(n347), 
        .Q(phitOut0[1]) );
  HS65_LS_DFPRQX9 \phitOut0_reg[0]  ( .D(mux_out[0]), .CP(na_clk), .RN(n341), 
        .Q(phitOut0[0]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[34]  ( .D(phitOut0[34]), .CP(na_clk), .RN(n345), .Q(phitOut1[34]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[33]  ( .D(phitOut0[33]), .CP(na_clk), .RN(n341), .Q(phitOut1[33]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[32]  ( .D(phitOut0[32]), .CP(na_clk), .RN(n341), .Q(phitOut1[32]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[31]  ( .D(phitOut0[31]), .CP(na_clk), .RN(n341), .Q(phitOut1[31]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[30]  ( .D(phitOut0[30]), .CP(na_clk), .RN(n341), .Q(phitOut1[30]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[29]  ( .D(phitOut0[29]), .CP(na_clk), .RN(n341), .Q(phitOut1[29]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[28]  ( .D(phitOut0[28]), .CP(na_clk), .RN(n341), .Q(phitOut1[28]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[27]  ( .D(phitOut0[27]), .CP(na_clk), .RN(n341), .Q(phitOut1[27]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[26]  ( .D(phitOut0[26]), .CP(na_clk), .RN(n341), .Q(phitOut1[26]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[25]  ( .D(phitOut0[25]), .CP(na_clk), .RN(n341), .Q(phitOut1[25]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[24]  ( .D(phitOut0[24]), .CP(na_clk), .RN(n341), .Q(phitOut1[24]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[23]  ( .D(phitOut0[23]), .CP(na_clk), .RN(n341), .Q(phitOut1[23]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[22]  ( .D(phitOut0[22]), .CP(na_clk), .RN(n341), .Q(phitOut1[22]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[21]  ( .D(phitOut0[21]), .CP(na_clk), .RN(n355), .Q(phitOut1[21]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[20]  ( .D(phitOut0[20]), .CP(na_clk), .RN(n350), .Q(phitOut1[20]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[19]  ( .D(phitOut0[19]), .CP(na_clk), .RN(n352), .Q(phitOut1[19]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[18]  ( .D(phitOut0[18]), .CP(na_clk), .RN(n348), .Q(phitOut1[18]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[17]  ( .D(phitOut0[17]), .CP(na_clk), .RN(n341), .Q(phitOut1[17]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[16]  ( .D(phitOut0[16]), .CP(na_clk), .RN(n353), .Q(phitOut1[16]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[15]  ( .D(phitOut0[15]), .CP(na_clk), .RN(n354), .Q(phitOut1[15]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[14]  ( .D(phitOut0[14]), .CP(na_clk), .RN(n349), .Q(phitOut1[14]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[13]  ( .D(phitOut0[13]), .CP(na_clk), .RN(n345), .Q(phitOut1[13]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[12]  ( .D(phitOut0[12]), .CP(na_clk), .RN(n355), .Q(phitOut1[12]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[11]  ( .D(phitOut0[11]), .CP(na_clk), .RN(n351), .Q(phitOut1[11]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[10]  ( .D(phitOut0[10]), .CP(na_clk), .RN(n347), .Q(phitOut1[10]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[9]  ( .D(phitOut0[9]), .CP(na_clk), .RN(n345), 
        .Q(phitOut1[9]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[8]  ( .D(phitOut0[8]), .CP(na_clk), .RN(n350), 
        .Q(phitOut1[8]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[7]  ( .D(phitOut0[7]), .CP(na_clk), .RN(n352), 
        .Q(phitOut1[7]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[6]  ( .D(phitOut0[6]), .CP(na_clk), .RN(n342), 
        .Q(phitOut1[6]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[5]  ( .D(phitOut0[5]), .CP(na_clk), .RN(n342), 
        .Q(phitOut1[5]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[4]  ( .D(phitOut0[4]), .CP(na_clk), .RN(n342), 
        .Q(phitOut1[4]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[3]  ( .D(phitOut0[3]), .CP(na_clk), .RN(n342), 
        .Q(phitOut1[3]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[2]  ( .D(phitOut0[2]), .CP(na_clk), .RN(n342), 
        .Q(phitOut1[2]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[1]  ( .D(phitOut0[1]), .CP(na_clk), .RN(n342), 
        .Q(phitOut1[1]) );
  HS65_LS_DFPRQX9 \phitOut1_reg[0]  ( .D(phitOut0[0]), .CP(na_clk), .RN(n342), 
        .Q(phitOut1[0]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[34]  ( .D(phitOut1[34]), .CP(na_clk), .RN(n342), .Q(phitOut2[34]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[33]  ( .D(phitOut1[33]), .CP(na_clk), .RN(n342), .Q(phitOut2[33]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[32]  ( .D(phitOut1[32]), .CP(na_clk), .RN(n342), .Q(phitOut2[32]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[31]  ( .D(phitOut1[31]), .CP(na_clk), .RN(n342), .Q(phitOut2[31]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[30]  ( .D(phitOut1[30]), .CP(na_clk), .RN(n342), .Q(phitOut2[30]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[29]  ( .D(phitOut1[29]), .CP(na_clk), .RN(n342), .Q(phitOut2[29]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[28]  ( .D(phitOut1[28]), .CP(na_clk), .RN(n342), .Q(phitOut2[28]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[27]  ( .D(phitOut1[27]), .CP(na_clk), .RN(n342), .Q(phitOut2[27]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[26]  ( .D(phitOut1[26]), .CP(na_clk), .RN(n343), .Q(phitOut2[26]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[25]  ( .D(phitOut1[25]), .CP(na_clk), .RN(n343), .Q(phitOut2[25]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[24]  ( .D(phitOut1[24]), .CP(na_clk), .RN(n343), .Q(phitOut2[24]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[23]  ( .D(phitOut1[23]), .CP(na_clk), .RN(n343), .Q(phitOut2[23]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[22]  ( .D(phitOut1[22]), .CP(na_clk), .RN(n343), .Q(phitOut2[22]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[21]  ( .D(phitOut1[21]), .CP(na_clk), .RN(n343), .Q(phitOut2[21]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[20]  ( .D(phitOut1[20]), .CP(na_clk), .RN(n343), .Q(phitOut2[20]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[19]  ( .D(phitOut1[19]), .CP(na_clk), .RN(n343), .Q(phitOut2[19]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[18]  ( .D(phitOut1[18]), .CP(na_clk), .RN(n343), .Q(phitOut2[18]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[17]  ( .D(phitOut1[17]), .CP(na_clk), .RN(n343), .Q(phitOut2[17]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[16]  ( .D(phitOut1[16]), .CP(na_clk), .RN(n343), .Q(phitOut2[16]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[15]  ( .D(phitOut1[15]), .CP(na_clk), .RN(n343), .Q(phitOut2[15]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[14]  ( .D(phitOut1[14]), .CP(na_clk), .RN(n343), .Q(phitOut2[14]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[13]  ( .D(phitOut1[13]), .CP(na_clk), .RN(n343), .Q(phitOut2[13]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[12]  ( .D(phitOut1[12]), .CP(na_clk), .RN(n343), .Q(phitOut2[12]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[11]  ( .D(phitOut1[11]), .CP(na_clk), .RN(n344), .Q(phitOut2[11]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[10]  ( .D(phitOut1[10]), .CP(na_clk), .RN(n344), .Q(phitOut2[10]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[9]  ( .D(phitOut1[9]), .CP(na_clk), .RN(n344), 
        .Q(phitOut2[9]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[8]  ( .D(phitOut1[8]), .CP(na_clk), .RN(n344), 
        .Q(phitOut2[8]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[7]  ( .D(phitOut1[7]), .CP(na_clk), .RN(n344), 
        .Q(phitOut2[7]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[6]  ( .D(phitOut1[6]), .CP(na_clk), .RN(n344), 
        .Q(phitOut2[6]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[5]  ( .D(phitOut1[5]), .CP(na_clk), .RN(n344), 
        .Q(phitOut2[5]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[4]  ( .D(phitOut1[4]), .CP(na_clk), .RN(n344), 
        .Q(phitOut2[4]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[3]  ( .D(phitOut1[3]), .CP(na_clk), .RN(n344), 
        .Q(phitOut2[3]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[2]  ( .D(phitOut1[2]), .CP(na_clk), .RN(n344), 
        .Q(phitOut2[2]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[1]  ( .D(phitOut1[1]), .CP(na_clk), .RN(n344), 
        .Q(phitOut2[1]) );
  HS65_LS_DFPRQX9 \phitOut2_reg[0]  ( .D(phitOut1[0]), .CP(na_clk), .RN(n344), 
        .Q(phitOut2[0]) );
  HS65_LS_DFPRQX9 \config_reg_reg[4]  ( .D(\proc_in[MCMD][1] ), .CP(na_clk), 
        .RN(n344), .Q(config_reg[4]) );
  HS65_LS_DFPRQX9 \config_reg_reg[3]  ( .D(n675), .CP(na_clk), .RN(n344), .Q(
        config_reg[3]) );
  HS65_LS_DFPRQX9 \config_reg_reg[2]  ( .D(n652), .CP(na_clk), .RN(n344), .Q(
        config_reg[2]) );
  HS65_LS_DFPRQX9 \config_reg_reg[1]  ( .D(n653), .CP(na_clk), .RN(n345), .Q(
        config_reg[1]) );
  HS65_LS_DFPRQX9 \config_reg_reg[0]  ( .D(n651), .CP(na_clk), .RN(n345), .Q(
        config_reg[0]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[70]  ( .D(n757), .CP(na_clk), .RN(n345), .Q(
        flit_buf[70]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[69]  ( .D(n758), .CP(na_clk), .RN(n345), .Q(
        flit_buf[69]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[68]  ( .D(n759), .CP(na_clk), .RN(n345), .Q(
        flit_buf[68]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[67]  ( .D(n760), .CP(na_clk), .RN(n345), .Q(
        flit_buf[67]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[66]  ( .D(n761), .CP(na_clk), .RN(n345), .Q(
        flit_buf[66]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[65]  ( .D(n762), .CP(na_clk), .RN(n345), .Q(
        flit_buf[65]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[64]  ( .D(n763), .CP(na_clk), .RN(n345), .Q(
        flit_buf[64]) );
  HS65_LS_DFPRQX9 \flit_buf_reg[63]  ( .D(n764), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][63] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[62]  ( .D(n765), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][62] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[61]  ( .D(n766), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][61] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[60]  ( .D(n767), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][60] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[59]  ( .D(n768), .CP(na_clk), .RN(n345), .Q(
        \spm_out[MDATA][59] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[58]  ( .D(n769), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][58] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[57]  ( .D(n770), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][57] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[56]  ( .D(n771), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][56] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[55]  ( .D(n772), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][55] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[54]  ( .D(n773), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][54] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[53]  ( .D(n774), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][53] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[52]  ( .D(n775), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][52] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[51]  ( .D(n776), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][51] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[50]  ( .D(n777), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][50] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[49]  ( .D(n778), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][49] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[48]  ( .D(n779), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][48] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[47]  ( .D(n780), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][47] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[46]  ( .D(n781), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][46] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[45]  ( .D(n782), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][45] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[44]  ( .D(n783), .CP(na_clk), .RN(n346), .Q(
        \spm_out[MDATA][44] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[43]  ( .D(n784), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][43] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[42]  ( .D(n785), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][42] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[41]  ( .D(n786), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][41] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[40]  ( .D(n787), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][40] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[39]  ( .D(n788), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][39] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[38]  ( .D(n789), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][38] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[37]  ( .D(n790), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][37] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[36]  ( .D(n791), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][36] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[35]  ( .D(n792), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][35] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[34]  ( .D(n793), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][34] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[33]  ( .D(n794), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][33] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[32]  ( .D(n795), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][32] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[31]  ( .D(n796), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][31] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[30]  ( .D(n797), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][30] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[29]  ( .D(n798), .CP(na_clk), .RN(n347), .Q(
        \spm_out[MDATA][29] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[28]  ( .D(n799), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][28] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[27]  ( .D(n800), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][27] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[26]  ( .D(n801), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][26] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[25]  ( .D(n802), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][25] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[24]  ( .D(n803), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][24] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[23]  ( .D(n804), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][23] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[22]  ( .D(n805), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][22] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[21]  ( .D(n806), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][21] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[20]  ( .D(n807), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][20] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[19]  ( .D(n808), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][19] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[18]  ( .D(n809), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][18] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[17]  ( .D(n810), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][17] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[16]  ( .D(n811), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][16] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[15]  ( .D(n812), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][15] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[14]  ( .D(n813), .CP(na_clk), .RN(n348), .Q(
        \spm_out[MDATA][14] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[13]  ( .D(n814), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][13] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[12]  ( .D(n815), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][12] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[11]  ( .D(n816), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][11] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[10]  ( .D(n817), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][10] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[9]  ( .D(n818), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][9] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[8]  ( .D(n819), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][8] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[7]  ( .D(n820), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][7] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[6]  ( .D(n821), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][6] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[5]  ( .D(n822), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][5] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[4]  ( .D(n823), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][4] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[3]  ( .D(n824), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][3] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[2]  ( .D(n825), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][2] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[1]  ( .D(n826), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][1] ) );
  HS65_LS_DFPRQX9 \flit_buf_reg[0]  ( .D(n827), .CP(na_clk), .RN(n349), .Q(
        \spm_out[MDATA][0] ) );
  HS65_LS_DFPRQX9 \phase_prev_reg[0]  ( .D(n682), .CP(na_clk), .RN(n349), .Q(
        \phase_prev[0] ) );
  counter_WIDTH3_1 slt_cnt ( .clk(na_clk), .reset(n356), .enable(n647), .cnt(
        slt_index) );
  dma_sdp_DATA64_ADDR2_1 dma_table ( .clk(na_clk), .reset(n357), .ren(dma_ren), 
        .wen(dma_wen), .waddr(dma_waddr), .wdata(dma_wdata), .raddr(dma_raddr), 
        .rdata(dma_rdata) );
  bram_DATA5_ADDR3_1 slt_table ( .clk(na_clk), .reset(n356), .rd_addr(
        slt_index), .wr_addr({\proc_in[MADDR][2] , \proc_in[MADDR][1] , 
        \proc_in[MADDR][0] }), .wr_data({\proc_in[MDATA][4] , 
        \proc_in[MDATA][3] , \proc_in[MDATA][2] , \proc_in[MDATA][1] , 
        \proc_in[MDATA][0] }), .wr_ena(n650), .rd_data(slt_entry) );
  HS65_LS_DFPRQNX9 vld_buf_reg ( .D(n680), .CP(na_clk), .RN(n353), .QN(n683)
         );
  HS65_LS_DFPRQNX9 dma_ctrl_reg_reg ( .D(n678), .CP(na_clk), .RN(n354), .QN(
        n684) );
  HS65_LS_DFPRQX9 \state_cnt_reg[0]  ( .D(n142), .CP(na_clk), .RN(n341), .Q(
        state_cnt[0]) );
  HS65_LS_DFPRQX9 \state_cnt_reg[1]  ( .D(n597), .CP(na_clk), .RN(n351), .Q(
        state_cnt[1]) );
  HS65_LS_DFPRQNX4 \phase_next_reg[0]  ( .D(n677), .CP(na_clk), .RN(n349), 
        .QN(n685) );
  HS65_LS_DFPRQX9 \phase_prev_reg[1]  ( .D(n681), .CP(na_clk), .RN(n341), .Q(
        n21) );
  HS65_LH_IVX2 U3 ( .A(n18), .Z(n1) );
  HS65_LS_IVX4 U4 ( .A(n17), .Z(n18) );
  HS65_LS_IVX2 U5 ( .A(n35), .Z(n17) );
  HS65_LS_OAI212X5 U6 ( .A(n552), .B(n125), .C(n42), .D(n551), .E(n550), .Z(
        pkt_out[27]) );
  HS65_LS_IVX7 U7 ( .A(n458), .Z(n2) );
  HS65_LS_IVX9 U8 ( .A(n2), .Z(n3) );
  HS65_LS_NAND2X5 U9 ( .A(n20), .B(n448), .Z(n451) );
  HS65_LS_IVX31 U10 ( .A(n575), .Z(n122) );
  HS65_LS_IVX27 U11 ( .A(n122), .Z(n125) );
  HS65_LH_OAI222X2 U12 ( .A(n657), .B(n850), .C(n645), .D(n451), .E(n656), .F(
        n852), .Z(dma_waddr[1]) );
  HS65_LH_OAI222X2 U13 ( .A(n658), .B(n850), .C(n646), .D(n451), .E(n657), .F(
        n852), .Z(dma_waddr[0]) );
  HS65_LS_NAND2X4 U14 ( .A(n448), .B(n452), .Z(n449) );
  HS65_LS_AND2X4 U15 ( .A(\proc_in[MCMD][0] ), .B(n592), .Z(n4) );
  HS65_LS_AND2X4 U16 ( .A(n611), .B(n57), .Z(n5) );
  HS65_LS_AND2X4 U17 ( .A(\add_545/A[14] ), .B(n78), .Z(n6) );
  HS65_LS_AND2X4 U18 ( .A(n142), .B(n415), .Z(n15) );
  HS65_LS_NAND3X13 U19 ( .A(n127), .B(n455), .C(n454), .Z(n456) );
  HS65_LS_NAND2X14 U20 ( .A(n22), .B(n35), .Z(n39) );
  HS65_LS_OAI212X5 U21 ( .A(n571), .B(n125), .C(n42), .D(n569), .E(n568), .Z(
        pkt_out[33]) );
  HS65_LS_NAND2X2 U22 ( .A(phitOut2[10]), .B(n513), .Z(n498) );
  HS65_LS_NAND2X7 U23 ( .A(n27), .B(n111), .Z(n570) );
  HS65_LS_IVX9 U24 ( .A(n460), .Z(n463) );
  HS65_LS_CBI4I1X11 U25 ( .A(n3), .B(n112), .C(n457), .D(n456), .Z(n459) );
  HS65_LS_IVX2 U26 ( .A(n22), .Z(n19) );
  HS65_LS_IVX2 U27 ( .A(n452), .Z(n20) );
  HS65_LS_AND2X27 U28 ( .A(n27), .B(n572), .Z(n45) );
  HS65_LH_NAND2X2 U29 ( .A(n21), .B(n453), .Z(n460) );
  HS65_LS_IVX9 U30 ( .A(n21), .Z(n22) );
  HS65_LS_IVX18 U31 ( .A(n453), .Z(n35) );
  HS65_LS_BFX27 U32 ( .A(n113), .Z(n127) );
  HS65_LS_IVX27 U33 ( .A(n41), .Z(n31) );
  HS65_LS_IVX13 U34 ( .A(n25), .Z(n42) );
  HS65_LS_AND2X27 U35 ( .A(n118), .B(n30), .Z(n27) );
  HS65_LS_NAND2X4 U36 ( .A(phitOut2[26]), .B(n45), .Z(n547) );
  HS65_LS_IVX35 U37 ( .A(n25), .Z(n23) );
  HS65_LH_IVX2 U38 ( .A(n448), .Z(n24) );
  HS65_LS_IVX9 U39 ( .A(n25), .Z(n26) );
  HS65_LH_AND2X4 U40 ( .A(n24), .B(n415), .Z(phit_togo[32]) );
  HS65_LS_IVX18 U41 ( .A(n570), .Z(n25) );
  HS65_LS_NAND2X4 U42 ( .A(state_cnt[0]), .B(state_cnt[1]), .Z(n461) );
  HS65_LS_NAND2X4 U43 ( .A(n17), .B(n465), .Z(n450) );
  HS65_LS_NAND2X2 U44 ( .A(phitOut2[22]), .B(n44), .Z(n535) );
  HS65_LS_IVX18 U45 ( .A(n32), .Z(n34) );
  HS65_LS_NAND2X5 U46 ( .A(phitOut2[21]), .B(n45), .Z(n532) );
  HS65_LS_NAND2X5 U47 ( .A(phitOut2[23]), .B(n45), .Z(n538) );
  HS65_LS_NAND2X5 U48 ( .A(phitOut2[28]), .B(n45), .Z(n553) );
  HS65_LS_NAND2X5 U49 ( .A(phitOut2[18]), .B(n45), .Z(n523) );
  HS65_LS_NAND2X5 U50 ( .A(phitOut2[2]), .B(n45), .Z(n472) );
  HS65_LS_NAND2X5 U51 ( .A(phitOut2[16]), .B(n45), .Z(n517) );
  HS65_LS_NAND2X5 U52 ( .A(phitOut2[20]), .B(n45), .Z(n529) );
  HS65_LS_NAND2X5 U53 ( .A(phitOut2[24]), .B(n45), .Z(n541) );
  HS65_LS_NAND2X5 U54 ( .A(phitOut2[25]), .B(n45), .Z(n544) );
  HS65_LS_NAND2X5 U55 ( .A(phitOut2[31]), .B(n45), .Z(n562) );
  HS65_LS_NAND2X5 U56 ( .A(phitOut2[32]), .B(n45), .Z(n565) );
  HS65_LS_NAND2X5 U57 ( .A(phitOut2[29]), .B(n45), .Z(n556) );
  HS65_LS_IVX13 U58 ( .A(n122), .Z(n28) );
  HS65_LS_IVX13 U59 ( .A(n122), .Z(n29) );
  HS65_LS_CB4I1X18 U60 ( .A(n3), .B(n112), .C(n685), .D(n461), .Z(n30) );
  HS65_LS_NAND2X4 U61 ( .A(state_cnt[0]), .B(n37), .Z(n458) );
  HS65_LS_NAND2X14 U62 ( .A(n129), .B(n111), .Z(n575) );
  HS65_LS_NAND2X7 U63 ( .A(n118), .B(n30), .Z(n129) );
  HS65_LS_OAI21X6 U64 ( .A(n574), .B(n125), .C(n573), .Z(pkt_out[34]) );
  HS65_LS_IVX9 U65 ( .A(n117), .Z(n32) );
  HS65_LS_NAND2X2 U66 ( .A(phitOut2[7]), .B(n513), .Z(n489) );
  HS65_LS_NAND2X2 U67 ( .A(phitOut2[3]), .B(n513), .Z(n477) );
  HS65_LS_NAND2X2 U68 ( .A(phitOut2[11]), .B(n513), .Z(n501) );
  HS65_LS_OAI212X5 U69 ( .A(n500), .B(n43), .C(n23), .D(n499), .E(n498), .Z(
        pkt_out[10]) );
  HS65_LS_OAI212X5 U70 ( .A(n494), .B(n43), .C(n23), .D(n493), .E(n492), .Z(
        pkt_out[8]) );
  HS65_LS_AND2X18 U71 ( .A(n27), .B(n572), .Z(n44) );
  HS65_LS_NAND2X7 U72 ( .A(n27), .B(n572), .Z(n476) );
  HS65_LS_NAND2X14 U73 ( .A(n475), .B(n34), .Z(n572) );
  HS65_LS_IVX18 U74 ( .A(n459), .Z(n475) );
  HS65_LS_AND2X18 U75 ( .A(n475), .B(n34), .Z(n111) );
  HS65_LS_NAND2X7 U76 ( .A(n21), .B(n453), .Z(n37) );
  HS65_LS_NAND2X14 U77 ( .A(n37), .B(n39), .Z(n465) );
  HS65_LS_AOI312X4 U78 ( .A(n19), .B(n113), .C(n465), .D(n463), .E(n24), .F(
        n462), .Z(n117) );
  HS65_LS_AND2X18 U79 ( .A(n452), .B(n465), .Z(n112) );
  HS65_LS_AOI33X5 U80 ( .A(n464), .B(n465), .C(n18), .D(\phase_next[1] ), .E(
        n451), .F(n450), .Z(n118) );
  HS65_LS_IVX4 U81 ( .A(n465), .Z(n455) );
  HS65_LS_IVX9 U82 ( .A(n570), .Z(n41) );
  HS65_LS_IVX9 U83 ( .A(n122), .Z(n43) );
  HS65_LH_MUX21I1X3 U84 ( .D0(n22), .D1(\phase_next[1] ), .S0(n647), .Z(n681)
         );
  HS65_LS_NAND2X2 U85 ( .A(phitOut2[17]), .B(n44), .Z(n520) );
  HS65_LS_NAND2X2 U86 ( .A(phitOut2[19]), .B(n44), .Z(n526) );
  HS65_LS_NAND2X2 U87 ( .A(phitOut2[27]), .B(n44), .Z(n550) );
  HS65_LS_NAND2X2 U88 ( .A(phitOut2[30]), .B(n44), .Z(n559) );
  HS65_LS_OAI212X3 U89 ( .A(n561), .B(n125), .C(n42), .D(n560), .E(n559), .Z(
        pkt_out[30]) );
  HS65_LS_OAI212X3 U90 ( .A(n522), .B(n125), .C(n26), .D(n521), .E(n520), .Z(
        pkt_out[17]) );
  HS65_LS_OAI212X3 U91 ( .A(n528), .B(n125), .C(n26), .D(n527), .E(n526), .Z(
        pkt_out[19]) );
  HS65_LS_NAND2X4 U92 ( .A(phitOut2[33]), .B(n513), .Z(n568) );
  HS65_LS_OAI212X3 U93 ( .A(n537), .B(n125), .C(n42), .D(n536), .E(n535), .Z(
        pkt_out[22]) );
  HS65_LS_BFX9 U94 ( .A(n335), .Z(n331) );
  HS65_LS_BFX9 U95 ( .A(n335), .Z(n330) );
  HS65_LS_BFX9 U96 ( .A(n324), .Z(n310) );
  HS65_LS_BFX9 U97 ( .A(n324), .Z(n311) );
  HS65_LS_AND2X18 U98 ( .A(n448), .B(n452), .Z(n113) );
  HS65_LS_BFX9 U99 ( .A(n298), .Z(n301) );
  HS65_LS_BFX9 U100 ( .A(n340), .Z(n358) );
  HS65_LS_BFX9 U101 ( .A(n339), .Z(n357) );
  HS65_LS_BFX9 U102 ( .A(n339), .Z(n356) );
  HS65_LH_NAND2X2 U103 ( .A(n452), .B(n24), .Z(n365) );
  HS65_LH_MUXI21X2 U104 ( .D0(n457), .D1(n116), .S0(n647), .Z(n676) );
  HS65_LS_IVX9 U105 ( .A(n331), .Z(n325) );
  HS65_LS_IVX9 U106 ( .A(n331), .Z(n326) );
  HS65_LS_IVX9 U107 ( .A(n330), .Z(n327) );
  HS65_LS_IVX9 U108 ( .A(n330), .Z(n328) );
  HS65_LS_IVX9 U109 ( .A(n330), .Z(n329) );
  HS65_LS_AND2X4 U110 ( .A(n614), .B(n613), .Z(n46) );
  HS65_LS_AND2X4 U111 ( .A(n600), .B(n79), .Z(n47) );
  HS65_LS_AND2X4 U112 ( .A(n601), .B(n47), .Z(n48) );
  HS65_LS_AND2X4 U113 ( .A(n602), .B(n48), .Z(n49) );
  HS65_LS_AND2X4 U114 ( .A(n603), .B(n49), .Z(n50) );
  HS65_LS_AND2X4 U115 ( .A(n604), .B(n50), .Z(n51) );
  HS65_LS_AND2X4 U116 ( .A(n605), .B(n51), .Z(n52) );
  HS65_LS_AND2X4 U117 ( .A(n606), .B(n52), .Z(n53) );
  HS65_LS_AND2X4 U118 ( .A(n607), .B(n53), .Z(n54) );
  HS65_LS_AND2X4 U119 ( .A(n608), .B(n54), .Z(n55) );
  HS65_LS_AND2X4 U120 ( .A(n609), .B(n55), .Z(n56) );
  HS65_LS_AND2X4 U121 ( .A(n610), .B(n56), .Z(n57) );
  HS65_LS_AND2X4 U122 ( .A(n619), .B(n80), .Z(n58) );
  HS65_LS_AND2X4 U123 ( .A(n615), .B(n46), .Z(n59) );
  HS65_LS_AND2X4 U124 ( .A(n616), .B(n59), .Z(n62) );
  HS65_LS_AND2X4 U125 ( .A(n617), .B(n62), .Z(n64) );
  HS65_LS_AND2X4 U126 ( .A(\add_545/A[8] ), .B(n58), .Z(n72) );
  HS65_LS_AND2X4 U127 ( .A(\add_545/A[9] ), .B(n72), .Z(n73) );
  HS65_LS_AND2X4 U128 ( .A(\add_545/A[10] ), .B(n73), .Z(n74) );
  HS65_LS_AND2X4 U129 ( .A(\add_545/A[11] ), .B(n74), .Z(n75) );
  HS65_LS_AND2X4 U130 ( .A(\add_545/A[12] ), .B(n75), .Z(n77) );
  HS65_LS_AND2X4 U131 ( .A(\add_545/A[13] ), .B(n77), .Z(n78) );
  HS65_LS_AND2X4 U132 ( .A(n599), .B(n598), .Z(n79) );
  HS65_LS_AND2X4 U133 ( .A(n618), .B(n64), .Z(n80) );
  HS65_LS_BFX9 U134 ( .A(n334), .Z(n332) );
  HS65_LS_BFX9 U135 ( .A(n334), .Z(n333) );
  HS65_LS_IVX9 U136 ( .A(n310), .Z(n306) );
  HS65_LS_IVX9 U137 ( .A(n311), .Z(n305) );
  HS65_LS_IVX9 U138 ( .A(n311), .Z(n304) );
  HS65_LS_OAI21X3 U139 ( .A(n866), .B(n854), .C(n325), .Z(dma_wen[2]) );
  HS65_LS_NOR2AX3 U140 ( .A(n852), .B(n596), .Z(n866) );
  HS65_LS_IVX9 U141 ( .A(n850), .Z(n596) );
  HS65_LSS_XNOR2X6 U142 ( .A(n102), .B(\sub_544/A[10] ), .Z(dma_cnt_new[10])
         );
  HS65_LSS_XNOR2X6 U143 ( .A(n91), .B(\sub_544/A[5] ), .Z(dma_cnt_new[5]) );
  HS65_LSS_XNOR2X6 U144 ( .A(n101), .B(\sub_544/A[9] ), .Z(dma_cnt_new[9]) );
  HS65_LSS_XNOR2X6 U145 ( .A(n90), .B(\sub_544/A[4] ), .Z(dma_cnt_new[4]) );
  HS65_LSS_XNOR2X6 U146 ( .A(n95), .B(\sub_544/A[8] ), .Z(dma_cnt_new[8]) );
  HS65_LS_NOR4ABX2 U147 ( .A(n105), .B(n106), .C(n862), .D(dma_cnt_new[13]), 
        .Z(n844) );
  HS65_LSS_XOR2X6 U148 ( .A(n94), .B(\sub_544/A[7] ), .Z(n84) );
  HS65_LSS_XOR2X6 U149 ( .A(n89), .B(\sub_544/A[3] ), .Z(n87) );
  HS65_LSS_XOR2X6 U150 ( .A(n93), .B(\sub_544/A[6] ), .Z(n88) );
  HS65_LS_IVX9 U151 ( .A(n876), .Z(\add_545/A[8] ) );
  HS65_LS_IVX9 U152 ( .A(n877), .Z(\add_545/A[9] ) );
  HS65_LS_IVX9 U153 ( .A(n878), .Z(\add_545/A[10] ) );
  HS65_LS_IVX9 U154 ( .A(n871), .Z(\add_545/A[11] ) );
  HS65_LS_IVX9 U155 ( .A(n872), .Z(\add_545/A[12] ) );
  HS65_LS_IVX9 U156 ( .A(n873), .Z(\add_545/A[13] ) );
  HS65_LS_IVX9 U157 ( .A(n122), .Z(n124) );
  HS65_LS_BFX9 U158 ( .A(n109), .Z(n334) );
  HS65_LS_BFX9 U159 ( .A(n109), .Z(n335) );
  HS65_LS_OR2X9 U160 ( .A(\sub_544/A[2] ), .B(\sub_544/A[1] ), .Z(n89) );
  HS65_LS_OR2X9 U161 ( .A(\sub_544/A[3] ), .B(n89), .Z(n90) );
  HS65_LS_OR2X9 U162 ( .A(\sub_544/A[4] ), .B(n90), .Z(n91) );
  HS65_LS_OR2X9 U163 ( .A(\sub_544/A[5] ), .B(n91), .Z(n93) );
  HS65_LS_OR2X9 U164 ( .A(\sub_544/A[6] ), .B(n93), .Z(n94) );
  HS65_LS_OR2X9 U165 ( .A(\sub_544/A[7] ), .B(n94), .Z(n95) );
  HS65_LS_OR2X9 U166 ( .A(\sub_544/A[8] ), .B(n95), .Z(n101) );
  HS65_LS_OR2X9 U167 ( .A(\sub_544/A[9] ), .B(n101), .Z(n102) );
  HS65_LS_OR2X9 U168 ( .A(\sub_544/A[10] ), .B(n102), .Z(n103) );
  HS65_LS_OR2X9 U169 ( .A(\sub_544/A[11] ), .B(n103), .Z(n104) );
  HS65_LSS_XOR2X6 U170 ( .A(n103), .B(\sub_544/A[11] ), .Z(n105) );
  HS65_LSS_XOR2X6 U171 ( .A(n104), .B(\sub_544/A[12] ), .Z(n106) );
  HS65_LS_BFX9 U172 ( .A(n620), .Z(n144) );
  HS65_LS_BFX9 U173 ( .A(n620), .Z(n149) );
  HS65_LS_BFX9 U174 ( .A(n620), .Z(n293) );
  HS65_LS_IVX9 U175 ( .A(n874), .Z(\add_545/A[14] ) );
  HS65_LS_IVX9 U176 ( .A(n301), .Z(n299) );
  HS65_LS_IVX9 U177 ( .A(n301), .Z(n300) );
  HS65_LSS_XOR2X6 U178 ( .A(\sub_544/A[1] ), .B(\sub_544/A[2] ), .Z(n108) );
  HS65_LS_BFX9 U179 ( .A(n324), .Z(n312) );
  HS65_LS_BFX9 U180 ( .A(n324), .Z(n314) );
  HS65_LS_BFX9 U181 ( .A(n324), .Z(n313) );
  HS65_LS_BFX9 U182 ( .A(n294), .Z(n296) );
  HS65_LS_BFX9 U183 ( .A(n294), .Z(n295) );
  HS65_LS_BFX9 U184 ( .A(n324), .Z(n323) );
  HS65_LS_BFX9 U185 ( .A(n134), .Z(n136) );
  HS65_LS_BFX9 U186 ( .A(n134), .Z(n137) );
  HS65_LS_BFX9 U187 ( .A(n15), .Z(n130) );
  HS65_LS_BFX9 U188 ( .A(n15), .Z(n132) );
  HS65_LS_BFX9 U189 ( .A(n294), .Z(n297) );
  HS65_LS_BFX9 U190 ( .A(n134), .Z(n138) );
  HS65_LS_BFX9 U191 ( .A(n15), .Z(n133) );
  HS65_LS_IVX9 U192 ( .A(n854), .Z(n652) );
  HS65_LS_IVX9 U193 ( .A(\proc_out[SRESP] ), .Z(n336) );
  HS65_LS_IVX9 U194 ( .A(n358), .Z(n349) );
  HS65_LS_IVX9 U195 ( .A(n358), .Z(n348) );
  HS65_LS_IVX9 U196 ( .A(n358), .Z(n352) );
  HS65_LS_IVX9 U197 ( .A(n358), .Z(n350) );
  HS65_LS_IVX9 U198 ( .A(n358), .Z(n351) );
  HS65_LS_IVX9 U199 ( .A(n357), .Z(n347) );
  HS65_LS_IVX9 U200 ( .A(n357), .Z(n346) );
  HS65_LS_IVX9 U201 ( .A(n357), .Z(n344) );
  HS65_LS_IVX9 U202 ( .A(n357), .Z(n343) );
  HS65_LS_IVX9 U203 ( .A(n357), .Z(n342) );
  HS65_LS_IVX9 U204 ( .A(n357), .Z(n345) );
  HS65_LS_IVX9 U205 ( .A(n359), .Z(n355) );
  HS65_LS_IVX9 U206 ( .A(n359), .Z(n354) );
  HS65_LS_IVX9 U207 ( .A(n359), .Z(n353) );
  HS65_LS_IVX9 U208 ( .A(n356), .Z(n341) );
  HS65_LS_NOR2X6 U209 ( .A(n359), .B(n876), .Z(\spm_out[MADDR][7] ) );
  HS65_LS_NOR2X6 U210 ( .A(n359), .B(n877), .Z(\spm_out[MADDR][8] ) );
  HS65_LS_NOR2X6 U211 ( .A(n359), .B(n878), .Z(\spm_out[MADDR][9] ) );
  HS65_LS_NOR2X6 U212 ( .A(n359), .B(n871), .Z(\spm_out[MADDR][10] ) );
  HS65_LS_NOR2X6 U213 ( .A(n359), .B(n872), .Z(\spm_out[MADDR][11] ) );
  HS65_LS_NOR2X6 U214 ( .A(n359), .B(n873), .Z(\spm_out[MADDR][12] ) );
  HS65_LS_NOR2X6 U215 ( .A(n359), .B(n874), .Z(\spm_out[MADDR][13] ) );
  HS65_LS_NOR2X6 U216 ( .A(n359), .B(n875), .Z(\spm_out[MADDR][14] ) );
  HS65_LS_NOR2X6 U217 ( .A(n336), .B(n642), .Z(\proc_out[SDATA][0] ) );
  HS65_LS_NOR2X6 U218 ( .A(n336), .B(n641), .Z(\proc_out[SDATA][1] ) );
  HS65_LS_NOR2X6 U219 ( .A(n336), .B(n640), .Z(\proc_out[SDATA][2] ) );
  HS65_LS_NOR2X6 U220 ( .A(n870), .B(n639), .Z(\proc_out[SDATA][3] ) );
  HS65_LS_NOR2X6 U221 ( .A(n336), .B(n638), .Z(\proc_out[SDATA][4] ) );
  HS65_LS_NOR2X6 U222 ( .A(n870), .B(n637), .Z(\proc_out[SDATA][5] ) );
  HS65_LS_NOR2X6 U223 ( .A(n870), .B(n636), .Z(\proc_out[SDATA][6] ) );
  HS65_LS_NOR2X6 U224 ( .A(n870), .B(n635), .Z(\proc_out[SDATA][7] ) );
  HS65_LS_NOR2X6 U225 ( .A(n336), .B(n634), .Z(\proc_out[SDATA][8] ) );
  HS65_LS_NOR2X6 U226 ( .A(n336), .B(n633), .Z(\proc_out[SDATA][9] ) );
  HS65_LS_NOR2X6 U227 ( .A(n336), .B(n632), .Z(\proc_out[SDATA][10] ) );
  HS65_LS_NOR2X6 U228 ( .A(n336), .B(n631), .Z(\proc_out[SDATA][11] ) );
  HS65_LS_NOR2X6 U229 ( .A(n336), .B(n630), .Z(\proc_out[SDATA][12] ) );
  HS65_LS_NOR2X6 U230 ( .A(n336), .B(n629), .Z(\proc_out[SDATA][13] ) );
  HS65_LS_NOR2X6 U231 ( .A(n336), .B(n628), .Z(\proc_out[SDATA][14] ) );
  HS65_LS_NOR2X6 U232 ( .A(n336), .B(n627), .Z(\proc_out[SDATA][15] ) );
  HS65_LS_AND3X9 U233 ( .A(dma_rdata[63]), .B(n644), .C(n293), .Z(n109) );
  HS65_LS_OAI222X2 U234 ( .A(n331), .B(n836), .C(n849), .D(n674), .E(n325), 
        .F(n836), .Z(dma_wdata[48]) );
  HS65_LS_NOR2X6 U235 ( .A(n866), .B(n853), .Z(dma_wen[0]) );
  HS65_LS_OAI222X2 U236 ( .A(n331), .B(n837), .C(n849), .D(n671), .E(n325), 
        .F(n87), .Z(dma_wdata[51]) );
  HS65_LS_OAI222X2 U237 ( .A(n331), .B(n838), .C(n849), .D(n670), .E(n325), 
        .F(n626), .Z(dma_wdata[52]) );
  HS65_LS_IVX9 U238 ( .A(dma_cnt_new[4]), .Z(n626) );
  HS65_LS_OAI222X2 U239 ( .A(n331), .B(n839), .C(n667), .D(n849), .E(n325), 
        .F(n84), .Z(dma_wdata[55]) );
  HS65_LS_OAI222X2 U240 ( .A(n331), .B(n840), .C(n666), .D(n849), .E(n325), 
        .F(n624), .Z(dma_wdata[56]) );
  HS65_LS_IVX9 U241 ( .A(dma_cnt_new[8]), .Z(n624) );
  HS65_LS_OAI222X2 U242 ( .A(n331), .B(n841), .C(n849), .D(n664), .E(n326), 
        .F(n622), .Z(dma_wdata[58]) );
  HS65_LS_IVX9 U243 ( .A(dma_cnt_new[10]), .Z(n622) );
  HS65_LS_OAI222X2 U244 ( .A(n330), .B(n842), .C(n849), .D(n662), .E(n326), 
        .F(n106), .Z(dma_wdata[60]) );
  HS65_LS_OAI222X2 U245 ( .A(n331), .B(n843), .C(n849), .D(n661), .E(n325), 
        .F(n621), .Z(dma_wdata[61]) );
  HS65_LS_IVX9 U246 ( .A(dma_cnt_new[13]), .Z(n621) );
  HS65_LS_OAI222X2 U247 ( .A(n331), .B(n862), .C(n849), .D(n673), .E(n325), 
        .F(\sub_544/A[1] ), .Z(dma_wdata[49]) );
  HS65_LS_OAI222X2 U248 ( .A(n331), .B(n861), .C(n849), .D(n672), .E(n325), 
        .F(n108), .Z(dma_wdata[50]) );
  HS65_LS_OAI222X2 U249 ( .A(n331), .B(n860), .C(n849), .D(n669), .E(n325), 
        .F(n625), .Z(dma_wdata[53]) );
  HS65_LS_IVX9 U250 ( .A(dma_cnt_new[5]), .Z(n625) );
  HS65_LS_OAI222X2 U251 ( .A(n331), .B(n859), .C(n668), .D(n849), .E(n325), 
        .F(n88), .Z(dma_wdata[54]) );
  HS65_LS_OAI222X2 U252 ( .A(n331), .B(n858), .C(n665), .D(n849), .E(n325), 
        .F(n623), .Z(dma_wdata[57]) );
  HS65_LS_IVX9 U253 ( .A(dma_cnt_new[9]), .Z(n623) );
  HS65_LS_OAI222X2 U254 ( .A(n331), .B(n857), .C(n849), .D(n663), .E(n325), 
        .F(n105), .Z(dma_wdata[59]) );
  HS65_LS_OAI212X5 U255 ( .A(n849), .B(n660), .C(n851), .D(n644), .E(n848), 
        .Z(dma_wdata[62]) );
  HS65_LS_NAND4ABX3 U256 ( .A(n847), .B(n846), .C(n845), .D(n844), .Z(n848) );
  HS65_LS_NAND4ABX3 U257 ( .A(dma_cnt_new[5]), .B(dma_cnt_new[4]), .C(n108), 
        .D(n87), .Z(n846) );
  HS65_LS_NAND4ABX3 U258 ( .A(dma_cnt_new[9]), .B(dma_cnt_new[8]), .C(n88), 
        .D(n84), .Z(n847) );
  HS65_LS_NAND2X7 U259 ( .A(n651), .B(n4), .Z(n850) );
  HS65_LS_OAI21X3 U260 ( .A(n866), .B(n856), .C(n325), .Z(dma_wen[1]) );
  HS65_LS_NAND2X7 U261 ( .A(n365), .B(n128), .Z(n592) );
  HS65_LSS_XNOR2X6 U262 ( .A(n843), .B(n120), .Z(dma_cnt_new[13]) );
  HS65_LS_NOR2X6 U263 ( .A(\sub_544/A[12] ), .B(n104), .Z(n120) );
  HS65_LS_NOR3X4 U264 ( .A(n325), .B(dma_cnt_new[10]), .C(dma_cnt_new[0]), .Z(
        n845) );
  HS65_LS_IVX9 U265 ( .A(n836), .Z(dma_cnt_new[0]) );
  HS65_LS_IVX9 U266 ( .A(n862), .Z(\sub_544/A[1] ) );
  HS65_LS_NAND2X7 U267 ( .A(dma_rdata[40]), .B(n144), .Z(n876) );
  HS65_LS_NAND2X7 U268 ( .A(dma_rdata[41]), .B(n144), .Z(n877) );
  HS65_LS_NAND2X7 U269 ( .A(dma_rdata[42]), .B(n144), .Z(n878) );
  HS65_LS_NAND2X7 U270 ( .A(dma_rdata[43]), .B(n144), .Z(n871) );
  HS65_LS_NAND2X7 U271 ( .A(dma_rdata[44]), .B(n144), .Z(n872) );
  HS65_LS_NAND2X7 U272 ( .A(dma_rdata[45]), .B(n149), .Z(n873) );
  HS65_LS_IVX9 U273 ( .A(n837), .Z(\sub_544/A[3] ) );
  HS65_LS_IVX9 U274 ( .A(n838), .Z(\sub_544/A[4] ) );
  HS65_LS_IVX9 U275 ( .A(n839), .Z(\sub_544/A[7] ) );
  HS65_LS_IVX9 U276 ( .A(n840), .Z(\sub_544/A[8] ) );
  HS65_LS_IVX9 U277 ( .A(n841), .Z(\sub_544/A[10] ) );
  HS65_LS_IVX9 U278 ( .A(n861), .Z(\sub_544/A[2] ) );
  HS65_LS_IVX9 U279 ( .A(n860), .Z(\sub_544/A[5] ) );
  HS65_LS_IVX9 U280 ( .A(n859), .Z(\sub_544/A[6] ) );
  HS65_LS_IVX9 U281 ( .A(n858), .Z(\sub_544/A[9] ) );
  HS65_LS_IVX9 U282 ( .A(n857), .Z(\sub_544/A[11] ) );
  HS65_LS_OAI22X6 U283 ( .A(n851), .B(n643), .C(n849), .D(n659), .Z(
        dma_wdata[63]) );
  HS65_LS_IVX9 U284 ( .A(dma_rdata[63]), .Z(n643) );
  HS65_LS_OAI22X6 U285 ( .A(n851), .B(n642), .C(n850), .D(n674), .Z(
        dma_wdata[0]) );
  HS65_LS_OAI22X6 U286 ( .A(n851), .B(n641), .C(n850), .D(n673), .Z(
        dma_wdata[1]) );
  HS65_LS_OAI22X6 U287 ( .A(n851), .B(n640), .C(n850), .D(n672), .Z(
        dma_wdata[2]) );
  HS65_LS_OAI22X6 U288 ( .A(n851), .B(n639), .C(n850), .D(n671), .Z(
        dma_wdata[3]) );
  HS65_LS_OAI22X6 U289 ( .A(n851), .B(n638), .C(n850), .D(n670), .Z(
        dma_wdata[4]) );
  HS65_LS_OAI22X6 U290 ( .A(n851), .B(n637), .C(n850), .D(n669), .Z(
        dma_wdata[5]) );
  HS65_LS_OAI22X6 U291 ( .A(n851), .B(n636), .C(n850), .D(n668), .Z(
        dma_wdata[6]) );
  HS65_LS_OAI22X6 U292 ( .A(n851), .B(n635), .C(n850), .D(n667), .Z(
        dma_wdata[7]) );
  HS65_LS_OAI22X6 U293 ( .A(n851), .B(n634), .C(n850), .D(n666), .Z(
        dma_wdata[8]) );
  HS65_LS_OAI22X6 U294 ( .A(n851), .B(n633), .C(n850), .D(n665), .Z(
        dma_wdata[9]) );
  HS65_LS_OAI22X6 U295 ( .A(n851), .B(n632), .C(n850), .D(n664), .Z(
        dma_wdata[10]) );
  HS65_LS_OAI22X6 U296 ( .A(n851), .B(n631), .C(n850), .D(n663), .Z(
        dma_wdata[11]) );
  HS65_LS_OAI22X6 U297 ( .A(n851), .B(n630), .C(n850), .D(n662), .Z(
        dma_wdata[12]) );
  HS65_LS_OAI22X6 U298 ( .A(n851), .B(n629), .C(n850), .D(n661), .Z(
        dma_wdata[13]) );
  HS65_LS_OAI22X6 U299 ( .A(n851), .B(n628), .C(n850), .D(n660), .Z(
        dma_wdata[14]) );
  HS65_LS_OAI22X6 U300 ( .A(n851), .B(n627), .C(n850), .D(n659), .Z(
        dma_wdata[15]) );
  HS65_LS_OAI21X3 U301 ( .A(n651), .B(n834), .C(n361), .Z(n593) );
  HS65_LS_NAND2X7 U302 ( .A(n652), .B(n4), .Z(n849) );
  HS65_LS_IVX9 U303 ( .A(n863), .Z(n648) );
  HS65_LS_OAI21X3 U304 ( .A(n853), .B(n593), .C(n365), .Z(dma_ren[0]) );
  HS65_LH_OAI21X2 U305 ( .A(n856), .B(n593), .C(n365), .Z(dma_ren[1]) );
  HS65_LH_OAI21X2 U306 ( .A(n854), .B(n593), .C(n365), .Z(dma_ren[2]) );
  HS65_LS_NAND2X7 U307 ( .A(dma_rdata[46]), .B(n149), .Z(n874) );
  HS65_LS_NAND2X7 U308 ( .A(dma_rdata[47]), .B(n149), .Z(n875) );
  HS65_LS_IVX9 U309 ( .A(dma_rdata[0]), .Z(n642) );
  HS65_LS_IVX9 U310 ( .A(dma_rdata[1]), .Z(n641) );
  HS65_LS_IVX9 U311 ( .A(dma_rdata[2]), .Z(n640) );
  HS65_LS_IVX9 U312 ( .A(dma_rdata[3]), .Z(n639) );
  HS65_LS_IVX9 U313 ( .A(dma_rdata[4]), .Z(n638) );
  HS65_LS_IVX9 U314 ( .A(dma_rdata[5]), .Z(n637) );
  HS65_LS_IVX9 U315 ( .A(dma_rdata[6]), .Z(n636) );
  HS65_LS_IVX9 U316 ( .A(dma_rdata[7]), .Z(n635) );
  HS65_LS_IVX9 U317 ( .A(dma_rdata[8]), .Z(n634) );
  HS65_LS_IVX9 U318 ( .A(dma_rdata[9]), .Z(n633) );
  HS65_LS_IVX9 U319 ( .A(dma_rdata[10]), .Z(n632) );
  HS65_LS_IVX9 U320 ( .A(dma_rdata[11]), .Z(n631) );
  HS65_LS_IVX9 U321 ( .A(dma_rdata[12]), .Z(n630) );
  HS65_LS_IVX9 U322 ( .A(dma_rdata[13]), .Z(n629) );
  HS65_LS_IVX9 U323 ( .A(dma_rdata[14]), .Z(n628) );
  HS65_LS_IVX9 U324 ( .A(dma_rdata[15]), .Z(n627) );
  HS65_LS_IVX9 U325 ( .A(n842), .Z(\sub_544/A[12] ) );
  HS65_LS_BFX9 U326 ( .A(n414), .Z(n134) );
  HS65_LS_BFX9 U327 ( .A(n835), .Z(n294) );
  HS65_LS_NOR2AX3 U328 ( .A(n4), .B(n856), .Z(n835) );
  HS65_LS_BFX9 U329 ( .A(n298), .Z(n302) );
  HS65_LS_IVX9 U330 ( .A(n865), .Z(n324) );
  HS65_LS_BFX9 U331 ( .A(n298), .Z(n303) );
  HS65_LS_NAND3X5 U332 ( .A(n142), .B(n576), .C(n341), .Z(n591) );
  HS65_LS_IVX9 U333 ( .A(n853), .Z(n651) );
  HS65_LS_NAND2X7 U334 ( .A(n854), .B(n856), .Z(n834) );
  HS65_LS_NAND2X7 U335 ( .A(n831), .B(n658), .Z(n854) );
  HS65_LS_BFX9 U336 ( .A(n338), .Z(\proc_out[SRESP] ) );
  HS65_LS_IVX9 U337 ( .A(n870), .Z(n338) );
  HS65_LS_BFX9 U338 ( .A(n340), .Z(n359) );
  HS65_LS_IVX9 U339 ( .A(n867), .Z(n650) );
  HS65_LS_NOR2AX3 U340 ( .A(dma_rdata[16]), .B(n870), .Z(\proc_out[SDATA][16] ) );
  HS65_LS_NOR2AX3 U341 ( .A(dma_rdata[17]), .B(n870), .Z(\proc_out[SDATA][17] ) );
  HS65_LS_NOR2AX3 U342 ( .A(dma_rdata[18]), .B(n870), .Z(\proc_out[SDATA][18] ) );
  HS65_LS_NOR2AX3 U343 ( .A(dma_rdata[19]), .B(n870), .Z(\proc_out[SDATA][19] ) );
  HS65_LS_NOR2AX3 U344 ( .A(dma_rdata[20]), .B(n870), .Z(\proc_out[SDATA][20] ) );
  HS65_LS_NOR2AX3 U345 ( .A(dma_rdata[21]), .B(n870), .Z(\proc_out[SDATA][21] ) );
  HS65_LS_NOR2AX3 U346 ( .A(dma_rdata[22]), .B(n870), .Z(\proc_out[SDATA][22] ) );
  HS65_LS_NOR2AX3 U347 ( .A(dma_rdata[23]), .B(n870), .Z(\proc_out[SDATA][23] ) );
  HS65_LS_NOR2AX3 U348 ( .A(dma_rdata[24]), .B(n870), .Z(\proc_out[SDATA][24] ) );
  HS65_LS_NOR2AX3 U349 ( .A(dma_rdata[25]), .B(n870), .Z(\proc_out[SDATA][25] ) );
  HS65_LS_NOR2AX3 U350 ( .A(dma_rdata[26]), .B(n336), .Z(\proc_out[SDATA][26] ) );
  HS65_LS_NOR2AX3 U351 ( .A(dma_rdata[27]), .B(n870), .Z(\proc_out[SDATA][27] ) );
  HS65_LS_NOR2AX3 U352 ( .A(dma_rdata[28]), .B(n870), .Z(\proc_out[SDATA][28] ) );
  HS65_LS_NOR2AX3 U353 ( .A(dma_rdata[29]), .B(n336), .Z(\proc_out[SDATA][29] ) );
  HS65_LS_NOR2AX3 U354 ( .A(dma_rdata[30]), .B(n870), .Z(\proc_out[SDATA][30] ) );
  HS65_LS_NOR2AX3 U355 ( .A(dma_rdata[31]), .B(n870), .Z(\proc_out[SDATA][31] ) );
  HS65_LS_IVX9 U356 ( .A(n856), .Z(n653) );
  HS65_LS_AOI22X6 U357 ( .A(\proc_in[MADDR][1] ), .B(n651), .C(
        \proc_in[MADDR][2] ), .D(n834), .Z(n833) );
  HS65_LS_IVX9 U358 ( .A(\proc_in[MADDR][2] ), .Z(n656) );
  HS65_LS_NAND2X7 U359 ( .A(slt_entry[4]), .B(n647), .Z(n851) );
  HS65_LH_MUXI21X2 U360 ( .D0(n685), .D1(n114), .S0(n647), .Z(n677) );
  HS65_LS_NOR2X6 U361 ( .A(slt_entry[0]), .B(n327), .Z(n114) );
  HS65_LS_NOR2X6 U362 ( .A(slt_entry[1]), .B(n327), .Z(n116) );
  HS65_LS_OAI21X3 U363 ( .A(n684), .B(n647), .C(n327), .Z(n678) );
  HS65_LS_MX41X7 U364 ( .D0(n595), .S0(n332), .D1(n595), .S1(n326), .D2(
        \proc_in[MDATA][16] ), .S2(n596), .D3(n295), .S3(\proc_in[MDATA][0] ), 
        .Z(dma_wdata[16]) );
  HS65_LS_MX41X7 U365 ( .D0(n385), .S0(n331), .D1(n598), .S1(n326), .D2(
        \proc_in[MDATA][17] ), .S2(n596), .D3(n295), .S3(\proc_in[MDATA][1] ), 
        .Z(dma_wdata[17]) );
  HS65_LS_MX41X7 U366 ( .D0(dma_wp_new[2]), .S0(n331), .D1(n599), .S1(n326), 
        .D2(\proc_in[MDATA][18] ), .S2(n596), .D3(n295), .S3(
        \proc_in[MDATA][2] ), .Z(dma_wdata[18]) );
  HS65_LSS_XOR2X6 U367 ( .A(n598), .B(n599), .Z(dma_wp_new[2]) );
  HS65_LS_MX41X7 U368 ( .D0(dma_wp_new[3]), .S0(n331), .D1(n600), .S1(n326), 
        .D2(\proc_in[MDATA][19] ), .S2(n596), .D3(n295), .S3(
        \proc_in[MDATA][3] ), .Z(dma_wdata[19]) );
  HS65_LSS_XOR2X6 U369 ( .A(n79), .B(n600), .Z(dma_wp_new[3]) );
  HS65_LS_MX41X7 U370 ( .D0(dma_wp_new[4]), .S0(n331), .D1(n601), .S1(n326), 
        .D2(\proc_in[MDATA][20] ), .S2(n596), .D3(n295), .S3(
        \proc_in[MDATA][4] ), .Z(dma_wdata[20]) );
  HS65_LSS_XOR2X6 U371 ( .A(n47), .B(n601), .Z(dma_wp_new[4]) );
  HS65_LS_MX41X7 U372 ( .D0(dma_wp_new[5]), .S0(n331), .D1(n602), .S1(n326), 
        .D2(\proc_in[MDATA][21] ), .S2(n596), .D3(n295), .S3(
        \proc_in[MDATA][5] ), .Z(dma_wdata[21]) );
  HS65_LSS_XOR2X6 U373 ( .A(n48), .B(n602), .Z(dma_wp_new[5]) );
  HS65_LS_MX41X7 U374 ( .D0(dma_wp_new[6]), .S0(n332), .D1(n603), .S1(n326), 
        .D2(\proc_in[MDATA][22] ), .S2(n596), .D3(n295), .S3(
        \proc_in[MDATA][6] ), .Z(dma_wdata[22]) );
  HS65_LSS_XOR2X6 U375 ( .A(n49), .B(n603), .Z(dma_wp_new[6]) );
  HS65_LS_MX41X7 U376 ( .D0(dma_wp_new[7]), .S0(n332), .D1(n604), .S1(n326), 
        .D2(\proc_in[MDATA][23] ), .S2(n596), .D3(n295), .S3(
        \proc_in[MDATA][7] ), .Z(dma_wdata[23]) );
  HS65_LSS_XOR2X6 U377 ( .A(n50), .B(n604), .Z(dma_wp_new[7]) );
  HS65_LS_MX41X7 U378 ( .D0(dma_wp_new[8]), .S0(n332), .D1(n605), .S1(n326), 
        .D2(\proc_in[MDATA][24] ), .S2(n596), .D3(n295), .S3(
        \proc_in[MDATA][8] ), .Z(dma_wdata[24]) );
  HS65_LSS_XOR2X6 U379 ( .A(n51), .B(n605), .Z(dma_wp_new[8]) );
  HS65_LS_MX41X7 U380 ( .D0(dma_wp_new[9]), .S0(n332), .D1(n606), .S1(n326), 
        .D2(\proc_in[MDATA][25] ), .S2(n596), .D3(n295), .S3(
        \proc_in[MDATA][9] ), .Z(dma_wdata[25]) );
  HS65_LSS_XOR2X6 U381 ( .A(n52), .B(n606), .Z(dma_wp_new[9]) );
  HS65_LS_MX41X7 U382 ( .D0(dma_wp_new[10]), .S0(n332), .D1(n607), .S1(n326), 
        .D2(\proc_in[MDATA][26] ), .S2(n596), .D3(n295), .S3(
        \proc_in[MDATA][10] ), .Z(dma_wdata[26]) );
  HS65_LSS_XOR2X6 U383 ( .A(n53), .B(n607), .Z(dma_wp_new[10]) );
  HS65_LS_MX41X7 U384 ( .D0(dma_wp_new[11]), .S0(n332), .D1(n608), .S1(n326), 
        .D2(\proc_in[MDATA][27] ), .S2(n596), .D3(n295), .S3(
        \proc_in[MDATA][11] ), .Z(dma_wdata[27]) );
  HS65_LSS_XOR2X6 U385 ( .A(n54), .B(n608), .Z(dma_wp_new[11]) );
  HS65_LS_MX41X7 U386 ( .D0(dma_wp_new[12]), .S0(n332), .D1(n609), .S1(n326), 
        .D2(\proc_in[MDATA][28] ), .S2(n596), .D3(n296), .S3(
        \proc_in[MDATA][12] ), .Z(dma_wdata[28]) );
  HS65_LSS_XOR2X6 U387 ( .A(n55), .B(n609), .Z(dma_wp_new[12]) );
  HS65_LS_MX41X7 U388 ( .D0(dma_wp_new[13]), .S0(n332), .D1(n610), .S1(n326), 
        .D2(\proc_in[MDATA][29] ), .S2(n596), .D3(n296), .S3(
        \proc_in[MDATA][13] ), .Z(dma_wdata[29]) );
  HS65_LSS_XOR2X6 U389 ( .A(n56), .B(n610), .Z(dma_wp_new[13]) );
  HS65_LS_MX41X7 U390 ( .D0(dma_wp_new[14]), .S0(n332), .D1(n611), .S1(n326), 
        .D2(\proc_in[MDATA][30] ), .S2(n596), .D3(n296), .S3(
        \proc_in[MDATA][14] ), .Z(dma_wdata[30]) );
  HS65_LSS_XOR2X6 U391 ( .A(n57), .B(n611), .Z(dma_wp_new[14]) );
  HS65_LS_MX41X7 U392 ( .D0(dma_wp_new[15]), .S0(n332), .D1(n612), .S1(n326), 
        .D2(\proc_in[MDATA][31] ), .S2(n596), .D3(n296), .S3(
        \proc_in[MDATA][15] ), .Z(dma_wdata[31]) );
  HS65_LSS_XOR2X6 U393 ( .A(n612), .B(n5), .Z(dma_wp_new[15]) );
  HS65_LS_AO222X4 U394 ( .A(n613), .B(n327), .C(\proc_in[MDATA][17] ), .D(n296), .E(n578), .F(n332), .Z(dma_wdata[33]) );
  HS65_LS_AO222X4 U395 ( .A(n614), .B(n327), .C(\proc_in[MDATA][18] ), .D(n296), .E(dma_rp_new[2]), .F(n332), .Z(dma_wdata[34]) );
  HS65_LSS_XOR2X6 U396 ( .A(n613), .B(n614), .Z(dma_rp_new[2]) );
  HS65_LS_AO222X4 U397 ( .A(n615), .B(n327), .C(\proc_in[MDATA][19] ), .D(n296), .E(dma_rp_new[3]), .F(n332), .Z(dma_wdata[35]) );
  HS65_LSS_XOR2X6 U398 ( .A(n46), .B(n615), .Z(dma_rp_new[3]) );
  HS65_LS_AO222X4 U399 ( .A(n616), .B(n326), .C(\proc_in[MDATA][20] ), .D(n296), .E(dma_rp_new[4]), .F(n332), .Z(dma_wdata[36]) );
  HS65_LSS_XOR2X6 U400 ( .A(n59), .B(n616), .Z(dma_rp_new[4]) );
  HS65_LS_AO222X4 U401 ( .A(n617), .B(n327), .C(\proc_in[MDATA][21] ), .D(n296), .E(dma_rp_new[5]), .F(n332), .Z(dma_wdata[37]) );
  HS65_LSS_XOR2X6 U402 ( .A(n62), .B(n617), .Z(dma_rp_new[5]) );
  HS65_LS_AO222X4 U403 ( .A(n618), .B(n327), .C(\proc_in[MDATA][22] ), .D(n296), .E(dma_rp_new[6]), .F(n332), .Z(dma_wdata[38]) );
  HS65_LSS_XOR2X6 U404 ( .A(n64), .B(n618), .Z(dma_rp_new[6]) );
  HS65_LS_AO222X4 U405 ( .A(n619), .B(n327), .C(\proc_in[MDATA][23] ), .D(n296), .E(dma_rp_new[7]), .F(n332), .Z(dma_wdata[39]) );
  HS65_LSS_XOR2X6 U406 ( .A(n80), .B(n619), .Z(dma_rp_new[7]) );
  HS65_LS_AO222X4 U407 ( .A(\add_545/A[8] ), .B(n327), .C(\proc_in[MDATA][24] ), .D(n296), .E(dma_rp_new[8]), .F(n332), .Z(dma_wdata[40]) );
  HS65_LSS_XOR2X6 U408 ( .A(n58), .B(\add_545/A[8] ), .Z(dma_rp_new[8]) );
  HS65_LS_AO222X4 U409 ( .A(\add_545/A[9] ), .B(n327), .C(\proc_in[MDATA][25] ), .D(n297), .E(dma_rp_new[9]), .F(n333), .Z(dma_wdata[41]) );
  HS65_LSS_XOR2X6 U410 ( .A(n72), .B(\add_545/A[9] ), .Z(dma_rp_new[9]) );
  HS65_LS_AO222X4 U411 ( .A(\add_545/A[10] ), .B(n327), .C(
        \proc_in[MDATA][26] ), .D(n297), .E(dma_rp_new[10]), .F(n333), .Z(
        dma_wdata[42]) );
  HS65_LSS_XOR2X6 U412 ( .A(n73), .B(\add_545/A[10] ), .Z(dma_rp_new[10]) );
  HS65_LS_AO222X4 U413 ( .A(\add_545/A[11] ), .B(n327), .C(
        \proc_in[MDATA][27] ), .D(n297), .E(dma_rp_new[11]), .F(n333), .Z(
        dma_wdata[43]) );
  HS65_LSS_XOR2X6 U414 ( .A(n74), .B(\add_545/A[11] ), .Z(dma_rp_new[11]) );
  HS65_LS_AO222X4 U415 ( .A(\add_545/A[12] ), .B(n327), .C(
        \proc_in[MDATA][28] ), .D(n297), .E(dma_rp_new[12]), .F(n333), .Z(
        dma_wdata[44]) );
  HS65_LSS_XOR2X6 U416 ( .A(n75), .B(\add_545/A[12] ), .Z(dma_rp_new[12]) );
  HS65_LS_AO222X4 U417 ( .A(\add_545/A[13] ), .B(n327), .C(
        \proc_in[MDATA][29] ), .D(n297), .E(dma_rp_new[13]), .F(n333), .Z(
        dma_wdata[45]) );
  HS65_LSS_XOR2X6 U418 ( .A(n77), .B(\add_545/A[13] ), .Z(dma_rp_new[13]) );
  HS65_LS_AO222X4 U419 ( .A(\add_545/A[14] ), .B(n326), .C(
        \proc_in[MDATA][30] ), .D(n297), .E(dma_rp_new[14]), .F(n333), .Z(
        dma_wdata[46]) );
  HS65_LSS_XOR2X6 U420 ( .A(n78), .B(\add_545/A[14] ), .Z(dma_rp_new[14]) );
  HS65_LS_AO222X4 U421 ( .A(dma_rp_new[0]), .B(n327), .C(\proc_in[MDATA][16] ), 
        .D(n296), .E(dma_rp_new[0]), .F(n332), .Z(dma_wdata[32]) );
  HS65_LS_NOR2AX3 U422 ( .A(dma_rdata[32]), .B(n851), .Z(dma_rp_new[0]) );
  HS65_LS_AO222X4 U423 ( .A(\add_545/A[15] ), .B(n327), .C(
        \proc_in[MDATA][31] ), .D(n297), .E(dma_rp_new[15]), .F(n333), .Z(
        dma_wdata[47]) );
  HS65_LSS_XOR2X6 U424 ( .A(\add_545/A[15] ), .B(n6), .Z(dma_rp_new[15]) );
  HS65_LS_IVX9 U425 ( .A(n875), .Z(\add_545/A[15] ) );
  HS65_LS_IVX18 U426 ( .A(\phase_prev[0] ), .Z(n453) );
  HS65_LS_NAND2X7 U427 ( .A(dma_rdata[51]), .B(n144), .Z(n837) );
  HS65_LS_NAND2X7 U428 ( .A(dma_rdata[52]), .B(n144), .Z(n838) );
  HS65_LS_NAND2X7 U429 ( .A(dma_rdata[55]), .B(n144), .Z(n839) );
  HS65_LS_NAND2X7 U430 ( .A(dma_rdata[56]), .B(n144), .Z(n840) );
  HS65_LS_NAND2X7 U431 ( .A(dma_rdata[58]), .B(n144), .Z(n841) );
  HS65_LS_NAND2X7 U432 ( .A(dma_rdata[49]), .B(n149), .Z(n862) );
  HS65_LS_NAND2X7 U433 ( .A(dma_rdata[50]), .B(n149), .Z(n861) );
  HS65_LS_NAND2X7 U434 ( .A(dma_rdata[53]), .B(n149), .Z(n860) );
  HS65_LS_NAND2X7 U435 ( .A(dma_rdata[54]), .B(n149), .Z(n859) );
  HS65_LS_NAND2X7 U436 ( .A(dma_rdata[57]), .B(n149), .Z(n858) );
  HS65_LS_NAND2X7 U437 ( .A(dma_rdata[59]), .B(n149), .Z(n857) );
  HS65_LH_OAI12X2 U438 ( .A(n20), .B(n684), .C(n325), .Z(phit_togo[34]) );
  HS65_LS_OAI21X3 U439 ( .A(n647), .B(n142), .C(n360), .Z(n362) );
  HS65_LS_IVX18 U440 ( .A(state_cnt[1]), .Z(n452) );
  HS65_LS_IVX9 U441 ( .A(dma_rdata[62]), .Z(n644) );
  HS65_LS_IVX18 U442 ( .A(state_cnt[0]), .Z(n448) );
  HS65_LS_AOI22X6 U443 ( .A(\proc_in[MADDR][0] ), .B(n651), .C(
        \proc_in[MADDR][1] ), .D(n834), .Z(n832) );
  HS65_LS_NAND2X7 U444 ( .A(phitIn[33]), .B(phitIn[34]), .Z(n863) );
  HS65_LS_NAND3X5 U445 ( .A(n128), .B(n576), .C(n306), .Z(n363) );
  HS65_LS_NAND3AX6 U446 ( .A(phitIn[33]), .B(phitIn[32]), .C(phitIn[34]), .Z(
        n865) );
  HS65_LS_NAND2X7 U447 ( .A(dma_rdata[48]), .B(n144), .Z(n836) );
  HS65_LS_NAND2X7 U448 ( .A(dma_rdata[60]), .B(n144), .Z(n842) );
  HS65_LS_NAND2X7 U449 ( .A(dma_rdata[61]), .B(n144), .Z(n843) );
  HS65_LS_BFX9 U450 ( .A(n864), .Z(n298) );
  HS65_LS_NOR3AX2 U451 ( .A(phitIn[34]), .B(phitIn[32]), .C(phitIn[33]), .Z(
        n864) );
  HS65_LS_AO22X9 U452 ( .A(n863), .B(address[0]), .C(phitIn[17]), .D(n648), 
        .Z(n738) );
  HS65_LS_AO22X9 U453 ( .A(n863), .B(address[1]), .C(phitIn[18]), .D(n648), 
        .Z(n736) );
  HS65_LS_AO22X9 U454 ( .A(n863), .B(address[2]), .C(phitIn[19]), .D(n648), 
        .Z(n734) );
  HS65_LS_AO22X9 U455 ( .A(n863), .B(address[3]), .C(phitIn[20]), .D(n648), 
        .Z(n732) );
  HS65_LS_AO22X9 U456 ( .A(n863), .B(address[4]), .C(phitIn[21]), .D(n648), 
        .Z(n730) );
  HS65_LS_AO22X9 U457 ( .A(n863), .B(address[5]), .C(phitIn[22]), .D(n648), 
        .Z(n728) );
  HS65_LS_AO22X9 U458 ( .A(n863), .B(address[6]), .C(phitIn[23]), .D(n648), 
        .Z(n726) );
  HS65_LS_IVX9 U459 ( .A(slt_entry[3]), .Z(n645) );
  HS65_LS_IVX9 U460 ( .A(slt_entry[2]), .Z(n646) );
  HS65_LS_AO22X9 U461 ( .A(phitIn[0]), .B(n312), .C(\spm_out[MDATA][0] ), .D(
        n306), .Z(n827) );
  HS65_LS_AO22X9 U462 ( .A(phitIn[1]), .B(n323), .C(\spm_out[MDATA][1] ), .D(
        n306), .Z(n826) );
  HS65_LS_AO22X9 U463 ( .A(phitIn[2]), .B(n323), .C(\spm_out[MDATA][2] ), .D(
        n306), .Z(n825) );
  HS65_LS_AO22X9 U464 ( .A(phitIn[3]), .B(n323), .C(\spm_out[MDATA][3] ), .D(
        n305), .Z(n824) );
  HS65_LS_AO22X9 U465 ( .A(phitIn[4]), .B(n323), .C(\spm_out[MDATA][4] ), .D(
        n304), .Z(n823) );
  HS65_LS_AO22X9 U466 ( .A(phitIn[5]), .B(n323), .C(\spm_out[MDATA][5] ), .D(
        n865), .Z(n822) );
  HS65_LS_AO22X9 U467 ( .A(phitIn[6]), .B(n323), .C(\spm_out[MDATA][6] ), .D(
        n306), .Z(n821) );
  HS65_LS_AO22X9 U468 ( .A(phitIn[7]), .B(n323), .C(\spm_out[MDATA][7] ), .D(
        n865), .Z(n820) );
  HS65_LS_AO22X9 U469 ( .A(phitIn[8]), .B(n323), .C(\spm_out[MDATA][8] ), .D(
        n865), .Z(n819) );
  HS65_LS_AO22X9 U470 ( .A(phitIn[9]), .B(n323), .C(\spm_out[MDATA][9] ), .D(
        n865), .Z(n818) );
  HS65_LS_AO22X9 U471 ( .A(phitIn[10]), .B(n314), .C(\spm_out[MDATA][10] ), 
        .D(n865), .Z(n817) );
  HS65_LS_AO22X9 U472 ( .A(phitIn[11]), .B(n314), .C(\spm_out[MDATA][11] ), 
        .D(n865), .Z(n816) );
  HS65_LS_AO22X9 U473 ( .A(phitIn[12]), .B(n314), .C(\spm_out[MDATA][12] ), 
        .D(n865), .Z(n815) );
  HS65_LS_AO22X9 U474 ( .A(phitIn[13]), .B(n314), .C(\spm_out[MDATA][13] ), 
        .D(n865), .Z(n814) );
  HS65_LS_AO22X9 U475 ( .A(phitIn[14]), .B(n314), .C(\spm_out[MDATA][14] ), 
        .D(n865), .Z(n813) );
  HS65_LS_AO22X9 U476 ( .A(phitIn[15]), .B(n314), .C(\spm_out[MDATA][15] ), 
        .D(n865), .Z(n812) );
  HS65_LS_AO22X9 U477 ( .A(phitIn[16]), .B(n314), .C(\spm_out[MDATA][16] ), 
        .D(n865), .Z(n811) );
  HS65_LS_AO22X9 U478 ( .A(phitIn[17]), .B(n314), .C(\spm_out[MDATA][17] ), 
        .D(n865), .Z(n810) );
  HS65_LS_AO22X9 U479 ( .A(phitIn[18]), .B(n314), .C(\spm_out[MDATA][18] ), 
        .D(n865), .Z(n809) );
  HS65_LS_AO22X9 U480 ( .A(phitIn[19]), .B(n314), .C(\spm_out[MDATA][19] ), 
        .D(n306), .Z(n808) );
  HS65_LS_AO22X9 U481 ( .A(phitIn[20]), .B(n314), .C(\spm_out[MDATA][20] ), 
        .D(n306), .Z(n807) );
  HS65_LS_AO22X9 U482 ( .A(phitIn[21]), .B(n314), .C(\spm_out[MDATA][21] ), 
        .D(n306), .Z(n806) );
  HS65_LS_AO22X9 U483 ( .A(phitIn[22]), .B(n314), .C(\spm_out[MDATA][22] ), 
        .D(n306), .Z(n805) );
  HS65_LS_AO22X9 U484 ( .A(phitIn[23]), .B(n314), .C(\spm_out[MDATA][23] ), 
        .D(n306), .Z(n804) );
  HS65_LS_AO22X9 U485 ( .A(phitIn[24]), .B(n314), .C(\spm_out[MDATA][24] ), 
        .D(n306), .Z(n803) );
  HS65_LS_AO22X9 U486 ( .A(phitIn[25]), .B(n314), .C(\spm_out[MDATA][25] ), 
        .D(n306), .Z(n802) );
  HS65_LS_AO22X9 U487 ( .A(phitIn[26]), .B(n314), .C(\spm_out[MDATA][26] ), 
        .D(n306), .Z(n801) );
  HS65_LS_AO22X9 U488 ( .A(phitIn[27]), .B(n314), .C(\spm_out[MDATA][27] ), 
        .D(n306), .Z(n800) );
  HS65_LS_AO22X9 U489 ( .A(phitIn[28]), .B(n314), .C(\spm_out[MDATA][28] ), 
        .D(n306), .Z(n799) );
  HS65_LS_AO22X9 U490 ( .A(phitIn[29]), .B(n314), .C(\spm_out[MDATA][29] ), 
        .D(n306), .Z(n798) );
  HS65_LS_AO22X9 U491 ( .A(phitIn[30]), .B(n313), .C(\spm_out[MDATA][30] ), 
        .D(n306), .Z(n797) );
  HS65_LS_AO22X9 U492 ( .A(phitIn[31]), .B(n313), .C(\spm_out[MDATA][31] ), 
        .D(n306), .Z(n796) );
  HS65_LS_AO22X9 U493 ( .A(dIn_h[0]), .B(n313), .C(\spm_out[MDATA][32] ), .D(
        n305), .Z(n795) );
  HS65_LS_AO22X9 U494 ( .A(dIn_h[1]), .B(n313), .C(\spm_out[MDATA][33] ), .D(
        n305), .Z(n794) );
  HS65_LS_AO22X9 U495 ( .A(dIn_h[2]), .B(n313), .C(\spm_out[MDATA][34] ), .D(
        n305), .Z(n793) );
  HS65_LS_AO22X9 U496 ( .A(dIn_h[3]), .B(n313), .C(\spm_out[MDATA][35] ), .D(
        n305), .Z(n792) );
  HS65_LS_AO22X9 U497 ( .A(dIn_h[4]), .B(n313), .C(\spm_out[MDATA][36] ), .D(
        n305), .Z(n791) );
  HS65_LS_AO22X9 U498 ( .A(dIn_h[5]), .B(n313), .C(\spm_out[MDATA][37] ), .D(
        n305), .Z(n790) );
  HS65_LS_AO22X9 U499 ( .A(dIn_h[6]), .B(n313), .C(\spm_out[MDATA][38] ), .D(
        n305), .Z(n789) );
  HS65_LS_AO22X9 U500 ( .A(dIn_h[7]), .B(n313), .C(\spm_out[MDATA][39] ), .D(
        n305), .Z(n788) );
  HS65_LS_AO22X9 U501 ( .A(dIn_h[8]), .B(n313), .C(\spm_out[MDATA][40] ), .D(
        n305), .Z(n787) );
  HS65_LS_AO22X9 U502 ( .A(dIn_h[9]), .B(n313), .C(\spm_out[MDATA][41] ), .D(
        n305), .Z(n786) );
  HS65_LS_AO22X9 U503 ( .A(dIn_h[10]), .B(n313), .C(\spm_out[MDATA][42] ), .D(
        n305), .Z(n785) );
  HS65_LS_AO22X9 U504 ( .A(dIn_h[11]), .B(n313), .C(\spm_out[MDATA][43] ), .D(
        n305), .Z(n784) );
  HS65_LS_AO22X9 U505 ( .A(dIn_h[12]), .B(n313), .C(\spm_out[MDATA][44] ), .D(
        n304), .Z(n783) );
  HS65_LS_AO22X9 U506 ( .A(dIn_h[13]), .B(n313), .C(\spm_out[MDATA][45] ), .D(
        n304), .Z(n782) );
  HS65_LS_AO22X9 U507 ( .A(dIn_h[14]), .B(n313), .C(\spm_out[MDATA][46] ), .D(
        n304), .Z(n781) );
  HS65_LS_AO22X9 U508 ( .A(dIn_h[15]), .B(n313), .C(\spm_out[MDATA][47] ), .D(
        n304), .Z(n780) );
  HS65_LS_AO22X9 U509 ( .A(dIn_h[16]), .B(n313), .C(\spm_out[MDATA][48] ), .D(
        n304), .Z(n779) );
  HS65_LS_AO22X9 U510 ( .A(dIn_h[17]), .B(n312), .C(\spm_out[MDATA][49] ), .D(
        n304), .Z(n778) );
  HS65_LS_AO22X9 U511 ( .A(dIn_h[18]), .B(n312), .C(\spm_out[MDATA][50] ), .D(
        n304), .Z(n777) );
  HS65_LS_AO22X9 U512 ( .A(dIn_h[19]), .B(n312), .C(\spm_out[MDATA][51] ), .D(
        n304), .Z(n776) );
  HS65_LS_AO22X9 U513 ( .A(dIn_h[20]), .B(n313), .C(\spm_out[MDATA][52] ), .D(
        n304), .Z(n775) );
  HS65_LS_AO22X9 U514 ( .A(dIn_h[21]), .B(n312), .C(\spm_out[MDATA][53] ), .D(
        n305), .Z(n774) );
  HS65_LS_AO22X9 U515 ( .A(dIn_h[22]), .B(n312), .C(\spm_out[MDATA][54] ), .D(
        n304), .Z(n773) );
  HS65_LS_AO22X9 U516 ( .A(dIn_h[23]), .B(n312), .C(\spm_out[MDATA][55] ), .D(
        n304), .Z(n772) );
  HS65_LS_AO22X9 U517 ( .A(dIn_h[24]), .B(n312), .C(\spm_out[MDATA][56] ), .D(
        n304), .Z(n771) );
  HS65_LS_AO22X9 U518 ( .A(dIn_h[25]), .B(n312), .C(\spm_out[MDATA][57] ), .D(
        n304), .Z(n770) );
  HS65_LS_AO22X9 U519 ( .A(dIn_h[26]), .B(n312), .C(\spm_out[MDATA][58] ), .D(
        n304), .Z(n769) );
  HS65_LS_AO22X9 U520 ( .A(dIn_h[27]), .B(n312), .C(\spm_out[MDATA][59] ), .D(
        n305), .Z(n768) );
  HS65_LS_AO22X9 U521 ( .A(dIn_h[28]), .B(n312), .C(\spm_out[MDATA][60] ), .D(
        n304), .Z(n767) );
  HS65_LS_AO22X9 U522 ( .A(dIn_h[29]), .B(n312), .C(\spm_out[MDATA][61] ), .D(
        n305), .Z(n766) );
  HS65_LS_AO22X9 U523 ( .A(dIn_h[30]), .B(n312), .C(\spm_out[MDATA][62] ), .D(
        n304), .Z(n765) );
  HS65_LS_AO22X9 U524 ( .A(dIn_h[31]), .B(n312), .C(\spm_out[MDATA][63] ), .D(
        n306), .Z(n764) );
  HS65_LS_AO22X9 U525 ( .A(phitIn[17]), .B(n302), .C(n300), .D(dIn_h[17]), .Z(
        n739) );
  HS65_LS_AO22X9 U526 ( .A(phitIn[18]), .B(n302), .C(n300), .D(dIn_h[18]), .Z(
        n737) );
  HS65_LS_AO22X9 U527 ( .A(phitIn[19]), .B(n302), .C(n300), .D(dIn_h[19]), .Z(
        n735) );
  HS65_LS_AO22X9 U528 ( .A(phitIn[20]), .B(n302), .C(n300), .D(dIn_h[20]), .Z(
        n733) );
  HS65_LS_AO22X9 U529 ( .A(phitIn[21]), .B(n303), .C(n300), .D(dIn_h[21]), .Z(
        n731) );
  HS65_LS_AO22X9 U530 ( .A(phitIn[22]), .B(n303), .C(n300), .D(dIn_h[22]), .Z(
        n729) );
  HS65_LS_AO22X9 U531 ( .A(phitIn[23]), .B(n303), .C(n300), .D(dIn_h[23]), .Z(
        n727) );
  HS65_LS_AO22X9 U532 ( .A(phitIn[0]), .B(n301), .C(n299), .D(dIn_h[0]), .Z(
        n756) );
  HS65_LS_AO22X9 U533 ( .A(phitIn[1]), .B(n302), .C(n299), .D(dIn_h[1]), .Z(
        n755) );
  HS65_LS_AO22X9 U534 ( .A(phitIn[2]), .B(n302), .C(n299), .D(dIn_h[2]), .Z(
        n754) );
  HS65_LS_AO22X9 U535 ( .A(phitIn[3]), .B(n302), .C(n299), .D(dIn_h[3]), .Z(
        n753) );
  HS65_LS_AO22X9 U536 ( .A(phitIn[4]), .B(n302), .C(n299), .D(dIn_h[4]), .Z(
        n752) );
  HS65_LS_AO22X9 U537 ( .A(phitIn[5]), .B(n302), .C(n299), .D(dIn_h[5]), .Z(
        n751) );
  HS65_LS_AO22X9 U538 ( .A(phitIn[6]), .B(n302), .C(n299), .D(dIn_h[6]), .Z(
        n750) );
  HS65_LS_AO22X9 U539 ( .A(phitIn[7]), .B(n302), .C(n299), .D(dIn_h[7]), .Z(
        n749) );
  HS65_LS_AO22X9 U540 ( .A(phitIn[8]), .B(n302), .C(n299), .D(dIn_h[8]), .Z(
        n748) );
  HS65_LS_AO22X9 U541 ( .A(phitIn[9]), .B(n302), .C(n299), .D(dIn_h[9]), .Z(
        n747) );
  HS65_LS_AO22X9 U542 ( .A(phitIn[10]), .B(n302), .C(n299), .D(dIn_h[10]), .Z(
        n746) );
  HS65_LS_AO22X9 U543 ( .A(phitIn[11]), .B(n302), .C(n299), .D(dIn_h[11]), .Z(
        n745) );
  HS65_LS_AO22X9 U544 ( .A(phitIn[12]), .B(n302), .C(n299), .D(dIn_h[12]), .Z(
        n744) );
  HS65_LS_AO22X9 U545 ( .A(phitIn[13]), .B(n302), .C(n300), .D(dIn_h[13]), .Z(
        n743) );
  HS65_LS_AO22X9 U546 ( .A(phitIn[14]), .B(n302), .C(n300), .D(dIn_h[14]), .Z(
        n742) );
  HS65_LS_AO22X9 U547 ( .A(phitIn[15]), .B(n302), .C(n300), .D(dIn_h[15]), .Z(
        n741) );
  HS65_LS_AO22X9 U548 ( .A(phitIn[16]), .B(n302), .C(n300), .D(dIn_h[16]), .Z(
        n740) );
  HS65_LS_AO22X9 U549 ( .A(phitIn[24]), .B(n303), .C(n300), .D(dIn_h[24]), .Z(
        n725) );
  HS65_LS_AO22X9 U550 ( .A(phitIn[25]), .B(n303), .C(n300), .D(dIn_h[25]), .Z(
        n724) );
  HS65_LS_AO22X9 U551 ( .A(phitIn[26]), .B(n303), .C(n299), .D(dIn_h[26]), .Z(
        n723) );
  HS65_LS_AO22X9 U552 ( .A(phitIn[27]), .B(n303), .C(n300), .D(dIn_h[27]), .Z(
        n722) );
  HS65_LS_AO22X9 U553 ( .A(phitIn[28]), .B(n303), .C(n299), .D(dIn_h[28]), .Z(
        n721) );
  HS65_LS_AO22X9 U554 ( .A(phitIn[29]), .B(n303), .C(n300), .D(dIn_h[29]), .Z(
        n720) );
  HS65_LS_AO22X9 U555 ( .A(phitIn[30]), .B(n303), .C(n299), .D(dIn_h[30]), .Z(
        n719) );
  HS65_LS_AO22X9 U556 ( .A(phitIn[31]), .B(n303), .C(n300), .D(dIn_h[31]), .Z(
        n718) );
  HS65_LS_AO22X9 U557 ( .A(n312), .B(address[0]), .C(n305), .D(flit_buf[64]), 
        .Z(n763) );
  HS65_LS_AO22X9 U558 ( .A(n312), .B(address[1]), .C(n304), .D(flit_buf[65]), 
        .Z(n762) );
  HS65_LS_AO22X9 U559 ( .A(n312), .B(address[2]), .C(n305), .D(flit_buf[66]), 
        .Z(n761) );
  HS65_LS_AO22X9 U560 ( .A(n312), .B(address[3]), .C(n304), .D(flit_buf[67]), 
        .Z(n760) );
  HS65_LS_AO22X9 U561 ( .A(n311), .B(address[4]), .C(n305), .D(flit_buf[68]), 
        .Z(n759) );
  HS65_LS_AO22X9 U562 ( .A(n310), .B(address[5]), .C(n304), .D(flit_buf[69]), 
        .Z(n758) );
  HS65_LS_AO22X9 U563 ( .A(n312), .B(address[6]), .C(n305), .D(flit_buf[70]), 
        .Z(n757) );
  HS65_LS_OR2X9 U564 ( .A(vld_pkt), .B(n648), .Z(n679) );
  HS65_LS_NAND2X7 U565 ( .A(\proc_in[MADDR][0] ), .B(n831), .Z(n856) );
  HS65_LS_NOR4ABX2 U566 ( .A(n655), .B(n828), .C(\proc_in[MADDR][26] ), .D(
        \proc_in[MADDR][24] ), .Z(n855) );
  HS65_LS_IVX9 U567 ( .A(\proc_in[MADDR][25] ), .Z(n655) );
  HS65_LS_NOR3X4 U568 ( .A(\proc_in[MADDR][27] ), .B(\proc_in[MADDR][31] ), 
        .C(\proc_in[MADDR][30] ), .Z(n828) );
  HS65_LS_NAND4ABX3 U569 ( .A(\proc_in[MADDR][29] ), .B(\proc_in[MADDR][26] ), 
        .C(n830), .D(n829), .Z(n853) );
  HS65_LS_NOR2X6 U570 ( .A(\proc_in[MADDR][31] ), .B(\proc_in[MADDR][30] ), 
        .Z(n830) );
  HS65_LS_NOR4ABX2 U571 ( .A(\proc_in[MADDR][28] ), .B(\proc_in[MADDR][27] ), 
        .C(\proc_in[MADDR][25] ), .D(\proc_in[MADDR][24] ), .Z(n829) );
  HS65_LS_NOR3AX2 U572 ( .A(n855), .B(n654), .C(\proc_in[MADDR][29] ), .Z(n675) );
  HS65_LS_NAND4ABX3 U573 ( .A(config_reg[3]), .B(n869), .C(config_reg[4]), .D(
        n592), .Z(n870) );
  HS65_LS_OA32X4 U574 ( .A(config_reg[0]), .B(config_reg[1]), .C(n649), .D(
        n868), .E(config_reg[2]), .Z(n869) );
  HS65_LS_IVX9 U575 ( .A(config_reg[2]), .Z(n649) );
  HS65_LSS_XNOR2X6 U576 ( .A(config_reg[1]), .B(config_reg[0]), .Z(n868) );
  HS65_LS_BFX9 U577 ( .A(na_reset), .Z(n339) );
  HS65_LS_BFX9 U578 ( .A(na_reset), .Z(n340) );
  HS65_LS_NAND2X7 U579 ( .A(n675), .B(\proc_in[MCMD][0] ), .Z(n867) );
  HS65_LS_IVX9 U580 ( .A(\proc_in[MDATA][15] ), .Z(n659) );
  HS65_LS_IVX9 U581 ( .A(\proc_in[MDATA][6] ), .Z(n668) );
  HS65_LS_IVX9 U582 ( .A(\proc_in[MDATA][7] ), .Z(n667) );
  HS65_LS_IVX9 U583 ( .A(\proc_in[MDATA][8] ), .Z(n666) );
  HS65_LS_IVX9 U584 ( .A(\proc_in[MDATA][9] ), .Z(n665) );
  HS65_LS_IVX9 U585 ( .A(\proc_in[MADDR][28] ), .Z(n654) );
  HS65_LS_AND3X9 U586 ( .A(n855), .B(n654), .C(\proc_in[MADDR][29] ), .Z(n831)
         );
  HS65_LS_IVX9 U587 ( .A(\proc_in[MDATA][14] ), .Z(n660) );
  HS65_LS_IVX9 U588 ( .A(\proc_in[MDATA][0] ), .Z(n674) );
  HS65_LS_IVX9 U589 ( .A(\proc_in[MDATA][1] ), .Z(n673) );
  HS65_LS_IVX9 U590 ( .A(\proc_in[MDATA][2] ), .Z(n672) );
  HS65_LS_IVX9 U591 ( .A(\proc_in[MDATA][3] ), .Z(n671) );
  HS65_LS_IVX9 U592 ( .A(\proc_in[MDATA][4] ), .Z(n670) );
  HS65_LS_IVX9 U593 ( .A(\proc_in[MDATA][5] ), .Z(n669) );
  HS65_LS_IVX9 U594 ( .A(\proc_in[MDATA][10] ), .Z(n664) );
  HS65_LS_IVX9 U595 ( .A(\proc_in[MDATA][11] ), .Z(n663) );
  HS65_LS_IVX9 U596 ( .A(\proc_in[MDATA][12] ), .Z(n662) );
  HS65_LS_IVX9 U597 ( .A(\proc_in[MDATA][13] ), .Z(n661) );
  HS65_LS_IVX9 U598 ( .A(\proc_in[MADDR][0] ), .Z(n658) );
  HS65_LS_IVX9 U599 ( .A(\proc_in[MADDR][1] ), .Z(n657) );
  HS65_LH_MUX21I1X3 U600 ( .D0(n1), .D1(n454), .S0(n647), .Z(n682) );
  HS65_LS_IVX18 U601 ( .A(n476), .Z(n513) );
  HS65_LS_NAND2X2 U602 ( .A(phitOut2[8]), .B(n513), .Z(n492) );
  HS65_LS_NAND2X2 U603 ( .A(phitOut2[9]), .B(n44), .Z(n495) );
  HS65_LS_NAND2X2 U604 ( .A(phitOut2[6]), .B(n513), .Z(n486) );
  HS65_LS_NAND2X2 U605 ( .A(phitOut2[5]), .B(n513), .Z(n483) );
  HS65_LS_NAND2X2 U606 ( .A(phitOut2[4]), .B(n513), .Z(n480) );
  HS65_LS_NAND2X2 U607 ( .A(phitOut2[12]), .B(n513), .Z(n504) );
  HS65_LS_NAND2X2 U608 ( .A(phitOut2[13]), .B(n513), .Z(n507) );
  HS65_LS_NAND2X2 U609 ( .A(phitOut2[14]), .B(n513), .Z(n510) );
  HS65_LS_NAND2X2 U610 ( .A(phitOut2[15]), .B(n513), .Z(n514) );
  HS65_LS_AOI33X2 U611 ( .A(n572), .B(n27), .C(phitOut2[34]), .D(n111), .E(n27), .F(phitOut0[34]), .Z(n573) );
  HS65_LS_IVX9 U612 ( .A(n139), .Z(n128) );
  HS65_LH_BFX2 U613 ( .A(n113), .Z(n139) );
  HS65_LS_BFX9 U614 ( .A(n139), .Z(n142) );
  HS65_LS_BFX9 U615 ( .A(n139), .Z(n140) );
  HS65_LH_CBI4I1X3 U616 ( .A(n128), .B(n364), .C(n306), .D(n363), .Z(n680) );
  HS65_LS_IVX9 U617 ( .A(n451), .Z(n647) );
  HS65_LS_IVX9 U618 ( .A(n851), .Z(n620) );
  HS65_LS_NAND2X7 U619 ( .A(dma_rdata[39]), .B(n149), .Z(n590) );
  HS65_LS_IVX9 U620 ( .A(n590), .Z(n619) );
  HS65_LS_NAND2X7 U621 ( .A(dma_rdata[38]), .B(n149), .Z(n588) );
  HS65_LS_IVX9 U622 ( .A(n588), .Z(n618) );
  HS65_LS_NAND2X7 U623 ( .A(dma_rdata[37]), .B(n293), .Z(n586) );
  HS65_LS_IVX9 U624 ( .A(n586), .Z(n617) );
  HS65_LS_NAND2X7 U625 ( .A(dma_rdata[36]), .B(n293), .Z(n584) );
  HS65_LS_IVX9 U626 ( .A(n584), .Z(n616) );
  HS65_LS_NAND2X7 U627 ( .A(dma_rdata[35]), .B(n293), .Z(n582) );
  HS65_LS_IVX9 U628 ( .A(n582), .Z(n615) );
  HS65_LS_NAND2X7 U629 ( .A(dma_rdata[34]), .B(n293), .Z(n580) );
  HS65_LS_IVX9 U630 ( .A(n580), .Z(n614) );
  HS65_LS_NAND2X7 U631 ( .A(dma_rdata[33]), .B(n293), .Z(n578) );
  HS65_LS_IVX9 U632 ( .A(n578), .Z(n613) );
  HS65_LS_NAND2X7 U633 ( .A(dma_rdata[31]), .B(n293), .Z(n413) );
  HS65_LS_IVX9 U634 ( .A(n413), .Z(n612) );
  HS65_LS_NAND2X7 U635 ( .A(dma_rdata[30]), .B(n293), .Z(n411) );
  HS65_LS_IVX9 U636 ( .A(n411), .Z(n611) );
  HS65_LS_NAND2X7 U637 ( .A(dma_rdata[29]), .B(n293), .Z(n409) );
  HS65_LS_IVX9 U638 ( .A(n409), .Z(n610) );
  HS65_LS_NAND2X7 U639 ( .A(dma_rdata[28]), .B(n293), .Z(n407) );
  HS65_LS_IVX9 U640 ( .A(n407), .Z(n609) );
  HS65_LS_NAND2X7 U641 ( .A(dma_rdata[27]), .B(n293), .Z(n405) );
  HS65_LS_IVX9 U642 ( .A(n405), .Z(n608) );
  HS65_LS_NAND2X7 U643 ( .A(dma_rdata[26]), .B(n293), .Z(n403) );
  HS65_LS_IVX9 U644 ( .A(n403), .Z(n607) );
  HS65_LS_NAND2X7 U645 ( .A(dma_rdata[25]), .B(n293), .Z(n401) );
  HS65_LS_IVX9 U646 ( .A(n401), .Z(n606) );
  HS65_LS_NAND2X7 U647 ( .A(dma_rdata[24]), .B(n293), .Z(n399) );
  HS65_LS_IVX9 U648 ( .A(n399), .Z(n605) );
  HS65_LS_NAND2X7 U649 ( .A(dma_rdata[23]), .B(n293), .Z(n397) );
  HS65_LS_IVX9 U650 ( .A(n397), .Z(n604) );
  HS65_LS_NAND2X7 U651 ( .A(dma_rdata[22]), .B(n293), .Z(n395) );
  HS65_LS_IVX9 U652 ( .A(n395), .Z(n603) );
  HS65_LS_NAND2X7 U653 ( .A(dma_rdata[21]), .B(n293), .Z(n393) );
  HS65_LS_IVX9 U654 ( .A(n393), .Z(n602) );
  HS65_LS_NAND2X7 U655 ( .A(dma_rdata[20]), .B(n293), .Z(n391) );
  HS65_LS_IVX9 U656 ( .A(n391), .Z(n601) );
  HS65_LS_NAND2X7 U657 ( .A(dma_rdata[19]), .B(n149), .Z(n389) );
  HS65_LS_IVX9 U658 ( .A(n389), .Z(n600) );
  HS65_LS_NAND2X7 U659 ( .A(dma_rdata[18]), .B(n149), .Z(n387) );
  HS65_LS_IVX9 U660 ( .A(n387), .Z(n599) );
  HS65_LS_NAND2X7 U661 ( .A(dma_rdata[17]), .B(n149), .Z(n385) );
  HS65_LS_IVX9 U662 ( .A(n385), .Z(n598) );
  HS65_LS_IVX9 U663 ( .A(\proc_in[MCMD][0] ), .Z(n360) );
  HS65_LS_IVX9 U664 ( .A(n362), .Z(n361) );
  HS65_LS_NAND2X7 U665 ( .A(n834), .B(n4), .Z(n852) );
  HS65_LS_OAI22X6 U666 ( .A(n645), .B(n365), .C(n833), .D(n362), .Z(
        dma_raddr[1]) );
  HS65_LS_OAI22X6 U667 ( .A(n646), .B(n365), .C(n832), .D(n362), .Z(
        dma_raddr[0]) );
  HS65_LS_NAND2X7 U668 ( .A(dma_rdata[16]), .B(n149), .Z(n383) );
  HS65_LS_IVX9 U669 ( .A(n383), .Z(n595) );
  HS65_LS_IVX9 U670 ( .A(n685), .Z(n454) );
  HS65_LS_IVX9 U671 ( .A(vld_pkt), .Z(n364) );
  HS65_LS_IVX9 U672 ( .A(n683), .Z(n576) );
  HS65_LS_IVX9 U673 ( .A(n365), .Z(n597) );
  HS65_LS_IVX9 U674 ( .A(n684), .Z(n415) );
  HS65_LS_NAND2X7 U675 ( .A(n597), .B(n415), .Z(n414) );
  HS65_LS_IVX9 U676 ( .A(dOut_l[0]), .Z(n416) );
  HS65_LS_NAND2X7 U677 ( .A(\spm_in[SDATA][32] ), .B(n130), .Z(n366) );
  HS65_LS_OAI212X5 U678 ( .A(n136), .B(n416), .C(n329), .D(n642), .E(n366), 
        .Z(mux_out[0]) );
  HS65_LS_IVX9 U679 ( .A(dOut_l[1]), .Z(n417) );
  HS65_LS_NAND2X7 U680 ( .A(\spm_in[SDATA][33] ), .B(n130), .Z(n367) );
  HS65_LS_OAI212X5 U681 ( .A(n136), .B(n417), .C(n329), .D(n641), .E(n367), 
        .Z(mux_out[1]) );
  HS65_LS_IVX9 U682 ( .A(dOut_l[2]), .Z(n418) );
  HS65_LS_NAND2X7 U683 ( .A(\spm_in[SDATA][34] ), .B(n130), .Z(n368) );
  HS65_LS_OAI212X5 U684 ( .A(n136), .B(n418), .C(n329), .D(n640), .E(n368), 
        .Z(mux_out[2]) );
  HS65_LS_IVX9 U685 ( .A(dOut_l[3]), .Z(n419) );
  HS65_LS_NAND2X7 U686 ( .A(\spm_in[SDATA][35] ), .B(n130), .Z(n369) );
  HS65_LS_OAI212X5 U687 ( .A(n136), .B(n419), .C(n329), .D(n639), .E(n369), 
        .Z(mux_out[3]) );
  HS65_LS_IVX9 U688 ( .A(dOut_l[4]), .Z(n420) );
  HS65_LS_NAND2X7 U689 ( .A(\spm_in[SDATA][36] ), .B(n130), .Z(n370) );
  HS65_LS_OAI212X5 U690 ( .A(n136), .B(n420), .C(n329), .D(n638), .E(n370), 
        .Z(mux_out[4]) );
  HS65_LS_IVX9 U691 ( .A(dOut_l[5]), .Z(n421) );
  HS65_LS_NAND2X7 U692 ( .A(\spm_in[SDATA][37] ), .B(n130), .Z(n371) );
  HS65_LS_OAI212X5 U693 ( .A(n136), .B(n421), .C(n329), .D(n637), .E(n371), 
        .Z(mux_out[5]) );
  HS65_LS_IVX9 U694 ( .A(dOut_l[6]), .Z(n422) );
  HS65_LS_NAND2X7 U695 ( .A(\spm_in[SDATA][38] ), .B(n130), .Z(n372) );
  HS65_LS_OAI212X5 U696 ( .A(n136), .B(n422), .C(n329), .D(n636), .E(n372), 
        .Z(mux_out[6]) );
  HS65_LS_IVX9 U697 ( .A(dOut_l[7]), .Z(n423) );
  HS65_LS_NAND2X7 U698 ( .A(\spm_in[SDATA][39] ), .B(n130), .Z(n373) );
  HS65_LS_OAI212X5 U699 ( .A(n136), .B(n423), .C(n329), .D(n635), .E(n373), 
        .Z(mux_out[7]) );
  HS65_LS_IVX9 U700 ( .A(dOut_l[8]), .Z(n424) );
  HS65_LS_NAND2X7 U701 ( .A(\spm_in[SDATA][40] ), .B(n130), .Z(n374) );
  HS65_LS_OAI212X5 U702 ( .A(n136), .B(n424), .C(n329), .D(n634), .E(n374), 
        .Z(mux_out[8]) );
  HS65_LS_IVX9 U703 ( .A(dOut_l[9]), .Z(n425) );
  HS65_LS_NAND2X7 U704 ( .A(\spm_in[SDATA][41] ), .B(n130), .Z(n375) );
  HS65_LS_OAI212X5 U705 ( .A(n136), .B(n425), .C(n328), .D(n633), .E(n375), 
        .Z(mux_out[9]) );
  HS65_LS_IVX9 U706 ( .A(dOut_l[10]), .Z(n426) );
  HS65_LS_NAND2X7 U707 ( .A(\spm_in[SDATA][42] ), .B(n130), .Z(n376) );
  HS65_LS_OAI212X5 U708 ( .A(n136), .B(n426), .C(n328), .D(n632), .E(n376), 
        .Z(mux_out[10]) );
  HS65_LS_IVX9 U709 ( .A(dOut_l[11]), .Z(n427) );
  HS65_LS_NAND2X7 U710 ( .A(\spm_in[SDATA][43] ), .B(n130), .Z(n377) );
  HS65_LS_OAI212X5 U711 ( .A(n136), .B(n427), .C(n328), .D(n631), .E(n377), 
        .Z(mux_out[11]) );
  HS65_LS_IVX9 U712 ( .A(dOut_l[12]), .Z(n428) );
  HS65_LS_NAND2X7 U713 ( .A(\spm_in[SDATA][44] ), .B(n132), .Z(n378) );
  HS65_LS_OAI212X5 U714 ( .A(n137), .B(n428), .C(n328), .D(n630), .E(n378), 
        .Z(mux_out[12]) );
  HS65_LS_IVX9 U715 ( .A(dOut_l[13]), .Z(n429) );
  HS65_LS_NAND2X7 U716 ( .A(\spm_in[SDATA][45] ), .B(n132), .Z(n379) );
  HS65_LS_OAI212X5 U717 ( .A(n137), .B(n429), .C(n328), .D(n629), .E(n379), 
        .Z(mux_out[13]) );
  HS65_LS_IVX9 U718 ( .A(dOut_l[14]), .Z(n430) );
  HS65_LS_NAND2X7 U719 ( .A(\spm_in[SDATA][46] ), .B(n132), .Z(n380) );
  HS65_LS_OAI212X5 U720 ( .A(n137), .B(n430), .C(n328), .D(n628), .E(n380), 
        .Z(mux_out[14]) );
  HS65_LS_IVX9 U721 ( .A(dOut_l[15]), .Z(n431) );
  HS65_LS_NAND2X7 U722 ( .A(\spm_in[SDATA][47] ), .B(n132), .Z(n381) );
  HS65_LS_OAI212X5 U723 ( .A(n137), .B(n431), .C(n328), .D(n627), .E(n381), 
        .Z(mux_out[15]) );
  HS65_LS_IVX9 U724 ( .A(dOut_l[16]), .Z(n432) );
  HS65_LS_NAND2X7 U725 ( .A(\spm_in[SDATA][48] ), .B(n132), .Z(n382) );
  HS65_LS_OAI212X5 U726 ( .A(n137), .B(n432), .C(n328), .D(n383), .E(n382), 
        .Z(mux_out[16]) );
  HS65_LS_IVX9 U727 ( .A(dOut_l[17]), .Z(n433) );
  HS65_LS_NAND2X7 U728 ( .A(\spm_in[SDATA][49] ), .B(n132), .Z(n384) );
  HS65_LS_OAI212X5 U729 ( .A(n137), .B(n433), .C(n328), .D(n385), .E(n384), 
        .Z(mux_out[17]) );
  HS65_LS_IVX9 U730 ( .A(dOut_l[18]), .Z(n434) );
  HS65_LS_NAND2X7 U731 ( .A(\spm_in[SDATA][50] ), .B(n132), .Z(n386) );
  HS65_LS_OAI212X5 U732 ( .A(n137), .B(n434), .C(n328), .D(n387), .E(n386), 
        .Z(mux_out[18]) );
  HS65_LS_IVX9 U733 ( .A(dOut_l[19]), .Z(n435) );
  HS65_LS_NAND2X7 U734 ( .A(\spm_in[SDATA][51] ), .B(n132), .Z(n388) );
  HS65_LS_OAI212X5 U735 ( .A(n137), .B(n435), .C(n328), .D(n389), .E(n388), 
        .Z(mux_out[19]) );
  HS65_LS_IVX9 U736 ( .A(dOut_l[20]), .Z(n436) );
  HS65_LS_NAND2X7 U737 ( .A(\spm_in[SDATA][52] ), .B(n132), .Z(n390) );
  HS65_LS_OAI212X5 U738 ( .A(n137), .B(n436), .C(n328), .D(n391), .E(n390), 
        .Z(mux_out[20]) );
  HS65_LS_IVX9 U739 ( .A(dOut_l[21]), .Z(n437) );
  HS65_LS_NAND2X7 U740 ( .A(\spm_in[SDATA][53] ), .B(n132), .Z(n392) );
  HS65_LS_OAI212X5 U741 ( .A(n137), .B(n437), .C(n328), .D(n393), .E(n392), 
        .Z(mux_out[21]) );
  HS65_LS_IVX9 U742 ( .A(dOut_l[22]), .Z(n438) );
  HS65_LS_NAND2X7 U743 ( .A(\spm_in[SDATA][54] ), .B(n132), .Z(n394) );
  HS65_LS_OAI212X5 U744 ( .A(n137), .B(n438), .C(n328), .D(n395), .E(n394), 
        .Z(mux_out[22]) );
  HS65_LS_IVX9 U745 ( .A(dOut_l[23]), .Z(n439) );
  HS65_LS_NAND2X7 U746 ( .A(\spm_in[SDATA][55] ), .B(n132), .Z(n396) );
  HS65_LS_OAI212X5 U747 ( .A(n137), .B(n439), .C(n328), .D(n397), .E(n396), 
        .Z(mux_out[23]) );
  HS65_LS_IVX9 U748 ( .A(dOut_l[24]), .Z(n440) );
  HS65_LS_NAND2X7 U749 ( .A(\spm_in[SDATA][56] ), .B(n133), .Z(n398) );
  HS65_LS_OAI212X5 U750 ( .A(n138), .B(n440), .C(n328), .D(n399), .E(n398), 
        .Z(mux_out[24]) );
  HS65_LS_IVX9 U751 ( .A(dOut_l[25]), .Z(n441) );
  HS65_LS_NAND2X7 U752 ( .A(\spm_in[SDATA][57] ), .B(n133), .Z(n400) );
  HS65_LS_OAI212X5 U753 ( .A(n138), .B(n441), .C(n328), .D(n401), .E(n400), 
        .Z(mux_out[25]) );
  HS65_LS_IVX9 U754 ( .A(dOut_l[26]), .Z(n442) );
  HS65_LS_NAND2X7 U755 ( .A(\spm_in[SDATA][58] ), .B(n133), .Z(n402) );
  HS65_LS_OAI212X5 U756 ( .A(n138), .B(n442), .C(n328), .D(n403), .E(n402), 
        .Z(mux_out[26]) );
  HS65_LS_IVX9 U757 ( .A(dOut_l[27]), .Z(n443) );
  HS65_LS_NAND2X7 U758 ( .A(\spm_in[SDATA][59] ), .B(n133), .Z(n404) );
  HS65_LS_OAI212X5 U759 ( .A(n138), .B(n443), .C(n327), .D(n405), .E(n404), 
        .Z(mux_out[27]) );
  HS65_LS_IVX9 U760 ( .A(dOut_l[28]), .Z(n444) );
  HS65_LS_NAND2X7 U761 ( .A(\spm_in[SDATA][60] ), .B(n133), .Z(n406) );
  HS65_LS_OAI212X5 U762 ( .A(n138), .B(n444), .C(n328), .D(n407), .E(n406), 
        .Z(mux_out[28]) );
  HS65_LS_IVX9 U763 ( .A(dOut_l[29]), .Z(n445) );
  HS65_LS_NAND2X7 U764 ( .A(\spm_in[SDATA][61] ), .B(n133), .Z(n408) );
  HS65_LS_OAI212X5 U765 ( .A(n138), .B(n445), .C(n327), .D(n409), .E(n408), 
        .Z(mux_out[29]) );
  HS65_LS_IVX9 U766 ( .A(dOut_l[30]), .Z(n446) );
  HS65_LS_NAND2X7 U767 ( .A(\spm_in[SDATA][62] ), .B(n133), .Z(n410) );
  HS65_LS_OAI212X5 U768 ( .A(n138), .B(n446), .C(n328), .D(n411), .E(n410), 
        .Z(mux_out[30]) );
  HS65_LS_IVX9 U769 ( .A(dOut_l[31]), .Z(n447) );
  HS65_LS_NAND2X7 U770 ( .A(\spm_in[SDATA][63] ), .B(n133), .Z(n412) );
  HS65_LS_OAI212X5 U771 ( .A(n138), .B(n447), .C(n327), .D(n413), .E(n412), 
        .Z(mux_out[31]) );
  HS65_LS_MUX21I1X6 U772 ( .D0(n416), .D1(\spm_in[SDATA][0] ), .S0(n140), .Z(
        n717) );
  HS65_LS_MUX21I1X6 U773 ( .D0(n417), .D1(\spm_in[SDATA][1] ), .S0(n140), .Z(
        n716) );
  HS65_LS_MUX21I1X6 U774 ( .D0(n418), .D1(\spm_in[SDATA][2] ), .S0(n140), .Z(
        n715) );
  HS65_LS_MUX21I1X6 U775 ( .D0(n419), .D1(\spm_in[SDATA][3] ), .S0(n142), .Z(
        n714) );
  HS65_LS_MUX21I1X6 U776 ( .D0(n420), .D1(\spm_in[SDATA][4] ), .S0(n140), .Z(
        n713) );
  HS65_LS_MUX21I1X6 U777 ( .D0(n421), .D1(\spm_in[SDATA][5] ), .S0(n142), .Z(
        n712) );
  HS65_LS_MUX21I1X6 U778 ( .D0(n422), .D1(\spm_in[SDATA][6] ), .S0(n140), .Z(
        n711) );
  HS65_LS_MUX21I1X6 U779 ( .D0(n423), .D1(\spm_in[SDATA][7] ), .S0(n140), .Z(
        n710) );
  HS65_LS_MUX21I1X6 U780 ( .D0(n424), .D1(\spm_in[SDATA][8] ), .S0(n142), .Z(
        n709) );
  HS65_LS_MUX21I1X6 U781 ( .D0(n425), .D1(\spm_in[SDATA][9] ), .S0(n140), .Z(
        n708) );
  HS65_LS_MUX21I1X6 U782 ( .D0(n426), .D1(\spm_in[SDATA][10] ), .S0(n140), .Z(
        n707) );
  HS65_LS_MUX21I1X6 U783 ( .D0(n427), .D1(\spm_in[SDATA][11] ), .S0(n142), .Z(
        n706) );
  HS65_LS_MUX21I1X6 U784 ( .D0(n428), .D1(\spm_in[SDATA][12] ), .S0(n140), .Z(
        n705) );
  HS65_LS_MUX21I1X6 U785 ( .D0(n429), .D1(\spm_in[SDATA][13] ), .S0(n140), .Z(
        n704) );
  HS65_LS_MUX21I1X6 U786 ( .D0(n430), .D1(\spm_in[SDATA][14] ), .S0(n142), .Z(
        n703) );
  HS65_LS_MUX21I1X6 U787 ( .D0(n431), .D1(\spm_in[SDATA][15] ), .S0(n140), .Z(
        n702) );
  HS65_LS_MUX21I1X6 U788 ( .D0(n432), .D1(\spm_in[SDATA][16] ), .S0(n142), .Z(
        n701) );
  HS65_LS_MUX21I1X6 U789 ( .D0(n433), .D1(\spm_in[SDATA][17] ), .S0(n140), .Z(
        n700) );
  HS65_LS_MUX21I1X6 U790 ( .D0(n434), .D1(\spm_in[SDATA][18] ), .S0(n142), .Z(
        n699) );
  HS65_LS_MUX21I1X6 U791 ( .D0(n435), .D1(\spm_in[SDATA][19] ), .S0(n140), .Z(
        n698) );
  HS65_LS_MUX21I1X6 U792 ( .D0(n436), .D1(\spm_in[SDATA][20] ), .S0(n140), .Z(
        n697) );
  HS65_LS_MUX21I1X6 U793 ( .D0(n437), .D1(\spm_in[SDATA][21] ), .S0(n140), .Z(
        n696) );
  HS65_LS_MUX21I1X6 U794 ( .D0(n438), .D1(\spm_in[SDATA][22] ), .S0(n142), .Z(
        n695) );
  HS65_LS_MUX21I1X6 U795 ( .D0(n439), .D1(\spm_in[SDATA][23] ), .S0(n140), .Z(
        n694) );
  HS65_LS_MUX21I1X6 U796 ( .D0(n440), .D1(\spm_in[SDATA][24] ), .S0(n140), .Z(
        n693) );
  HS65_LS_MUX21I1X6 U797 ( .D0(n441), .D1(\spm_in[SDATA][25] ), .S0(n142), .Z(
        n692) );
  HS65_LS_MUX21I1X6 U798 ( .D0(n442), .D1(\spm_in[SDATA][26] ), .S0(n140), .Z(
        n691) );
  HS65_LS_MUX21I1X6 U799 ( .D0(n443), .D1(\spm_in[SDATA][27] ), .S0(n140), .Z(
        n690) );
  HS65_LS_MUX21I1X6 U800 ( .D0(n444), .D1(\spm_in[SDATA][28] ), .S0(n140), .Z(
        n689) );
  HS65_LS_MUX21I1X6 U801 ( .D0(n445), .D1(\spm_in[SDATA][29] ), .S0(n142), .Z(
        n688) );
  HS65_LS_MUX21I1X6 U802 ( .D0(n446), .D1(\spm_in[SDATA][30] ), .S0(n142), .Z(
        n687) );
  HS65_LS_MUX21I1X6 U803 ( .D0(n447), .D1(\spm_in[SDATA][31] ), .S0(n142), .Z(
        n686) );
  HS65_LS_IVX9 U804 ( .A(\phase_next[1] ), .Z(n457) );
  HS65_LS_IVX9 U805 ( .A(n449), .Z(n464) );
  HS65_LS_IVX9 U806 ( .A(n461), .Z(n462) );
  HS65_LS_IVX9 U807 ( .A(phitOut1[0]), .Z(n468) );
  HS65_LS_IVX9 U808 ( .A(phitOut0[0]), .Z(n467) );
  HS65_LS_NAND2X7 U809 ( .A(phitOut2[0]), .B(n45), .Z(n466) );
  HS65_LS_OAI212X5 U810 ( .A(n468), .B(n28), .C(n26), .D(n467), .E(n466), .Z(
        pkt_out[0]) );
  HS65_LS_IVX9 U811 ( .A(phitOut1[1]), .Z(n471) );
  HS65_LS_IVX9 U812 ( .A(phitOut0[1]), .Z(n470) );
  HS65_LS_NAND2X7 U813 ( .A(phitOut2[1]), .B(n45), .Z(n469) );
  HS65_LS_OAI212X5 U814 ( .A(n471), .B(n29), .C(n23), .D(n470), .E(n469), .Z(
        pkt_out[1]) );
  HS65_LS_IVX9 U815 ( .A(phitOut1[2]), .Z(n474) );
  HS65_LS_IVX9 U816 ( .A(phitOut0[2]), .Z(n473) );
  HS65_LS_OAI212X5 U817 ( .A(n474), .B(n28), .C(n23), .D(n473), .E(n472), .Z(
        pkt_out[2]) );
  HS65_LS_IVX9 U818 ( .A(phitOut1[3]), .Z(n479) );
  HS65_LS_IVX9 U819 ( .A(phitOut0[3]), .Z(n478) );
  HS65_LS_OAI212X5 U820 ( .A(n125), .B(n479), .C(n23), .D(n478), .E(n477), .Z(
        pkt_out[3]) );
  HS65_LS_IVX9 U821 ( .A(phitOut1[4]), .Z(n482) );
  HS65_LS_IVX9 U822 ( .A(phitOut0[4]), .Z(n481) );
  HS65_LS_OAI212X5 U823 ( .A(n482), .B(n124), .C(n23), .D(n481), .E(n480), .Z(
        pkt_out[4]) );
  HS65_LS_IVX9 U824 ( .A(phitOut1[5]), .Z(n485) );
  HS65_LS_IVX9 U825 ( .A(phitOut0[5]), .Z(n484) );
  HS65_LS_OAI212X5 U826 ( .A(n485), .B(n29), .C(n23), .D(n484), .E(n483), .Z(
        pkt_out[5]) );
  HS65_LS_IVX9 U827 ( .A(phitOut1[6]), .Z(n488) );
  HS65_LS_IVX9 U828 ( .A(phitOut0[6]), .Z(n487) );
  HS65_LS_OAI212X5 U829 ( .A(n488), .B(n28), .C(n23), .D(n487), .E(n486), .Z(
        pkt_out[6]) );
  HS65_LS_IVX9 U830 ( .A(phitOut1[7]), .Z(n491) );
  HS65_LS_IVX9 U831 ( .A(phitOut0[7]), .Z(n490) );
  HS65_LS_OAI212X5 U832 ( .A(n491), .B(n28), .C(n23), .D(n490), .E(n489), .Z(
        pkt_out[7]) );
  HS65_LS_IVX9 U833 ( .A(phitOut1[8]), .Z(n494) );
  HS65_LS_IVX9 U834 ( .A(phitOut0[8]), .Z(n493) );
  HS65_LS_IVX9 U835 ( .A(phitOut1[9]), .Z(n497) );
  HS65_LS_IVX9 U836 ( .A(phitOut0[9]), .Z(n496) );
  HS65_LS_OAI212X5 U837 ( .A(n497), .B(n29), .C(n496), .D(n23), .E(n495), .Z(
        pkt_out[9]) );
  HS65_LS_IVX9 U838 ( .A(phitOut1[10]), .Z(n500) );
  HS65_LS_IVX9 U839 ( .A(phitOut0[10]), .Z(n499) );
  HS65_LS_IVX9 U840 ( .A(phitOut1[11]), .Z(n503) );
  HS65_LS_IVX9 U841 ( .A(phitOut0[11]), .Z(n502) );
  HS65_LS_OAI212X5 U842 ( .A(n503), .B(n28), .C(n23), .D(n502), .E(n501), .Z(
        pkt_out[11]) );
  HS65_LS_IVX9 U843 ( .A(phitOut1[12]), .Z(n506) );
  HS65_LS_IVX9 U844 ( .A(phitOut0[12]), .Z(n505) );
  HS65_LS_OAI212X5 U845 ( .A(n506), .B(n28), .C(n23), .D(n505), .E(n504), .Z(
        pkt_out[12]) );
  HS65_LS_IVX9 U846 ( .A(phitOut1[13]), .Z(n509) );
  HS65_LS_IVX9 U847 ( .A(phitOut0[13]), .Z(n508) );
  HS65_LS_OAI212X5 U848 ( .A(n509), .B(n124), .C(n23), .D(n508), .E(n507), .Z(
        pkt_out[13]) );
  HS65_LS_IVX9 U849 ( .A(phitOut1[14]), .Z(n512) );
  HS65_LS_IVX9 U850 ( .A(phitOut0[14]), .Z(n511) );
  HS65_LS_OAI212X5 U851 ( .A(n512), .B(n43), .C(n23), .D(n511), .E(n510), .Z(
        pkt_out[14]) );
  HS65_LS_IVX9 U852 ( .A(phitOut1[15]), .Z(n516) );
  HS65_LS_IVX9 U853 ( .A(phitOut0[15]), .Z(n515) );
  HS65_LS_OAI212X5 U854 ( .A(n516), .B(n29), .C(n23), .D(n515), .E(n514), .Z(
        pkt_out[15]) );
  HS65_LS_IVX9 U855 ( .A(phitOut1[16]), .Z(n519) );
  HS65_LS_IVX9 U856 ( .A(phitOut0[16]), .Z(n518) );
  HS65_LS_OAI212X5 U857 ( .A(n519), .B(n29), .C(n518), .D(n23), .E(n517), .Z(
        pkt_out[16]) );
  HS65_LS_IVX9 U858 ( .A(phitOut1[17]), .Z(n522) );
  HS65_LS_IVX9 U859 ( .A(phitOut0[17]), .Z(n521) );
  HS65_LS_IVX9 U860 ( .A(phitOut1[18]), .Z(n525) );
  HS65_LS_IVX9 U861 ( .A(phitOut0[18]), .Z(n524) );
  HS65_LS_OAI212X5 U862 ( .A(n525), .B(n43), .C(n524), .D(n23), .E(n523), .Z(
        pkt_out[18]) );
  HS65_LS_IVX9 U863 ( .A(phitOut1[19]), .Z(n528) );
  HS65_LS_IVX9 U864 ( .A(phitOut0[19]), .Z(n527) );
  HS65_LS_IVX9 U865 ( .A(phitOut1[20]), .Z(n531) );
  HS65_LS_IVX9 U866 ( .A(phitOut0[20]), .Z(n530) );
  HS65_LS_OAI212X5 U867 ( .A(n531), .B(n124), .C(n31), .D(n530), .E(n529), .Z(
        pkt_out[20]) );
  HS65_LS_IVX9 U868 ( .A(phitOut1[21]), .Z(n534) );
  HS65_LS_IVX9 U869 ( .A(phitOut0[21]), .Z(n533) );
  HS65_LS_OAI212X5 U870 ( .A(n534), .B(n28), .C(n31), .D(n533), .E(n532), .Z(
        pkt_out[21]) );
  HS65_LS_IVX9 U871 ( .A(phitOut1[22]), .Z(n537) );
  HS65_LS_IVX9 U872 ( .A(phitOut0[22]), .Z(n536) );
  HS65_LS_IVX9 U873 ( .A(phitOut1[23]), .Z(n540) );
  HS65_LS_IVX9 U874 ( .A(phitOut0[23]), .Z(n539) );
  HS65_LS_OAI212X5 U875 ( .A(n540), .B(n124), .C(n31), .D(n539), .E(n538), .Z(
        pkt_out[23]) );
  HS65_LS_IVX9 U876 ( .A(phitOut1[24]), .Z(n543) );
  HS65_LS_IVX9 U877 ( .A(phitOut0[24]), .Z(n542) );
  HS65_LS_OAI212X5 U878 ( .A(n543), .B(n124), .C(n31), .D(n542), .E(n541), .Z(
        pkt_out[24]) );
  HS65_LS_IVX9 U879 ( .A(phitOut1[25]), .Z(n546) );
  HS65_LS_IVX9 U880 ( .A(phitOut0[25]), .Z(n545) );
  HS65_LS_OAI212X5 U881 ( .A(n546), .B(n43), .C(n31), .D(n545), .E(n544), .Z(
        pkt_out[25]) );
  HS65_LS_IVX9 U882 ( .A(phitOut1[26]), .Z(n549) );
  HS65_LS_IVX9 U883 ( .A(phitOut0[26]), .Z(n548) );
  HS65_LS_OAI212X5 U884 ( .A(n549), .B(n29), .C(n31), .D(n548), .E(n547), .Z(
        pkt_out[26]) );
  HS65_LS_IVX9 U885 ( .A(phitOut1[27]), .Z(n552) );
  HS65_LS_IVX9 U886 ( .A(phitOut0[27]), .Z(n551) );
  HS65_LS_IVX9 U887 ( .A(phitOut1[28]), .Z(n555) );
  HS65_LS_IVX9 U888 ( .A(phitOut0[28]), .Z(n554) );
  HS65_LS_OAI212X5 U889 ( .A(n555), .B(n125), .C(n31), .D(n554), .E(n553), .Z(
        pkt_out[28]) );
  HS65_LS_IVX9 U890 ( .A(phitOut1[29]), .Z(n558) );
  HS65_LS_IVX9 U891 ( .A(phitOut0[29]), .Z(n557) );
  HS65_LS_OAI212X5 U892 ( .A(n558), .B(n29), .C(n31), .D(n557), .E(n556), .Z(
        pkt_out[29]) );
  HS65_LS_IVX9 U893 ( .A(phitOut1[30]), .Z(n561) );
  HS65_LS_IVX9 U894 ( .A(phitOut0[30]), .Z(n560) );
  HS65_LS_IVX9 U895 ( .A(phitOut1[31]), .Z(n564) );
  HS65_LS_IVX9 U896 ( .A(phitOut0[31]), .Z(n563) );
  HS65_LS_OAI212X5 U897 ( .A(n564), .B(n28), .C(n31), .D(n563), .E(n562), .Z(
        pkt_out[31]) );
  HS65_LS_IVX9 U898 ( .A(phitOut1[32]), .Z(n567) );
  HS65_LS_IVX9 U899 ( .A(phitOut0[32]), .Z(n566) );
  HS65_LS_OAI212X5 U900 ( .A(n567), .B(n29), .C(n31), .D(n566), .E(n565), .Z(
        pkt_out[32]) );
  HS65_LS_IVX9 U901 ( .A(phitOut1[33]), .Z(n571) );
  HS65_LS_IVX9 U902 ( .A(phitOut0[33]), .Z(n569) );
  HS65_LS_IVX9 U903 ( .A(phitOut1[34]), .Z(n574) );
  HS65_LS_IVX9 U904 ( .A(flit_buf[64]), .Z(n577) );
  HS65_LS_OAI22X6 U905 ( .A(n359), .B(n578), .C(n591), .D(n577), .Z(
        \spm_out[MADDR][0] ) );
  HS65_LS_IVX9 U906 ( .A(flit_buf[65]), .Z(n579) );
  HS65_LS_OAI22X6 U907 ( .A(n359), .B(n580), .C(n591), .D(n579), .Z(
        \spm_out[MADDR][1] ) );
  HS65_LS_IVX9 U908 ( .A(flit_buf[66]), .Z(n581) );
  HS65_LS_OAI22X6 U909 ( .A(n359), .B(n582), .C(n591), .D(n581), .Z(
        \spm_out[MADDR][2] ) );
  HS65_LS_IVX9 U910 ( .A(flit_buf[67]), .Z(n583) );
  HS65_LS_OAI22X6 U911 ( .A(n359), .B(n584), .C(n591), .D(n583), .Z(
        \spm_out[MADDR][3] ) );
  HS65_LS_IVX9 U912 ( .A(flit_buf[68]), .Z(n585) );
  HS65_LS_OAI22X6 U913 ( .A(n359), .B(n586), .C(n591), .D(n585), .Z(
        \spm_out[MADDR][4] ) );
  HS65_LS_IVX9 U914 ( .A(flit_buf[69]), .Z(n587) );
  HS65_LS_OAI22X6 U915 ( .A(n359), .B(n588), .C(n591), .D(n587), .Z(
        \spm_out[MADDR][5] ) );
  HS65_LS_IVX9 U916 ( .A(flit_buf[70]), .Z(n589) );
  HS65_LS_OAI22X6 U917 ( .A(n590), .B(n359), .C(n591), .D(n589), .Z(
        \spm_out[MADDR][6] ) );
  HS65_LS_IVX9 U918 ( .A(n591), .Z(\spm_out[MCMD][0] ) );
  HS65_LS_IVX9 U919 ( .A(n592), .Z(n594) );
  HS65_LS_OAI112X5 U920 ( .A(n867), .B(n594), .C(n866), .D(n593), .Z(
        \proc_out[SCMDACCEPT] ) );
endmodule


module latch_controller_1_25 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_25 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n3, n4, n5, n6;
  assign N0 = preset;

  latch_controller_1_25 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n4), .RN(n3), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n3), .Z(n5) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n6), .B(n5), .Z(N5) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_IVX9 U3 ( .A(lt_enable), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(N0), .Z(n3) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n4), .Z(lt_gated) );
endmodule


module latch_controller_1_24 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_24 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n3, n4, n5, n6;
  assign N0 = preset;

  latch_controller_1_24 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n4), .RN(n3), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n3), .Z(n5) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n6), .B(n5), .Z(N5) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_IVX9 U3 ( .A(lt_enable), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(N0), .Z(n3) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n4), .Z(lt_gated) );
endmodule


module latch_controller_1_23 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_23 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n3, n4, n5, n6;
  assign N0 = preset;

  latch_controller_1_23 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n4), .RN(n3), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n3), .Z(n5) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n6), .B(n5), .Z(N5) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_IVX9 U3 ( .A(lt_enable), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(N0), .Z(n3) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n4), .Z(lt_gated) );
endmodule


module latch_controller_1_22 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_22 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n3, n4, n5, n6;
  assign N0 = preset;

  latch_controller_1_22 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n4), .RN(n3), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n3), .Z(n5) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n6), .B(n5), .Z(N5) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_IVX9 U3 ( .A(lt_enable), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(N0), .Z(n3) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n4), .Z(lt_gated) );
endmodule


module latch_controller_1_21 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_NOR2AX3 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_21 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n3, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_21 controller ( .preset(n3), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLRQX18 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(n3), .Z(n7) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_LDHQX4 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX4 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX18 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX18 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX18 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX18 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX18 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX18 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX18 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX18 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX18 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX18 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX18 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX18 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX18 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX18 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX18 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX18 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX18 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX4 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX4 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX18 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX18 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX18 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX18 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX18 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX18 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX18 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX18 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX18 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX18 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX18 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX18 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX18 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_IVX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_IVX9 U5 ( .A(N0), .Z(n4) );
  HS65_LS_NAND2X7 U9 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_comb_0_0_1 ( data_valid, data_in, preset, data_out, sel );
  input [34:0] data_in;
  output [34:0] data_out;
  output [4:0] sel;
  input data_valid, preset;
  wire   data_in_34, data_in_33, data_in_32, \data_in[31] , \data_in[30] ,
         \data_in[29] , \data_in[28] , \data_in[27] , \data_in[26] ,
         \data_in[25] , \data_in[24] , \data_in[23] , \data_in[22] ,
         \data_in[21] , \data_in[20] , \data_in[19] , \data_in[18] ,
         \data_in[17] , \data_in[16] , N23, N25, N26, N27, N28, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n22,
         n23, n24;
  assign data_out[34] = data_in_34;
  assign data_in_34 = data_in[34];
  assign data_out[33] = data_in_33;
  assign data_in_33 = data_in[33];
  assign data_out[32] = data_in_32;
  assign data_in_32 = data_in[32];
  assign data_out[31] = \data_in[31] ;
  assign \data_in[31]  = data_in[31];
  assign data_out[30] = \data_in[30] ;
  assign \data_in[30]  = data_in[30];
  assign data_out[29] = \data_in[29] ;
  assign \data_in[29]  = data_in[29];
  assign data_out[28] = \data_in[28] ;
  assign \data_in[28]  = data_in[28];
  assign data_out[27] = \data_in[27] ;
  assign \data_in[27]  = data_in[27];
  assign data_out[26] = \data_in[26] ;
  assign \data_in[26]  = data_in[26];
  assign data_out[25] = \data_in[25] ;
  assign \data_in[25]  = data_in[25];
  assign data_out[24] = \data_in[24] ;
  assign \data_in[24]  = data_in[24];
  assign data_out[23] = \data_in[23] ;
  assign \data_in[23]  = data_in[23];
  assign data_out[22] = \data_in[22] ;
  assign \data_in[22]  = data_in[22];
  assign data_out[21] = \data_in[21] ;
  assign \data_in[21]  = data_in[21];
  assign data_out[20] = \data_in[20] ;
  assign \data_in[20]  = data_in[20];
  assign data_out[19] = \data_in[19] ;
  assign \data_in[19]  = data_in[19];
  assign data_out[18] = \data_in[18] ;
  assign \data_in[18]  = data_in[18];
  assign data_out[17] = \data_in[17] ;
  assign \data_in[17]  = data_in[17];
  assign data_out[16] = \data_in[16] ;
  assign \data_in[16]  = data_in[16];
  assign sel[0] = 1'b0;

  HS65_LS_LDHQX9 \sel_reg[4]  ( .G(N23), .D(N28), .Q(sel[4]) );
  HS65_LS_LDHQX9 \sel_reg[3]  ( .G(N23), .D(N27), .Q(sel[3]) );
  HS65_LS_LDHQX9 \sel_reg[2]  ( .G(N23), .D(N26), .Q(sel[2]) );
  HS65_LS_LDHQX9 \sel_reg[1]  ( .G(N23), .D(N25), .Q(sel[1]) );
  HS65_LS_NAND3AX6 U4 ( .A(preset), .B(n23), .C(n2), .Z(n22) );
  HS65_LS_OAI22X6 U5 ( .A(n9), .B(n24), .C(n2), .D(n11), .Z(data_out[7]) );
  HS65_LS_OAI22X6 U6 ( .A(n24), .B(n16), .C(n2), .D(n18), .Z(data_out[0]) );
  HS65_LS_OAI22X6 U7 ( .A(n24), .B(n15), .C(n2), .D(n17), .Z(data_out[1]) );
  HS65_LS_OAI22X6 U8 ( .A(n24), .B(n14), .C(n2), .D(n16), .Z(data_out[2]) );
  HS65_LS_OAI22X6 U9 ( .A(n24), .B(n13), .C(n2), .D(n15), .Z(data_out[3]) );
  HS65_LS_OAI22X6 U10 ( .A(n24), .B(n12), .C(n2), .D(n14), .Z(data_out[4]) );
  HS65_LS_OAI22X6 U11 ( .A(n24), .B(n11), .C(n2), .D(n13), .Z(data_out[5]) );
  HS65_LS_OAI22X6 U12 ( .A(n24), .B(n10), .C(n2), .D(n12), .Z(data_out[6]) );
  HS65_LS_OAI22X6 U13 ( .A(n24), .B(n8), .C(n2), .D(n10), .Z(data_out[8]) );
  HS65_LS_OAI22X6 U14 ( .A(n24), .B(n7), .C(n2), .D(n9), .Z(data_out[9]) );
  HS65_LS_OAI22X6 U15 ( .A(n24), .B(n6), .C(n2), .D(n8), .Z(data_out[10]) );
  HS65_LS_OAI22X6 U16 ( .A(n24), .B(n5), .C(n2), .D(n7), .Z(data_out[11]) );
  HS65_LS_OAI22X6 U17 ( .A(n24), .B(n4), .C(n2), .D(n6), .Z(data_out[12]) );
  HS65_LS_OAI22X6 U18 ( .A(n24), .B(n3), .C(n2), .D(n5), .Z(data_out[13]) );
  HS65_LS_IVX9 U19 ( .A(n24), .Z(n2) );
  HS65_LS_NOR3X4 U20 ( .A(n23), .B(preset), .C(n24), .Z(N28) );
  HS65_LS_NOR3X4 U21 ( .A(n22), .B(n17), .C(n18), .Z(N27) );
  HS65_LS_NAND2X7 U22 ( .A(n17), .B(n18), .Z(n23) );
  HS65_LS_NOR2X6 U23 ( .A(n2), .B(n4), .Z(data_out[14]) );
  HS65_LS_NOR2X6 U24 ( .A(n2), .B(n3), .Z(data_out[15]) );
  HS65_LS_NAND2X14 U25 ( .A(data_in_34), .B(data_in_33), .Z(n24) );
  HS65_LS_IVX9 U26 ( .A(data_in[1]), .Z(n17) );
  HS65_LS_IVX9 U27 ( .A(data_in[0]), .Z(n18) );
  HS65_LS_NOR2X6 U28 ( .A(data_in[1]), .B(n22), .Z(N25) );
  HS65_LS_NOR2X6 U29 ( .A(data_in[0]), .B(n22), .Z(N26) );
  HS65_LS_IVX9 U30 ( .A(data_in[9]), .Z(n9) );
  HS65_LS_IVX9 U31 ( .A(data_in[2]), .Z(n16) );
  HS65_LS_IVX9 U32 ( .A(data_in[3]), .Z(n15) );
  HS65_LS_IVX9 U33 ( .A(data_in[4]), .Z(n14) );
  HS65_LS_IVX9 U34 ( .A(data_in[5]), .Z(n13) );
  HS65_LS_IVX9 U35 ( .A(data_in[6]), .Z(n12) );
  HS65_LS_IVX9 U36 ( .A(data_in[7]), .Z(n11) );
  HS65_LS_IVX9 U37 ( .A(data_in[8]), .Z(n10) );
  HS65_LS_IVX9 U38 ( .A(data_in[10]), .Z(n8) );
  HS65_LS_IVX9 U39 ( .A(data_in[11]), .Z(n7) );
  HS65_LS_IVX9 U40 ( .A(data_in[12]), .Z(n6) );
  HS65_LS_IVX9 U41 ( .A(data_in[13]), .Z(n5) );
  HS65_LS_IVX9 U42 ( .A(data_in[14]), .Z(n4) );
  HS65_LS_IVX9 U43 ( .A(data_in[15]), .Z(n3) );
  HS65_LS_CB4I6X9 U44 ( .A(n2), .B(n1), .C(data_valid), .D(preset), .Z(N23) );
  HS65_LS_IVX9 U45 ( .A(data_in_34), .Z(n1) );
endmodule


module latch_controller_1_5 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_5 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_5 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n7) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_IVX9 U3 ( .A(N0), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_0_0_1 ( preset, .chan_in_f({\chan_in_f[REQ] , \chan_in_f[DATA][34] , 
        \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , 
        \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , 
        \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , 
        \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , 
        \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , 
        \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , 
        \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , 
        \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , 
        \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , 
        \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , 
        \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , 
        \chan_in_f[DATA][0] }), .chan_in_b(\chan_in_b[ACK] ), .chan_out_f({
        \chan_out_f[REQ] , \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , 
        \chan_out_f[DATA][32] , \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , 
        \chan_out_f[DATA][29] , \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , 
        \chan_out_f[DATA][26] , \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , 
        \chan_out_f[DATA][23] , \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , 
        \chan_out_f[DATA][20] , \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , 
        \chan_out_f[DATA][17] , \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , 
        \chan_out_f[DATA][14] , \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , 
        \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , 
        \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , 
        \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , 
        \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), 
    .chan_out_b(\chan_out_b[ACK] ), sel );
  output [4:0] sel;
  input preset, \chan_in_f[REQ] , \chan_in_f[DATA][34] , \chan_in_f[DATA][33] ,
         \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , \chan_in_f[DATA][30] ,
         \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , \chan_in_f[DATA][27] ,
         \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , \chan_in_f[DATA][24] ,
         \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , \chan_in_f[DATA][21] ,
         \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , \chan_in_f[DATA][18] ,
         \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , \chan_in_f[DATA][15] ,
         \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , \chan_in_f[DATA][12] ,
         \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , \chan_in_f[DATA][9] ,
         \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , \chan_in_f[DATA][6] ,
         \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , \chan_in_f[DATA][3] ,
         \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , \chan_in_f[DATA][0] ,
         \chan_out_b[ACK] ;
  output \chan_in_b[ACK] , \chan_out_f[REQ] , \chan_out_f[DATA][34] ,
         \chan_out_f[DATA][33] , \chan_out_f[DATA][32] ,
         \chan_out_f[DATA][31] , \chan_out_f[DATA][30] ,
         \chan_out_f[DATA][29] , \chan_out_f[DATA][28] ,
         \chan_out_f[DATA][27] , \chan_out_f[DATA][26] ,
         \chan_out_f[DATA][25] , \chan_out_f[DATA][24] ,
         \chan_out_f[DATA][23] , \chan_out_f[DATA][22] ,
         \chan_out_f[DATA][21] , \chan_out_f[DATA][20] ,
         \chan_out_f[DATA][19] , \chan_out_f[DATA][18] ,
         \chan_out_f[DATA][17] , \chan_out_f[DATA][16] ,
         \chan_out_f[DATA][15] , \chan_out_f[DATA][14] ,
         \chan_out_f[DATA][13] , \chan_out_f[DATA][12] ,
         \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] ,
         \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] ,
         \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] ,
         \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] ;
  wire   \chan_internal_f[REQ] , \chan_internal_f[DATA][34] ,
         \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] ,
         \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] ,
         \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] ,
         \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] ,
         \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] ,
         \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] ,
         \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] ,
         \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] ,
         \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] ,
         \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] ,
         \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] ,
         \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] ,
         \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] ,
         \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] ,
         \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] ,
         \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] ,
         \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] , req_n, lt_en,
         n1, n2, n3, n4, n5, n6, n7;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign sel[0] = 1'b0;

  hpu_comb_0_0_1 hpu_combinatorial ( .data_valid(lt_en), .data_in({
        \chan_in_f[DATA][34] , \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , 
        \chan_in_f[DATA][31] , \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , 
        \chan_in_f[DATA][28] , \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , 
        \chan_in_f[DATA][25] , \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , 
        \chan_in_f[DATA][22] , \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , 
        \chan_in_f[DATA][19] , \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , 
        \chan_in_f[DATA][16] , \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , 
        \chan_in_f[DATA][13] , \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , 
        \chan_in_f[DATA][10] , \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , 
        \chan_in_f[DATA][7] , \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , 
        \chan_in_f[DATA][4] , \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , 
        \chan_in_f[DATA][1] , \chan_in_f[DATA][0] }), .preset(n7), .data_out({
        \chan_internal_f[DATA][34] , \chan_internal_f[DATA][33] , 
        \chan_internal_f[DATA][32] , \chan_internal_f[DATA][31] , 
        \chan_internal_f[DATA][30] , \chan_internal_f[DATA][29] , 
        \chan_internal_f[DATA][28] , \chan_internal_f[DATA][27] , 
        \chan_internal_f[DATA][26] , \chan_internal_f[DATA][25] , 
        \chan_internal_f[DATA][24] , \chan_internal_f[DATA][23] , 
        \chan_internal_f[DATA][22] , \chan_internal_f[DATA][21] , 
        \chan_internal_f[DATA][20] , \chan_internal_f[DATA][19] , 
        \chan_internal_f[DATA][18] , \chan_internal_f[DATA][17] , 
        \chan_internal_f[DATA][16] , \chan_internal_f[DATA][15] , 
        \chan_internal_f[DATA][14] , \chan_internal_f[DATA][13] , 
        \chan_internal_f[DATA][12] , \chan_internal_f[DATA][11] , 
        \chan_internal_f[DATA][10] , \chan_internal_f[DATA][9] , 
        \chan_internal_f[DATA][8] , \chan_internal_f[DATA][7] , 
        \chan_internal_f[DATA][6] , \chan_internal_f[DATA][5] , 
        \chan_internal_f[DATA][4] , \chan_internal_f[DATA][3] , 
        \chan_internal_f[DATA][2] , \chan_internal_f[DATA][1] , 
        \chan_internal_f[DATA][0] }), .sel({sel[4:1], SYNOPSYS_UNCONNECTED__0}) );
  channel_latch_1_xxxxxxxxx_5 token_latch ( .preset(n7), .left_in({
        \chan_internal_f[REQ] , \chan_internal_f[DATA][34] , 
        \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] , 
        \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] , 
        \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] , 
        \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] , 
        \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] , 
        \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] , 
        \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] , 
        \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] , 
        \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] , 
        \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] , 
        \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] , 
        \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] , 
        \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] , 
        \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] , 
        \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] , 
        \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] , 
        \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] }), .left_out(
        \chan_in_b[ACK] ), .right_out({\chan_out_f[REQ] , 
        \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , \chan_out_f[DATA][32] , 
        \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , \chan_out_f[DATA][29] , 
        \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , \chan_out_f[DATA][26] , 
        \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , \chan_out_f[DATA][23] , 
        \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , \chan_out_f[DATA][20] , 
        \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , \chan_out_f[DATA][17] , 
        \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , \chan_out_f[DATA][14] , 
        \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , \chan_out_f[DATA][11] , 
        \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , \chan_out_f[DATA][8] , 
        \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , \chan_out_f[DATA][5] , 
        \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , \chan_out_f[DATA][2] , 
        \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), .right_in(
        \chan_out_b[ACK] ), .lt_enable(lt_en) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chan_internal_f[REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(\chan_in_f[REQ] ), .Z(req_n) );
  HS65_LS_BFX9 U1 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U2 ( .A(n3), .Z(n2) );
  HS65_LS_BFX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_BFX9 U4 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U6 ( .A(req_n), .Z(n6) );
  HS65_LS_BFX9 U7 ( .A(preset), .Z(n7) );
endmodule


module hpu_comb_0_2_1 ( data_valid, data_in, preset, data_out, sel );
  input [34:0] data_in;
  output [34:0] data_out;
  output [4:0] sel;
  input data_valid, preset;
  wire   data_in_34, data_in_33, data_in_32, \data_in[31] , \data_in[30] ,
         \data_in[29] , \data_in[28] , \data_in[27] , \data_in[26] ,
         \data_in[25] , \data_in[24] , \data_in[23] , \data_in[22] ,
         \data_in[21] , \data_in[20] , \data_in[19] , \data_in[18] ,
         \data_in[17] , \data_in[16] , N26, N27, N28, N30, N31, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n15, n16, n17, n18;
  assign data_out[34] = data_in_34;
  assign data_in_34 = data_in[34];
  assign data_out[33] = data_in_33;
  assign data_in_33 = data_in[33];
  assign data_out[32] = data_in_32;
  assign data_in_32 = data_in[32];
  assign data_out[31] = \data_in[31] ;
  assign \data_in[31]  = data_in[31];
  assign data_out[30] = \data_in[30] ;
  assign \data_in[30]  = data_in[30];
  assign data_out[29] = \data_in[29] ;
  assign \data_in[29]  = data_in[29];
  assign data_out[28] = \data_in[28] ;
  assign \data_in[28]  = data_in[28];
  assign data_out[27] = \data_in[27] ;
  assign \data_in[27]  = data_in[27];
  assign data_out[26] = \data_in[26] ;
  assign \data_in[26]  = data_in[26];
  assign data_out[25] = \data_in[25] ;
  assign \data_in[25]  = data_in[25];
  assign data_out[24] = \data_in[24] ;
  assign \data_in[24]  = data_in[24];
  assign data_out[23] = \data_in[23] ;
  assign \data_in[23]  = data_in[23];
  assign data_out[22] = \data_in[22] ;
  assign \data_in[22]  = data_in[22];
  assign data_out[21] = \data_in[21] ;
  assign \data_in[21]  = data_in[21];
  assign data_out[20] = \data_in[20] ;
  assign \data_in[20]  = data_in[20];
  assign data_out[19] = \data_in[19] ;
  assign \data_in[19]  = data_in[19];
  assign data_out[18] = \data_in[18] ;
  assign \data_in[18]  = data_in[18];
  assign data_out[17] = \data_in[17] ;
  assign \data_in[17]  = data_in[17];
  assign data_out[16] = \data_in[16] ;
  assign \data_in[16]  = data_in[16];
  assign sel[2] = 1'b0;

  HS65_LS_LDHQX9 \sel_reg[4]  ( .G(N26), .D(N31), .Q(sel[4]) );
  HS65_LS_LDHQX9 \sel_reg[3]  ( .G(N26), .D(N30), .Q(sel[3]) );
  HS65_LS_LDHQX9 \sel_reg[1]  ( .G(N26), .D(N28), .Q(sel[1]) );
  HS65_LS_LDHQX9 \sel_reg[0]  ( .G(N26), .D(N27), .Q(sel[0]) );
  HS65_LS_OAI22X6 U4 ( .A(n18), .B(n9), .C(n2), .D(n10), .Z(data_out[0]) );
  HS65_LS_OAI22X6 U5 ( .A(n18), .B(n8), .C(n2), .D(n9), .Z(data_out[2]) );
  HS65_LS_OAI22X6 U6 ( .A(n18), .B(n7), .C(n2), .D(n8), .Z(data_out[4]) );
  HS65_LS_OAI22X6 U7 ( .A(n18), .B(n6), .C(n2), .D(n7), .Z(data_out[6]) );
  HS65_LS_OAI22X6 U8 ( .A(n18), .B(n5), .C(n2), .D(n6), .Z(data_out[8]) );
  HS65_LS_OAI22X6 U9 ( .A(n18), .B(n4), .C(n2), .D(n5), .Z(data_out[10]) );
  HS65_LS_OAI22X6 U10 ( .A(n18), .B(n3), .C(n2), .D(n4), .Z(data_out[12]) );
  HS65_LS_NAND3AX6 U11 ( .A(preset), .B(n17), .C(n2), .Z(n16) );
  HS65_LS_NOR3X4 U12 ( .A(n17), .B(preset), .C(n18), .Z(N31) );
  HS65_LS_IVX9 U13 ( .A(n18), .Z(n2) );
  HS65_LS_NOR3X4 U14 ( .A(n16), .B(n10), .C(n15), .Z(N30) );
  HS65_LS_NOR2AX3 U15 ( .A(n15), .B(n16), .Z(N28) );
  HS65_LS_NOR2X6 U16 ( .A(n2), .B(n3), .Z(data_out[14]) );
  HS65_LS_NAND2X14 U17 ( .A(data_in_34), .B(data_in_33), .Z(n18) );
  HS65_LS_IVX9 U18 ( .A(data_in[0]), .Z(n10) );
  HS65_LS_NAND2X7 U19 ( .A(data_in[1]), .B(n10), .Z(n17) );
  HS65_LS_NOR2X6 U20 ( .A(n10), .B(data_in[1]), .Z(n15) );
  HS65_LS_NOR2X6 U21 ( .A(data_in[0]), .B(n16), .Z(N27) );
  HS65_LS_IVX9 U22 ( .A(data_in[2]), .Z(n9) );
  HS65_LS_IVX9 U23 ( .A(data_in[4]), .Z(n8) );
  HS65_LS_IVX9 U24 ( .A(data_in[6]), .Z(n7) );
  HS65_LS_IVX9 U25 ( .A(data_in[8]), .Z(n6) );
  HS65_LS_IVX9 U26 ( .A(data_in[10]), .Z(n5) );
  HS65_LS_IVX9 U27 ( .A(data_in[12]), .Z(n4) );
  HS65_LS_IVX9 U28 ( .A(data_in[14]), .Z(n3) );
  HS65_LS_AO22X9 U29 ( .A(n2), .B(data_in[3]), .C(n18), .D(data_in[1]), .Z(
        data_out[1]) );
  HS65_LS_AO22X9 U30 ( .A(n2), .B(data_in[5]), .C(n18), .D(data_in[3]), .Z(
        data_out[3]) );
  HS65_LS_AO22X9 U31 ( .A(n2), .B(data_in[7]), .C(n18), .D(data_in[5]), .Z(
        data_out[5]) );
  HS65_LS_AO22X9 U32 ( .A(data_in[9]), .B(n2), .C(n18), .D(data_in[7]), .Z(
        data_out[7]) );
  HS65_LS_AO22X9 U33 ( .A(n2), .B(data_in[11]), .C(n18), .D(data_in[9]), .Z(
        data_out[9]) );
  HS65_LS_AO22X9 U34 ( .A(n2), .B(data_in[13]), .C(n18), .D(data_in[11]), .Z(
        data_out[11]) );
  HS65_LS_AO22X9 U35 ( .A(n2), .B(data_in[15]), .C(n18), .D(data_in[13]), .Z(
        data_out[13]) );
  HS65_LS_AND2X4 U36 ( .A(data_in[15]), .B(n18), .Z(data_out[15]) );
  HS65_LS_CB4I6X9 U37 ( .A(n2), .B(n1), .C(data_valid), .D(preset), .Z(N26) );
  HS65_LS_IVX9 U38 ( .A(data_in_34), .Z(n1) );
endmodule


module latch_controller_1_4 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_4 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_4 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n7) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_IVX9 U3 ( .A(N0), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_0_2_1 ( preset, .chan_in_f({\chan_in_f[REQ] , \chan_in_f[DATA][34] , 
        \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , 
        \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , 
        \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , 
        \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , 
        \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , 
        \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , 
        \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , 
        \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , 
        \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , 
        \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , 
        \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , 
        \chan_in_f[DATA][0] }), .chan_in_b(\chan_in_b[ACK] ), .chan_out_f({
        \chan_out_f[REQ] , \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , 
        \chan_out_f[DATA][32] , \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , 
        \chan_out_f[DATA][29] , \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , 
        \chan_out_f[DATA][26] , \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , 
        \chan_out_f[DATA][23] , \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , 
        \chan_out_f[DATA][20] , \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , 
        \chan_out_f[DATA][17] , \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , 
        \chan_out_f[DATA][14] , \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , 
        \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , 
        \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , 
        \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , 
        \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), 
    .chan_out_b(\chan_out_b[ACK] ), sel );
  output [4:0] sel;
  input preset, \chan_in_f[REQ] , \chan_in_f[DATA][34] , \chan_in_f[DATA][33] ,
         \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , \chan_in_f[DATA][30] ,
         \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , \chan_in_f[DATA][27] ,
         \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , \chan_in_f[DATA][24] ,
         \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , \chan_in_f[DATA][21] ,
         \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , \chan_in_f[DATA][18] ,
         \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , \chan_in_f[DATA][15] ,
         \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , \chan_in_f[DATA][12] ,
         \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , \chan_in_f[DATA][9] ,
         \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , \chan_in_f[DATA][6] ,
         \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , \chan_in_f[DATA][3] ,
         \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , \chan_in_f[DATA][0] ,
         \chan_out_b[ACK] ;
  output \chan_in_b[ACK] , \chan_out_f[REQ] , \chan_out_f[DATA][34] ,
         \chan_out_f[DATA][33] , \chan_out_f[DATA][32] ,
         \chan_out_f[DATA][31] , \chan_out_f[DATA][30] ,
         \chan_out_f[DATA][29] , \chan_out_f[DATA][28] ,
         \chan_out_f[DATA][27] , \chan_out_f[DATA][26] ,
         \chan_out_f[DATA][25] , \chan_out_f[DATA][24] ,
         \chan_out_f[DATA][23] , \chan_out_f[DATA][22] ,
         \chan_out_f[DATA][21] , \chan_out_f[DATA][20] ,
         \chan_out_f[DATA][19] , \chan_out_f[DATA][18] ,
         \chan_out_f[DATA][17] , \chan_out_f[DATA][16] ,
         \chan_out_f[DATA][15] , \chan_out_f[DATA][14] ,
         \chan_out_f[DATA][13] , \chan_out_f[DATA][12] ,
         \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] ,
         \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] ,
         \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] ,
         \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] ;
  wire   \chan_internal_f[REQ] , \chan_internal_f[DATA][34] ,
         \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] ,
         \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] ,
         \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] ,
         \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] ,
         \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] ,
         \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] ,
         \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] ,
         \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] ,
         \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] ,
         \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] ,
         \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] ,
         \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] ,
         \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] ,
         \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] ,
         \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] ,
         \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] ,
         \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] , req_n, lt_en,
         n1, n2, n3, n4, n5, n6, n7;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign sel[2] = 1'b0;

  hpu_comb_0_2_1 hpu_combinatorial ( .data_valid(lt_en), .data_in({
        \chan_in_f[DATA][34] , \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , 
        \chan_in_f[DATA][31] , \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , 
        \chan_in_f[DATA][28] , \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , 
        \chan_in_f[DATA][25] , \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , 
        \chan_in_f[DATA][22] , \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , 
        \chan_in_f[DATA][19] , \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , 
        \chan_in_f[DATA][16] , \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , 
        \chan_in_f[DATA][13] , \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , 
        \chan_in_f[DATA][10] , \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , 
        \chan_in_f[DATA][7] , \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , 
        \chan_in_f[DATA][4] , \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , 
        \chan_in_f[DATA][1] , \chan_in_f[DATA][0] }), .preset(n7), .data_out({
        \chan_internal_f[DATA][34] , \chan_internal_f[DATA][33] , 
        \chan_internal_f[DATA][32] , \chan_internal_f[DATA][31] , 
        \chan_internal_f[DATA][30] , \chan_internal_f[DATA][29] , 
        \chan_internal_f[DATA][28] , \chan_internal_f[DATA][27] , 
        \chan_internal_f[DATA][26] , \chan_internal_f[DATA][25] , 
        \chan_internal_f[DATA][24] , \chan_internal_f[DATA][23] , 
        \chan_internal_f[DATA][22] , \chan_internal_f[DATA][21] , 
        \chan_internal_f[DATA][20] , \chan_internal_f[DATA][19] , 
        \chan_internal_f[DATA][18] , \chan_internal_f[DATA][17] , 
        \chan_internal_f[DATA][16] , \chan_internal_f[DATA][15] , 
        \chan_internal_f[DATA][14] , \chan_internal_f[DATA][13] , 
        \chan_internal_f[DATA][12] , \chan_internal_f[DATA][11] , 
        \chan_internal_f[DATA][10] , \chan_internal_f[DATA][9] , 
        \chan_internal_f[DATA][8] , \chan_internal_f[DATA][7] , 
        \chan_internal_f[DATA][6] , \chan_internal_f[DATA][5] , 
        \chan_internal_f[DATA][4] , \chan_internal_f[DATA][3] , 
        \chan_internal_f[DATA][2] , \chan_internal_f[DATA][1] , 
        \chan_internal_f[DATA][0] }), .sel({sel[4:3], SYNOPSYS_UNCONNECTED__0, 
        sel[1:0]}) );
  channel_latch_1_xxxxxxxxx_4 token_latch ( .preset(n7), .left_in({
        \chan_internal_f[REQ] , \chan_internal_f[DATA][34] , 
        \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] , 
        \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] , 
        \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] , 
        \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] , 
        \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] , 
        \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] , 
        \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] , 
        \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] , 
        \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] , 
        \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] , 
        \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] , 
        \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] , 
        \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] , 
        \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] , 
        \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] , 
        \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] , 
        \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] }), .left_out(
        \chan_in_b[ACK] ), .right_out({\chan_out_f[REQ] , 
        \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , \chan_out_f[DATA][32] , 
        \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , \chan_out_f[DATA][29] , 
        \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , \chan_out_f[DATA][26] , 
        \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , \chan_out_f[DATA][23] , 
        \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , \chan_out_f[DATA][20] , 
        \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , \chan_out_f[DATA][17] , 
        \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , \chan_out_f[DATA][14] , 
        \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , \chan_out_f[DATA][11] , 
        \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , \chan_out_f[DATA][8] , 
        \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , \chan_out_f[DATA][5] , 
        \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , \chan_out_f[DATA][2] , 
        \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), .right_in(
        \chan_out_b[ACK] ), .lt_enable(lt_en) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chan_internal_f[REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(\chan_in_f[REQ] ), .Z(req_n) );
  HS65_LS_BFX9 U1 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U2 ( .A(n3), .Z(n2) );
  HS65_LS_BFX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_BFX9 U4 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U6 ( .A(req_n), .Z(n6) );
  HS65_LS_BFX9 U7 ( .A(preset), .Z(n7) );
endmodule


module hpu_comb_0_1_1 ( data_valid, data_in, preset, data_out, sel );
  input [34:0] data_in;
  output [34:0] data_out;
  output [4:0] sel;
  input data_valid, preset;
  wire   data_in_34, data_in_33, data_in_32, \data_in[31] , \data_in[30] ,
         \data_in[29] , \data_in[28] , \data_in[27] , \data_in[26] ,
         \data_in[25] , \data_in[24] , \data_in[23] , \data_in[22] ,
         \data_in[21] , \data_in[20] , \data_in[19] , \data_in[18] ,
         \data_in[17] , \data_in[16] , N23, N24, N26, N27, N28, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n15, n16, n17, n18;
  assign data_out[34] = data_in_34;
  assign data_in_34 = data_in[34];
  assign data_out[33] = data_in_33;
  assign data_in_33 = data_in[33];
  assign data_out[32] = data_in_32;
  assign data_in_32 = data_in[32];
  assign data_out[31] = \data_in[31] ;
  assign \data_in[31]  = data_in[31];
  assign data_out[30] = \data_in[30] ;
  assign \data_in[30]  = data_in[30];
  assign data_out[29] = \data_in[29] ;
  assign \data_in[29]  = data_in[29];
  assign data_out[28] = \data_in[28] ;
  assign \data_in[28]  = data_in[28];
  assign data_out[27] = \data_in[27] ;
  assign \data_in[27]  = data_in[27];
  assign data_out[26] = \data_in[26] ;
  assign \data_in[26]  = data_in[26];
  assign data_out[25] = \data_in[25] ;
  assign \data_in[25]  = data_in[25];
  assign data_out[24] = \data_in[24] ;
  assign \data_in[24]  = data_in[24];
  assign data_out[23] = \data_in[23] ;
  assign \data_in[23]  = data_in[23];
  assign data_out[22] = \data_in[22] ;
  assign \data_in[22]  = data_in[22];
  assign data_out[21] = \data_in[21] ;
  assign \data_in[21]  = data_in[21];
  assign data_out[20] = \data_in[20] ;
  assign \data_in[20]  = data_in[20];
  assign data_out[19] = \data_in[19] ;
  assign \data_in[19]  = data_in[19];
  assign data_out[18] = \data_in[18] ;
  assign \data_in[18]  = data_in[18];
  assign data_out[17] = \data_in[17] ;
  assign \data_in[17]  = data_in[17];
  assign data_out[16] = \data_in[16] ;
  assign \data_in[16]  = data_in[16];
  assign sel[1] = 1'b0;

  HS65_LS_LDHQX9 \sel_reg[4]  ( .G(N23), .D(N28), .Q(sel[4]) );
  HS65_LS_LDHQX9 \sel_reg[3]  ( .G(N23), .D(N27), .Q(sel[3]) );
  HS65_LS_LDHQX9 \sel_reg[2]  ( .G(N23), .D(N26), .Q(sel[2]) );
  HS65_LS_LDHQX9 \sel_reg[0]  ( .G(N23), .D(N24), .Q(sel[0]) );
  HS65_LS_OAI22X6 U4 ( .A(n6), .B(n18), .C(n2), .D(n7), .Z(data_out[7]) );
  HS65_LS_OAI22X6 U5 ( .A(n18), .B(n9), .C(n2), .D(n10), .Z(data_out[1]) );
  HS65_LS_OAI22X6 U6 ( .A(n18), .B(n8), .C(n2), .D(n9), .Z(data_out[3]) );
  HS65_LS_OAI22X6 U7 ( .A(n18), .B(n7), .C(n2), .D(n8), .Z(data_out[5]) );
  HS65_LS_OAI22X6 U8 ( .A(n18), .B(n5), .C(n2), .D(n6), .Z(data_out[9]) );
  HS65_LS_OAI22X6 U9 ( .A(n18), .B(n4), .C(n2), .D(n5), .Z(data_out[11]) );
  HS65_LS_OAI22X6 U10 ( .A(n18), .B(n3), .C(n2), .D(n4), .Z(data_out[13]) );
  HS65_LS_NAND3AX6 U11 ( .A(preset), .B(n17), .C(n2), .Z(n16) );
  HS65_LS_NOR3X4 U12 ( .A(n17), .B(preset), .C(n18), .Z(N28) );
  HS65_LS_IVX9 U13 ( .A(n18), .Z(n2) );
  HS65_LS_NOR3X4 U14 ( .A(n16), .B(n10), .C(n15), .Z(N27) );
  HS65_LS_NOR2AX3 U15 ( .A(n15), .B(n16), .Z(N26) );
  HS65_LS_NOR2X6 U16 ( .A(n2), .B(n3), .Z(data_out[15]) );
  HS65_LS_NAND2X14 U17 ( .A(data_in_34), .B(data_in_33), .Z(n18) );
  HS65_LS_IVX9 U18 ( .A(data_in[1]), .Z(n10) );
  HS65_LS_NAND2X7 U19 ( .A(data_in[0]), .B(n10), .Z(n17) );
  HS65_LS_NOR2X6 U20 ( .A(n10), .B(data_in[0]), .Z(n15) );
  HS65_LS_NOR2X6 U21 ( .A(data_in[1]), .B(n16), .Z(N24) );
  HS65_LS_IVX9 U22 ( .A(data_in[9]), .Z(n6) );
  HS65_LS_IVX9 U23 ( .A(data_in[3]), .Z(n9) );
  HS65_LS_IVX9 U24 ( .A(data_in[5]), .Z(n8) );
  HS65_LS_IVX9 U25 ( .A(data_in[7]), .Z(n7) );
  HS65_LS_IVX9 U26 ( .A(data_in[11]), .Z(n5) );
  HS65_LS_IVX9 U27 ( .A(data_in[13]), .Z(n4) );
  HS65_LS_IVX9 U28 ( .A(data_in[15]), .Z(n3) );
  HS65_LS_AO22X9 U29 ( .A(n2), .B(data_in[2]), .C(n18), .D(data_in[0]), .Z(
        data_out[0]) );
  HS65_LS_AO22X9 U30 ( .A(n2), .B(data_in[4]), .C(n18), .D(data_in[2]), .Z(
        data_out[2]) );
  HS65_LS_AO22X9 U31 ( .A(n2), .B(data_in[6]), .C(n18), .D(data_in[4]), .Z(
        data_out[4]) );
  HS65_LS_AO22X9 U32 ( .A(n2), .B(data_in[8]), .C(n18), .D(data_in[6]), .Z(
        data_out[6]) );
  HS65_LS_AO22X9 U33 ( .A(n2), .B(data_in[10]), .C(n18), .D(data_in[8]), .Z(
        data_out[8]) );
  HS65_LS_AO22X9 U34 ( .A(n2), .B(data_in[12]), .C(n18), .D(data_in[10]), .Z(
        data_out[10]) );
  HS65_LS_AO22X9 U35 ( .A(n2), .B(data_in[14]), .C(n18), .D(data_in[12]), .Z(
        data_out[12]) );
  HS65_LS_AND2X4 U36 ( .A(data_in[14]), .B(n18), .Z(data_out[14]) );
  HS65_LS_CB4I6X9 U37 ( .A(n2), .B(n1), .C(data_valid), .D(preset), .Z(N23) );
  HS65_LS_IVX9 U38 ( .A(data_in_34), .Z(n1) );
endmodule


module latch_controller_1_3 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_3 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_3 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n7) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_IVX9 U3 ( .A(N0), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_0_1_1 ( preset, .chan_in_f({\chan_in_f[REQ] , \chan_in_f[DATA][34] , 
        \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , 
        \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , 
        \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , 
        \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , 
        \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , 
        \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , 
        \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , 
        \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , 
        \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , 
        \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , 
        \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , 
        \chan_in_f[DATA][0] }), .chan_in_b(\chan_in_b[ACK] ), .chan_out_f({
        \chan_out_f[REQ] , \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , 
        \chan_out_f[DATA][32] , \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , 
        \chan_out_f[DATA][29] , \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , 
        \chan_out_f[DATA][26] , \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , 
        \chan_out_f[DATA][23] , \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , 
        \chan_out_f[DATA][20] , \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , 
        \chan_out_f[DATA][17] , \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , 
        \chan_out_f[DATA][14] , \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , 
        \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , 
        \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , 
        \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , 
        \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), 
    .chan_out_b(\chan_out_b[ACK] ), sel );
  output [4:0] sel;
  input preset, \chan_in_f[REQ] , \chan_in_f[DATA][34] , \chan_in_f[DATA][33] ,
         \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , \chan_in_f[DATA][30] ,
         \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , \chan_in_f[DATA][27] ,
         \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , \chan_in_f[DATA][24] ,
         \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , \chan_in_f[DATA][21] ,
         \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , \chan_in_f[DATA][18] ,
         \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , \chan_in_f[DATA][15] ,
         \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , \chan_in_f[DATA][12] ,
         \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , \chan_in_f[DATA][9] ,
         \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , \chan_in_f[DATA][6] ,
         \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , \chan_in_f[DATA][3] ,
         \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , \chan_in_f[DATA][0] ,
         \chan_out_b[ACK] ;
  output \chan_in_b[ACK] , \chan_out_f[REQ] , \chan_out_f[DATA][34] ,
         \chan_out_f[DATA][33] , \chan_out_f[DATA][32] ,
         \chan_out_f[DATA][31] , \chan_out_f[DATA][30] ,
         \chan_out_f[DATA][29] , \chan_out_f[DATA][28] ,
         \chan_out_f[DATA][27] , \chan_out_f[DATA][26] ,
         \chan_out_f[DATA][25] , \chan_out_f[DATA][24] ,
         \chan_out_f[DATA][23] , \chan_out_f[DATA][22] ,
         \chan_out_f[DATA][21] , \chan_out_f[DATA][20] ,
         \chan_out_f[DATA][19] , \chan_out_f[DATA][18] ,
         \chan_out_f[DATA][17] , \chan_out_f[DATA][16] ,
         \chan_out_f[DATA][15] , \chan_out_f[DATA][14] ,
         \chan_out_f[DATA][13] , \chan_out_f[DATA][12] ,
         \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] ,
         \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] ,
         \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] ,
         \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] ;
  wire   \chan_internal_f[REQ] , \chan_internal_f[DATA][34] ,
         \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] ,
         \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] ,
         \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] ,
         \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] ,
         \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] ,
         \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] ,
         \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] ,
         \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] ,
         \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] ,
         \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] ,
         \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] ,
         \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] ,
         \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] ,
         \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] ,
         \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] ,
         \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] ,
         \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] , req_n, lt_en,
         n1, n2, n3, n4, n5, n6, n7;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign sel[1] = 1'b0;

  hpu_comb_0_1_1 hpu_combinatorial ( .data_valid(lt_en), .data_in({
        \chan_in_f[DATA][34] , \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , 
        \chan_in_f[DATA][31] , \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , 
        \chan_in_f[DATA][28] , \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , 
        \chan_in_f[DATA][25] , \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , 
        \chan_in_f[DATA][22] , \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , 
        \chan_in_f[DATA][19] , \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , 
        \chan_in_f[DATA][16] , \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , 
        \chan_in_f[DATA][13] , \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , 
        \chan_in_f[DATA][10] , \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , 
        \chan_in_f[DATA][7] , \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , 
        \chan_in_f[DATA][4] , \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , 
        \chan_in_f[DATA][1] , \chan_in_f[DATA][0] }), .preset(n7), .data_out({
        \chan_internal_f[DATA][34] , \chan_internal_f[DATA][33] , 
        \chan_internal_f[DATA][32] , \chan_internal_f[DATA][31] , 
        \chan_internal_f[DATA][30] , \chan_internal_f[DATA][29] , 
        \chan_internal_f[DATA][28] , \chan_internal_f[DATA][27] , 
        \chan_internal_f[DATA][26] , \chan_internal_f[DATA][25] , 
        \chan_internal_f[DATA][24] , \chan_internal_f[DATA][23] , 
        \chan_internal_f[DATA][22] , \chan_internal_f[DATA][21] , 
        \chan_internal_f[DATA][20] , \chan_internal_f[DATA][19] , 
        \chan_internal_f[DATA][18] , \chan_internal_f[DATA][17] , 
        \chan_internal_f[DATA][16] , \chan_internal_f[DATA][15] , 
        \chan_internal_f[DATA][14] , \chan_internal_f[DATA][13] , 
        \chan_internal_f[DATA][12] , \chan_internal_f[DATA][11] , 
        \chan_internal_f[DATA][10] , \chan_internal_f[DATA][9] , 
        \chan_internal_f[DATA][8] , \chan_internal_f[DATA][7] , 
        \chan_internal_f[DATA][6] , \chan_internal_f[DATA][5] , 
        \chan_internal_f[DATA][4] , \chan_internal_f[DATA][3] , 
        \chan_internal_f[DATA][2] , \chan_internal_f[DATA][1] , 
        \chan_internal_f[DATA][0] }), .sel({sel[4:2], SYNOPSYS_UNCONNECTED__0, 
        sel[0]}) );
  channel_latch_1_xxxxxxxxx_3 token_latch ( .preset(n7), .left_in({
        \chan_internal_f[REQ] , \chan_internal_f[DATA][34] , 
        \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] , 
        \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] , 
        \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] , 
        \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] , 
        \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] , 
        \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] , 
        \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] , 
        \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] , 
        \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] , 
        \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] , 
        \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] , 
        \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] , 
        \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] , 
        \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] , 
        \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] , 
        \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] , 
        \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] }), .left_out(
        \chan_in_b[ACK] ), .right_out({\chan_out_f[REQ] , 
        \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , \chan_out_f[DATA][32] , 
        \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , \chan_out_f[DATA][29] , 
        \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , \chan_out_f[DATA][26] , 
        \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , \chan_out_f[DATA][23] , 
        \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , \chan_out_f[DATA][20] , 
        \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , \chan_out_f[DATA][17] , 
        \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , \chan_out_f[DATA][14] , 
        \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , \chan_out_f[DATA][11] , 
        \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , \chan_out_f[DATA][8] , 
        \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , \chan_out_f[DATA][5] , 
        \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , \chan_out_f[DATA][2] , 
        \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), .right_in(
        \chan_out_b[ACK] ), .lt_enable(lt_en) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chan_internal_f[REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(\chan_in_f[REQ] ), .Z(req_n) );
  HS65_LS_BFX9 U1 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U2 ( .A(n3), .Z(n2) );
  HS65_LS_BFX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_BFX9 U4 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U6 ( .A(req_n), .Z(n6) );
  HS65_LS_BFX9 U7 ( .A(preset), .Z(n7) );
endmodule


module hpu_comb_0_3_1 ( data_valid, data_in, preset, data_out, sel );
  input [34:0] data_in;
  output [34:0] data_out;
  output [4:0] sel;
  input data_valid, preset;
  wire   data_in_34, data_in_33, data_in_32, \data_in[31] , \data_in[30] ,
         \data_in[29] , \data_in[28] , \data_in[27] , \data_in[26] ,
         \data_in[25] , \data_in[24] , \data_in[23] , \data_in[22] ,
         \data_in[21] , \data_in[20] , \data_in[19] , \data_in[18] ,
         \data_in[17] , \data_in[16] , N25, N26, N27, N28, N30, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n15, n16, n17, n18;
  assign data_out[34] = data_in_34;
  assign data_in_34 = data_in[34];
  assign data_out[33] = data_in_33;
  assign data_in_33 = data_in[33];
  assign data_out[32] = data_in_32;
  assign data_in_32 = data_in[32];
  assign data_out[31] = \data_in[31] ;
  assign \data_in[31]  = data_in[31];
  assign data_out[30] = \data_in[30] ;
  assign \data_in[30]  = data_in[30];
  assign data_out[29] = \data_in[29] ;
  assign \data_in[29]  = data_in[29];
  assign data_out[28] = \data_in[28] ;
  assign \data_in[28]  = data_in[28];
  assign data_out[27] = \data_in[27] ;
  assign \data_in[27]  = data_in[27];
  assign data_out[26] = \data_in[26] ;
  assign \data_in[26]  = data_in[26];
  assign data_out[25] = \data_in[25] ;
  assign \data_in[25]  = data_in[25];
  assign data_out[24] = \data_in[24] ;
  assign \data_in[24]  = data_in[24];
  assign data_out[23] = \data_in[23] ;
  assign \data_in[23]  = data_in[23];
  assign data_out[22] = \data_in[22] ;
  assign \data_in[22]  = data_in[22];
  assign data_out[21] = \data_in[21] ;
  assign \data_in[21]  = data_in[21];
  assign data_out[20] = \data_in[20] ;
  assign \data_in[20]  = data_in[20];
  assign data_out[19] = \data_in[19] ;
  assign \data_in[19]  = data_in[19];
  assign data_out[18] = \data_in[18] ;
  assign \data_in[18]  = data_in[18];
  assign data_out[17] = \data_in[17] ;
  assign \data_in[17]  = data_in[17];
  assign data_out[16] = \data_in[16] ;
  assign \data_in[16]  = data_in[16];
  assign sel[3] = 1'b0;

  HS65_LS_LDHQX9 \sel_reg[4]  ( .G(N25), .D(N30), .Q(sel[4]) );
  HS65_LS_LDHQX9 \sel_reg[2]  ( .G(N25), .D(N28), .Q(sel[2]) );
  HS65_LS_LDHQX9 \sel_reg[1]  ( .G(N25), .D(N27), .Q(sel[1]) );
  HS65_LS_LDHQX9 \sel_reg[0]  ( .G(N25), .D(N26), .Q(sel[0]) );
  HS65_LS_OAI22X6 U4 ( .A(n18), .B(n9), .C(n2), .D(n10), .Z(data_out[0]) );
  HS65_LS_OAI22X6 U5 ( .A(n18), .B(n8), .C(n2), .D(n9), .Z(data_out[2]) );
  HS65_LS_OAI22X6 U6 ( .A(n18), .B(n7), .C(n2), .D(n8), .Z(data_out[4]) );
  HS65_LS_OAI22X6 U7 ( .A(n18), .B(n6), .C(n2), .D(n7), .Z(data_out[6]) );
  HS65_LS_OAI22X6 U8 ( .A(n18), .B(n5), .C(n2), .D(n6), .Z(data_out[8]) );
  HS65_LS_OAI22X6 U9 ( .A(n18), .B(n4), .C(n2), .D(n5), .Z(data_out[10]) );
  HS65_LS_OAI22X6 U10 ( .A(n18), .B(n3), .C(n2), .D(n4), .Z(data_out[12]) );
  HS65_LS_NAND3AX6 U11 ( .A(preset), .B(n17), .C(n2), .Z(n16) );
  HS65_LS_NOR3X4 U12 ( .A(n17), .B(preset), .C(n18), .Z(N30) );
  HS65_LS_IVX9 U13 ( .A(n18), .Z(n2) );
  HS65_LS_NOR2X6 U14 ( .A(n10), .B(n16), .Z(N27) );
  HS65_LS_NOR2AX3 U15 ( .A(n15), .B(n16), .Z(N26) );
  HS65_LS_NOR2X6 U16 ( .A(n2), .B(n3), .Z(data_out[14]) );
  HS65_LS_NAND2X14 U17 ( .A(data_in_34), .B(data_in_33), .Z(n18) );
  HS65_LS_NOR3X4 U18 ( .A(n16), .B(data_in[0]), .C(n15), .Z(N28) );
  HS65_LS_NAND2X7 U19 ( .A(data_in[0]), .B(data_in[1]), .Z(n17) );
  HS65_LS_NOR2X6 U20 ( .A(data_in[1]), .B(data_in[0]), .Z(n15) );
  HS65_LS_IVX9 U21 ( .A(data_in[0]), .Z(n10) );
  HS65_LS_IVX9 U22 ( .A(data_in[2]), .Z(n9) );
  HS65_LS_IVX9 U23 ( .A(data_in[4]), .Z(n8) );
  HS65_LS_IVX9 U24 ( .A(data_in[6]), .Z(n7) );
  HS65_LS_IVX9 U25 ( .A(data_in[8]), .Z(n6) );
  HS65_LS_IVX9 U26 ( .A(data_in[10]), .Z(n5) );
  HS65_LS_IVX9 U27 ( .A(data_in[12]), .Z(n4) );
  HS65_LS_IVX9 U28 ( .A(data_in[14]), .Z(n3) );
  HS65_LS_AO22X9 U29 ( .A(n2), .B(data_in[3]), .C(n18), .D(data_in[1]), .Z(
        data_out[1]) );
  HS65_LS_AO22X9 U30 ( .A(n2), .B(data_in[5]), .C(n18), .D(data_in[3]), .Z(
        data_out[3]) );
  HS65_LS_AO22X9 U31 ( .A(n2), .B(data_in[7]), .C(n18), .D(data_in[5]), .Z(
        data_out[5]) );
  HS65_LS_AO22X9 U32 ( .A(data_in[9]), .B(n2), .C(n18), .D(data_in[7]), .Z(
        data_out[7]) );
  HS65_LS_AO22X9 U33 ( .A(n2), .B(data_in[11]), .C(n18), .D(data_in[9]), .Z(
        data_out[9]) );
  HS65_LS_AO22X9 U34 ( .A(n2), .B(data_in[13]), .C(n18), .D(data_in[11]), .Z(
        data_out[11]) );
  HS65_LS_AO22X9 U35 ( .A(n2), .B(data_in[15]), .C(n18), .D(data_in[13]), .Z(
        data_out[13]) );
  HS65_LS_AND2X4 U36 ( .A(data_in[15]), .B(n18), .Z(data_out[15]) );
  HS65_LS_CB4I6X9 U37 ( .A(n2), .B(n1), .C(data_valid), .D(preset), .Z(N25) );
  HS65_LS_IVX9 U38 ( .A(data_in_34), .Z(n1) );
endmodule


module latch_controller_1_2 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_2 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_2 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n7) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_IVX9 U3 ( .A(N0), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_0_3_1 ( preset, .chan_in_f({\chan_in_f[REQ] , \chan_in_f[DATA][34] , 
        \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , 
        \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , 
        \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , 
        \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , 
        \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , 
        \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , 
        \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , 
        \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , 
        \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , 
        \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , 
        \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , 
        \chan_in_f[DATA][0] }), .chan_in_b(\chan_in_b[ACK] ), .chan_out_f({
        \chan_out_f[REQ] , \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , 
        \chan_out_f[DATA][32] , \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , 
        \chan_out_f[DATA][29] , \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , 
        \chan_out_f[DATA][26] , \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , 
        \chan_out_f[DATA][23] , \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , 
        \chan_out_f[DATA][20] , \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , 
        \chan_out_f[DATA][17] , \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , 
        \chan_out_f[DATA][14] , \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , 
        \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , 
        \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , 
        \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , 
        \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), 
    .chan_out_b(\chan_out_b[ACK] ), sel );
  output [4:0] sel;
  input preset, \chan_in_f[REQ] , \chan_in_f[DATA][34] , \chan_in_f[DATA][33] ,
         \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , \chan_in_f[DATA][30] ,
         \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , \chan_in_f[DATA][27] ,
         \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , \chan_in_f[DATA][24] ,
         \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , \chan_in_f[DATA][21] ,
         \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , \chan_in_f[DATA][18] ,
         \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , \chan_in_f[DATA][15] ,
         \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , \chan_in_f[DATA][12] ,
         \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , \chan_in_f[DATA][9] ,
         \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , \chan_in_f[DATA][6] ,
         \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , \chan_in_f[DATA][3] ,
         \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , \chan_in_f[DATA][0] ,
         \chan_out_b[ACK] ;
  output \chan_in_b[ACK] , \chan_out_f[REQ] , \chan_out_f[DATA][34] ,
         \chan_out_f[DATA][33] , \chan_out_f[DATA][32] ,
         \chan_out_f[DATA][31] , \chan_out_f[DATA][30] ,
         \chan_out_f[DATA][29] , \chan_out_f[DATA][28] ,
         \chan_out_f[DATA][27] , \chan_out_f[DATA][26] ,
         \chan_out_f[DATA][25] , \chan_out_f[DATA][24] ,
         \chan_out_f[DATA][23] , \chan_out_f[DATA][22] ,
         \chan_out_f[DATA][21] , \chan_out_f[DATA][20] ,
         \chan_out_f[DATA][19] , \chan_out_f[DATA][18] ,
         \chan_out_f[DATA][17] , \chan_out_f[DATA][16] ,
         \chan_out_f[DATA][15] , \chan_out_f[DATA][14] ,
         \chan_out_f[DATA][13] , \chan_out_f[DATA][12] ,
         \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] ,
         \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] ,
         \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] ,
         \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] ;
  wire   \chan_internal_f[REQ] , \chan_internal_f[DATA][34] ,
         \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] ,
         \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] ,
         \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] ,
         \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] ,
         \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] ,
         \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] ,
         \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] ,
         \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] ,
         \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] ,
         \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] ,
         \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] ,
         \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] ,
         \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] ,
         \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] ,
         \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] ,
         \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] ,
         \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] , req_n, lt_en,
         n1, n2, n3, n4, n5, n6, n7;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign sel[3] = 1'b0;

  hpu_comb_0_3_1 hpu_combinatorial ( .data_valid(lt_en), .data_in({
        \chan_in_f[DATA][34] , \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , 
        \chan_in_f[DATA][31] , \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , 
        \chan_in_f[DATA][28] , \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , 
        \chan_in_f[DATA][25] , \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , 
        \chan_in_f[DATA][22] , \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , 
        \chan_in_f[DATA][19] , \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , 
        \chan_in_f[DATA][16] , \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , 
        \chan_in_f[DATA][13] , \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , 
        \chan_in_f[DATA][10] , \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , 
        \chan_in_f[DATA][7] , \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , 
        \chan_in_f[DATA][4] , \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , 
        \chan_in_f[DATA][1] , \chan_in_f[DATA][0] }), .preset(n7), .data_out({
        \chan_internal_f[DATA][34] , \chan_internal_f[DATA][33] , 
        \chan_internal_f[DATA][32] , \chan_internal_f[DATA][31] , 
        \chan_internal_f[DATA][30] , \chan_internal_f[DATA][29] , 
        \chan_internal_f[DATA][28] , \chan_internal_f[DATA][27] , 
        \chan_internal_f[DATA][26] , \chan_internal_f[DATA][25] , 
        \chan_internal_f[DATA][24] , \chan_internal_f[DATA][23] , 
        \chan_internal_f[DATA][22] , \chan_internal_f[DATA][21] , 
        \chan_internal_f[DATA][20] , \chan_internal_f[DATA][19] , 
        \chan_internal_f[DATA][18] , \chan_internal_f[DATA][17] , 
        \chan_internal_f[DATA][16] , \chan_internal_f[DATA][15] , 
        \chan_internal_f[DATA][14] , \chan_internal_f[DATA][13] , 
        \chan_internal_f[DATA][12] , \chan_internal_f[DATA][11] , 
        \chan_internal_f[DATA][10] , \chan_internal_f[DATA][9] , 
        \chan_internal_f[DATA][8] , \chan_internal_f[DATA][7] , 
        \chan_internal_f[DATA][6] , \chan_internal_f[DATA][5] , 
        \chan_internal_f[DATA][4] , \chan_internal_f[DATA][3] , 
        \chan_internal_f[DATA][2] , \chan_internal_f[DATA][1] , 
        \chan_internal_f[DATA][0] }), .sel({sel[4], SYNOPSYS_UNCONNECTED__0, 
        sel[2:0]}) );
  channel_latch_1_xxxxxxxxx_2 token_latch ( .preset(n7), .left_in({
        \chan_internal_f[REQ] , \chan_internal_f[DATA][34] , 
        \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] , 
        \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] , 
        \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] , 
        \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] , 
        \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] , 
        \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] , 
        \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] , 
        \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] , 
        \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] , 
        \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] , 
        \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] , 
        \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] , 
        \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] , 
        \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] , 
        \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] , 
        \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] , 
        \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] }), .left_out(
        \chan_in_b[ACK] ), .right_out({\chan_out_f[REQ] , 
        \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , \chan_out_f[DATA][32] , 
        \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , \chan_out_f[DATA][29] , 
        \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , \chan_out_f[DATA][26] , 
        \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , \chan_out_f[DATA][23] , 
        \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , \chan_out_f[DATA][20] , 
        \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , \chan_out_f[DATA][17] , 
        \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , \chan_out_f[DATA][14] , 
        \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , \chan_out_f[DATA][11] , 
        \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , \chan_out_f[DATA][8] , 
        \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , \chan_out_f[DATA][5] , 
        \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , \chan_out_f[DATA][2] , 
        \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), .right_in(
        \chan_out_b[ACK] ), .lt_enable(lt_en) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chan_internal_f[REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(\chan_in_f[REQ] ), .Z(req_n) );
  HS65_LS_BFX9 U1 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U2 ( .A(n3), .Z(n2) );
  HS65_LS_BFX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_BFX9 U4 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U6 ( .A(req_n), .Z(n6) );
  HS65_LS_BFX9 U7 ( .A(preset), .Z(n7) );
endmodule


module hpu_comb_1_x_1 ( data_valid, data_in, preset, data_out, sel );
  input [34:0] data_in;
  output [34:0] data_out;
  output [4:0] sel;
  input data_valid, preset;
  wire   data_in_34, data_in_33, data_in_32, \data_in[31] , \data_in[30] ,
         \data_in[29] , \data_in[28] , \data_in[27] , \data_in[26] ,
         \data_in[25] , \data_in[24] , \data_in[23] , \data_in[22] ,
         \data_in[21] , \data_in[20] , \data_in[19] , \data_in[18] ,
         \data_in[17] , \data_in[16] , N19, N20, N21, N22, N23, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n22,
         n23, n24;
  assign data_out[34] = data_in_34;
  assign data_in_34 = data_in[34];
  assign data_out[33] = data_in_33;
  assign data_in_33 = data_in[33];
  assign data_out[32] = data_in_32;
  assign data_in_32 = data_in[32];
  assign data_out[31] = \data_in[31] ;
  assign \data_in[31]  = data_in[31];
  assign data_out[30] = \data_in[30] ;
  assign \data_in[30]  = data_in[30];
  assign data_out[29] = \data_in[29] ;
  assign \data_in[29]  = data_in[29];
  assign data_out[28] = \data_in[28] ;
  assign \data_in[28]  = data_in[28];
  assign data_out[27] = \data_in[27] ;
  assign \data_in[27]  = data_in[27];
  assign data_out[26] = \data_in[26] ;
  assign \data_in[26]  = data_in[26];
  assign data_out[25] = \data_in[25] ;
  assign \data_in[25]  = data_in[25];
  assign data_out[24] = \data_in[24] ;
  assign \data_in[24]  = data_in[24];
  assign data_out[23] = \data_in[23] ;
  assign \data_in[23]  = data_in[23];
  assign data_out[22] = \data_in[22] ;
  assign \data_in[22]  = data_in[22];
  assign data_out[21] = \data_in[21] ;
  assign \data_in[21]  = data_in[21];
  assign data_out[20] = \data_in[20] ;
  assign \data_in[20]  = data_in[20];
  assign data_out[19] = \data_in[19] ;
  assign \data_in[19]  = data_in[19];
  assign data_out[18] = \data_in[18] ;
  assign \data_in[18]  = data_in[18];
  assign data_out[17] = \data_in[17] ;
  assign \data_in[17]  = data_in[17];
  assign data_out[16] = \data_in[16] ;
  assign \data_in[16]  = data_in[16];
  assign sel[4] = 1'b0;

  HS65_LS_LDHQX9 \sel_reg[3]  ( .G(N19), .D(N23), .Q(sel[3]) );
  HS65_LS_LDHQX9 \sel_reg[2]  ( .G(N19), .D(N22), .Q(sel[2]) );
  HS65_LS_LDHQX9 \sel_reg[1]  ( .G(N19), .D(N21), .Q(sel[1]) );
  HS65_LS_LDHQX9 \sel_reg[0]  ( .G(N19), .D(N20), .Q(sel[0]) );
  HS65_LS_NAND2X21 U4 ( .A(data_in_34), .B(data_in_33), .Z(n24) );
  HS65_LS_NAND3AX6 U5 ( .A(preset), .B(n22), .C(n2), .Z(n23) );
  HS65_LS_OAI22X6 U6 ( .A(n9), .B(n24), .C(n2), .D(n11), .Z(data_out[7]) );
  HS65_LS_OAI22X6 U7 ( .A(n24), .B(n16), .C(n2), .D(n18), .Z(data_out[0]) );
  HS65_LS_OAI22X6 U8 ( .A(n24), .B(n15), .C(n2), .D(n17), .Z(data_out[1]) );
  HS65_LS_OAI22X6 U9 ( .A(n24), .B(n14), .C(n2), .D(n16), .Z(data_out[2]) );
  HS65_LS_OAI22X6 U10 ( .A(n24), .B(n13), .C(n2), .D(n15), .Z(data_out[3]) );
  HS65_LS_OAI22X6 U11 ( .A(n24), .B(n12), .C(n2), .D(n14), .Z(data_out[4]) );
  HS65_LS_OAI22X6 U12 ( .A(n24), .B(n11), .C(n2), .D(n13), .Z(data_out[5]) );
  HS65_LS_OAI22X6 U13 ( .A(n24), .B(n10), .C(n2), .D(n12), .Z(data_out[6]) );
  HS65_LS_OAI22X6 U14 ( .A(n24), .B(n8), .C(n2), .D(n10), .Z(data_out[8]) );
  HS65_LS_OAI22X6 U15 ( .A(n24), .B(n7), .C(n2), .D(n9), .Z(data_out[9]) );
  HS65_LS_OAI22X6 U16 ( .A(n24), .B(n6), .C(n2), .D(n8), .Z(data_out[10]) );
  HS65_LS_OAI22X6 U17 ( .A(n24), .B(n5), .C(n2), .D(n7), .Z(data_out[11]) );
  HS65_LS_OAI22X6 U18 ( .A(n24), .B(n4), .C(n2), .D(n6), .Z(data_out[12]) );
  HS65_LS_OAI22X6 U19 ( .A(n24), .B(n3), .C(n2), .D(n5), .Z(data_out[13]) );
  HS65_LS_IVX9 U20 ( .A(n24), .Z(n2) );
  HS65_LS_NOR3X4 U21 ( .A(n22), .B(preset), .C(n24), .Z(N20) );
  HS65_LS_NOR3X4 U22 ( .A(n23), .B(n17), .C(n18), .Z(N23) );
  HS65_LS_NAND2X7 U23 ( .A(n17), .B(n18), .Z(n22) );
  HS65_LS_NOR2X6 U24 ( .A(n2), .B(n4), .Z(data_out[14]) );
  HS65_LS_NOR2X6 U25 ( .A(n2), .B(n3), .Z(data_out[15]) );
  HS65_LS_IVX9 U26 ( .A(data_in[1]), .Z(n17) );
  HS65_LS_IVX9 U27 ( .A(data_in[0]), .Z(n18) );
  HS65_LS_NOR2X6 U28 ( .A(data_in[1]), .B(n23), .Z(N21) );
  HS65_LS_NOR2X6 U29 ( .A(data_in[0]), .B(n23), .Z(N22) );
  HS65_LS_IVX9 U30 ( .A(data_in[9]), .Z(n9) );
  HS65_LS_IVX9 U31 ( .A(data_in[2]), .Z(n16) );
  HS65_LS_IVX9 U32 ( .A(data_in[4]), .Z(n14) );
  HS65_LS_IVX9 U33 ( .A(data_in[5]), .Z(n13) );
  HS65_LS_IVX9 U34 ( .A(data_in[6]), .Z(n12) );
  HS65_LS_IVX9 U35 ( .A(data_in[8]), .Z(n10) );
  HS65_LS_IVX9 U36 ( .A(data_in[10]), .Z(n8) );
  HS65_LS_IVX9 U37 ( .A(data_in[12]), .Z(n6) );
  HS65_LS_IVX9 U38 ( .A(data_in[13]), .Z(n5) );
  HS65_LS_IVX9 U39 ( .A(data_in[14]), .Z(n4) );
  HS65_LS_IVX9 U40 ( .A(data_in[15]), .Z(n3) );
  HS65_LS_IVX9 U41 ( .A(data_in[3]), .Z(n15) );
  HS65_LS_IVX9 U42 ( .A(data_in[7]), .Z(n11) );
  HS65_LS_IVX9 U43 ( .A(data_in[11]), .Z(n7) );
  HS65_LS_CB4I6X9 U44 ( .A(n2), .B(n1), .C(data_valid), .D(preset), .Z(N19) );
  HS65_LS_IVX9 U45 ( .A(data_in_34), .Z(n1) );
endmodule


module latch_controller_1_1 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LS_NOR2AX3 U4 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_1_xxxxxxxxx_1 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, lt_gated, N5, n4, n5, n6, n7;
  assign N0 = preset;

  latch_controller_1_1 controller ( .preset(N0), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(\left_in[DATA][33] ), .Q(
        \right_out[DATA][33] ) );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(\left_in[DATA][32] ), .Q(
        \right_out[DATA][32] ) );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(\left_in[DATA][31] ), .Q(
        \right_out[DATA][31] ) );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(\left_in[DATA][30] ), .Q(
        \right_out[DATA][30] ) );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(\left_in[DATA][29] ), .Q(
        \right_out[DATA][29] ) );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(\left_in[DATA][28] ), .Q(
        \right_out[DATA][28] ) );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(\left_in[DATA][27] ), .Q(
        \right_out[DATA][27] ) );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(\left_in[DATA][26] ), .Q(
        \right_out[DATA][26] ) );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(\left_in[DATA][25] ), .Q(
        \right_out[DATA][25] ) );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(\left_in[DATA][24] ), .Q(
        \right_out[DATA][24] ) );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(\left_in[DATA][23] ), .Q(
        \right_out[DATA][23] ) );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(\left_in[DATA][22] ), .Q(
        \right_out[DATA][22] ) );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(\left_in[DATA][21] ), .Q(
        \right_out[DATA][21] ) );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(\left_in[DATA][20] ), .Q(
        \right_out[DATA][20] ) );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(\left_in[DATA][19] ), .Q(
        \right_out[DATA][19] ) );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(\left_in[DATA][18] ), .Q(
        \right_out[DATA][18] ) );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(\left_in[DATA][17] ), .Q(
        \right_out[DATA][17] ) );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(\left_in[DATA][16] ), .Q(
        \right_out[DATA][16] ) );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(\left_in[DATA][15] ), .Q(
        \right_out[DATA][15] ) );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(\left_in[DATA][14] ), .Q(
        \right_out[DATA][14] ) );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(\left_in[DATA][13] ), .Q(
        \right_out[DATA][13] ) );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(\left_in[DATA][12] ), .Q(
        \right_out[DATA][12] ) );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(\left_in[DATA][11] ), .Q(
        \right_out[DATA][11] ) );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(\left_in[DATA][10] ), .Q(
        \right_out[DATA][10] ) );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(\left_in[DATA][9] ), .Q(
        \right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(\left_in[DATA][8] ), .Q(
        \right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(\left_in[DATA][7] ), .Q(
        \right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(\left_in[DATA][6] ), .Q(
        \right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(\left_in[DATA][5] ), .Q(
        \right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(\left_in[DATA][4] ), .Q(
        \right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(\left_in[DATA][3] ), .Q(
        \right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(\left_in[DATA][2] ), .Q(
        \right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(\left_in[DATA][1] ), .Q(
        \right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(\left_in[DATA][0] ), .Q(
        \right_out[DATA][0] ) );
  HS65_LS_AND2X4 U6 ( .A(1'b1), .B(N0), .Z(n7) );
  HS65_LS_AND2X4 U7 ( .A(lt_gated), .B(n4), .Z(n6) );
  HS65_LS_OR2X9 U8 ( .A(n7), .B(n6), .Z(N5) );
  HS65_LS_LDLRQX9 type_out_reg ( .D(\left_in[DATA][34] ), .GN(n5), .RN(n4), 
        .Q(\right_out[DATA][34] ) );
  HS65_LS_IVX9 U3 ( .A(N0), .Z(n4) );
  HS65_LS_IVX9 U4 ( .A(lt_enable), .Z(n5) );
  HS65_LS_NAND2X7 U5 ( .A(\right_out[DATA][34] ), .B(n5), .Z(lt_gated) );
endmodule


module hpu_1_x_1 ( preset, .chan_in_f({\chan_in_f[REQ] , \chan_in_f[DATA][34] , 
        \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , 
        \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , 
        \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , 
        \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , 
        \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , 
        \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , 
        \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , 
        \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , 
        \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , 
        \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , 
        \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , 
        \chan_in_f[DATA][0] }), .chan_in_b(\chan_in_b[ACK] ), .chan_out_f({
        \chan_out_f[REQ] , \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , 
        \chan_out_f[DATA][32] , \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , 
        \chan_out_f[DATA][29] , \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , 
        \chan_out_f[DATA][26] , \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , 
        \chan_out_f[DATA][23] , \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , 
        \chan_out_f[DATA][20] , \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , 
        \chan_out_f[DATA][17] , \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , 
        \chan_out_f[DATA][14] , \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , 
        \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , 
        \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , 
        \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , 
        \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), 
    .chan_out_b(\chan_out_b[ACK] ), sel );
  output [4:0] sel;
  input preset, \chan_in_f[REQ] , \chan_in_f[DATA][34] , \chan_in_f[DATA][33] ,
         \chan_in_f[DATA][32] , \chan_in_f[DATA][31] , \chan_in_f[DATA][30] ,
         \chan_in_f[DATA][29] , \chan_in_f[DATA][28] , \chan_in_f[DATA][27] ,
         \chan_in_f[DATA][26] , \chan_in_f[DATA][25] , \chan_in_f[DATA][24] ,
         \chan_in_f[DATA][23] , \chan_in_f[DATA][22] , \chan_in_f[DATA][21] ,
         \chan_in_f[DATA][20] , \chan_in_f[DATA][19] , \chan_in_f[DATA][18] ,
         \chan_in_f[DATA][17] , \chan_in_f[DATA][16] , \chan_in_f[DATA][15] ,
         \chan_in_f[DATA][14] , \chan_in_f[DATA][13] , \chan_in_f[DATA][12] ,
         \chan_in_f[DATA][11] , \chan_in_f[DATA][10] , \chan_in_f[DATA][9] ,
         \chan_in_f[DATA][8] , \chan_in_f[DATA][7] , \chan_in_f[DATA][6] ,
         \chan_in_f[DATA][5] , \chan_in_f[DATA][4] , \chan_in_f[DATA][3] ,
         \chan_in_f[DATA][2] , \chan_in_f[DATA][1] , \chan_in_f[DATA][0] ,
         \chan_out_b[ACK] ;
  output \chan_in_b[ACK] , \chan_out_f[REQ] , \chan_out_f[DATA][34] ,
         \chan_out_f[DATA][33] , \chan_out_f[DATA][32] ,
         \chan_out_f[DATA][31] , \chan_out_f[DATA][30] ,
         \chan_out_f[DATA][29] , \chan_out_f[DATA][28] ,
         \chan_out_f[DATA][27] , \chan_out_f[DATA][26] ,
         \chan_out_f[DATA][25] , \chan_out_f[DATA][24] ,
         \chan_out_f[DATA][23] , \chan_out_f[DATA][22] ,
         \chan_out_f[DATA][21] , \chan_out_f[DATA][20] ,
         \chan_out_f[DATA][19] , \chan_out_f[DATA][18] ,
         \chan_out_f[DATA][17] , \chan_out_f[DATA][16] ,
         \chan_out_f[DATA][15] , \chan_out_f[DATA][14] ,
         \chan_out_f[DATA][13] , \chan_out_f[DATA][12] ,
         \chan_out_f[DATA][11] , \chan_out_f[DATA][10] , \chan_out_f[DATA][9] ,
         \chan_out_f[DATA][8] , \chan_out_f[DATA][7] , \chan_out_f[DATA][6] ,
         \chan_out_f[DATA][5] , \chan_out_f[DATA][4] , \chan_out_f[DATA][3] ,
         \chan_out_f[DATA][2] , \chan_out_f[DATA][1] , \chan_out_f[DATA][0] ;
  wire   \chan_internal_f[REQ] , \chan_internal_f[DATA][34] ,
         \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] ,
         \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] ,
         \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] ,
         \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] ,
         \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] ,
         \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] ,
         \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] ,
         \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] ,
         \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] ,
         \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] ,
         \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] ,
         \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] ,
         \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] ,
         \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] ,
         \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] ,
         \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] ,
         \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] , req_n, lt_en,
         n1, n2, n3, n4, n5, n6, n7;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign sel[4] = 1'b0;

  hpu_comb_1_x_1 hpu_combinatorial ( .data_valid(lt_en), .data_in({
        \chan_in_f[DATA][34] , \chan_in_f[DATA][33] , \chan_in_f[DATA][32] , 
        \chan_in_f[DATA][31] , \chan_in_f[DATA][30] , \chan_in_f[DATA][29] , 
        \chan_in_f[DATA][28] , \chan_in_f[DATA][27] , \chan_in_f[DATA][26] , 
        \chan_in_f[DATA][25] , \chan_in_f[DATA][24] , \chan_in_f[DATA][23] , 
        \chan_in_f[DATA][22] , \chan_in_f[DATA][21] , \chan_in_f[DATA][20] , 
        \chan_in_f[DATA][19] , \chan_in_f[DATA][18] , \chan_in_f[DATA][17] , 
        \chan_in_f[DATA][16] , \chan_in_f[DATA][15] , \chan_in_f[DATA][14] , 
        \chan_in_f[DATA][13] , \chan_in_f[DATA][12] , \chan_in_f[DATA][11] , 
        \chan_in_f[DATA][10] , \chan_in_f[DATA][9] , \chan_in_f[DATA][8] , 
        \chan_in_f[DATA][7] , \chan_in_f[DATA][6] , \chan_in_f[DATA][5] , 
        \chan_in_f[DATA][4] , \chan_in_f[DATA][3] , \chan_in_f[DATA][2] , 
        \chan_in_f[DATA][1] , \chan_in_f[DATA][0] }), .preset(n7), .data_out({
        \chan_internal_f[DATA][34] , \chan_internal_f[DATA][33] , 
        \chan_internal_f[DATA][32] , \chan_internal_f[DATA][31] , 
        \chan_internal_f[DATA][30] , \chan_internal_f[DATA][29] , 
        \chan_internal_f[DATA][28] , \chan_internal_f[DATA][27] , 
        \chan_internal_f[DATA][26] , \chan_internal_f[DATA][25] , 
        \chan_internal_f[DATA][24] , \chan_internal_f[DATA][23] , 
        \chan_internal_f[DATA][22] , \chan_internal_f[DATA][21] , 
        \chan_internal_f[DATA][20] , \chan_internal_f[DATA][19] , 
        \chan_internal_f[DATA][18] , \chan_internal_f[DATA][17] , 
        \chan_internal_f[DATA][16] , \chan_internal_f[DATA][15] , 
        \chan_internal_f[DATA][14] , \chan_internal_f[DATA][13] , 
        \chan_internal_f[DATA][12] , \chan_internal_f[DATA][11] , 
        \chan_internal_f[DATA][10] , \chan_internal_f[DATA][9] , 
        \chan_internal_f[DATA][8] , \chan_internal_f[DATA][7] , 
        \chan_internal_f[DATA][6] , \chan_internal_f[DATA][5] , 
        \chan_internal_f[DATA][4] , \chan_internal_f[DATA][3] , 
        \chan_internal_f[DATA][2] , \chan_internal_f[DATA][1] , 
        \chan_internal_f[DATA][0] }), .sel({SYNOPSYS_UNCONNECTED__0, sel[3:0]}) );
  channel_latch_1_xxxxxxxxx_1 token_latch ( .preset(n7), .left_in({
        \chan_internal_f[REQ] , \chan_internal_f[DATA][34] , 
        \chan_internal_f[DATA][33] , \chan_internal_f[DATA][32] , 
        \chan_internal_f[DATA][31] , \chan_internal_f[DATA][30] , 
        \chan_internal_f[DATA][29] , \chan_internal_f[DATA][28] , 
        \chan_internal_f[DATA][27] , \chan_internal_f[DATA][26] , 
        \chan_internal_f[DATA][25] , \chan_internal_f[DATA][24] , 
        \chan_internal_f[DATA][23] , \chan_internal_f[DATA][22] , 
        \chan_internal_f[DATA][21] , \chan_internal_f[DATA][20] , 
        \chan_internal_f[DATA][19] , \chan_internal_f[DATA][18] , 
        \chan_internal_f[DATA][17] , \chan_internal_f[DATA][16] , 
        \chan_internal_f[DATA][15] , \chan_internal_f[DATA][14] , 
        \chan_internal_f[DATA][13] , \chan_internal_f[DATA][12] , 
        \chan_internal_f[DATA][11] , \chan_internal_f[DATA][10] , 
        \chan_internal_f[DATA][9] , \chan_internal_f[DATA][8] , 
        \chan_internal_f[DATA][7] , \chan_internal_f[DATA][6] , 
        \chan_internal_f[DATA][5] , \chan_internal_f[DATA][4] , 
        \chan_internal_f[DATA][3] , \chan_internal_f[DATA][2] , 
        \chan_internal_f[DATA][1] , \chan_internal_f[DATA][0] }), .left_out(
        \chan_in_b[ACK] ), .right_out({\chan_out_f[REQ] , 
        \chan_out_f[DATA][34] , \chan_out_f[DATA][33] , \chan_out_f[DATA][32] , 
        \chan_out_f[DATA][31] , \chan_out_f[DATA][30] , \chan_out_f[DATA][29] , 
        \chan_out_f[DATA][28] , \chan_out_f[DATA][27] , \chan_out_f[DATA][26] , 
        \chan_out_f[DATA][25] , \chan_out_f[DATA][24] , \chan_out_f[DATA][23] , 
        \chan_out_f[DATA][22] , \chan_out_f[DATA][21] , \chan_out_f[DATA][20] , 
        \chan_out_f[DATA][19] , \chan_out_f[DATA][18] , \chan_out_f[DATA][17] , 
        \chan_out_f[DATA][16] , \chan_out_f[DATA][15] , \chan_out_f[DATA][14] , 
        \chan_out_f[DATA][13] , \chan_out_f[DATA][12] , \chan_out_f[DATA][11] , 
        \chan_out_f[DATA][10] , \chan_out_f[DATA][9] , \chan_out_f[DATA][8] , 
        \chan_out_f[DATA][7] , \chan_out_f[DATA][6] , \chan_out_f[DATA][5] , 
        \chan_out_f[DATA][4] , \chan_out_f[DATA][3] , \chan_out_f[DATA][2] , 
        \chan_out_f[DATA][1] , \chan_out_f[DATA][0] }), .right_in(
        \chan_out_b[ACK] ), .lt_enable(lt_en) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chan_internal_f[REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(\chan_in_f[REQ] ), .Z(req_n) );
  HS65_LS_BFX9 U1 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U2 ( .A(n3), .Z(n2) );
  HS65_LS_BFX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_BFX9 U4 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U6 ( .A(req_n), .Z(n6) );
  HS65_LS_BFX9 U7 ( .A(preset), .Z(n7) );
endmodule


module sr_latch_1_2 ( s, r, q, qn );
  input s, r;
  output q, qn;
  wire   N3, n1;

  HS65_LS_AND2X4 C9 ( .A(n1), .B(N3), .Z(qn) );
  HS65_LH_NOR2X3 U1 ( .A(r), .B(qn), .Z(q) );
  HS65_LS_IVX9 U2 ( .A(q), .Z(N3) );
  HS65_LS_IVX9 U3 ( .A(s), .Z(n1) );
endmodule


module c_gate_generic_1_5_2 ( preset, \input , \output  );
  input [4:0] \input ;
  input preset;
  output \output ;
  wire   set, reset, n1, n4, n5;

  sr_latch_1_2 latch ( .s(set), .r(reset), .q(\output ) );
  HS65_LS_NOR3X4 U3 ( .A(\input [3]), .B(preset), .C(\input [4]), .Z(n4) );
  HS65_LS_NOR4ABX2 U4 ( .A(n1), .B(n4), .C(\input [2]), .D(\input [1]), .Z(
        reset) );
  HS65_LS_AO31X9 U5 ( .A(n5), .B(\input [3]), .C(\input [4]), .D(preset), .Z(
        set) );
  HS65_LS_IVX9 U6 ( .A(\input [0]), .Z(n1) );
  HS65_LS_AND3X9 U7 ( .A(\input [1]), .B(\input [0]), .C(\input [2]), .Z(n5)
         );
endmodule


module sr_latch_1_1 ( s, r, q, qn );
  input s, r;
  output q, qn;
  wire   N3, n1;

  HS65_LS_AND2X4 C9 ( .A(n1), .B(N3), .Z(qn) );
  HS65_LS_IVX9 U1 ( .A(q), .Z(N3) );
  HS65_LS_IVX9 U2 ( .A(s), .Z(n1) );
  HS65_LS_NOR2X6 U3 ( .A(r), .B(qn), .Z(q) );
endmodule


module c_gate_generic_1_5_1 ( preset, \input , \output  );
  input [4:0] \input ;
  input preset;
  output \output ;
  wire   set, reset, n1, n4, n5;

  sr_latch_1_1 latch ( .s(set), .r(reset), .q(\output ) );
  HS65_LS_NOR3X4 U3 ( .A(\input [3]), .B(preset), .C(\input [4]), .Z(n4) );
  HS65_LS_NOR4ABX2 U4 ( .A(n1), .B(n4), .C(\input [2]), .D(\input [1]), .Z(
        reset) );
  HS65_LS_AO31X9 U5 ( .A(n5), .B(\input [3]), .C(\input [4]), .D(preset), .Z(
        set) );
  HS65_LS_IVX9 U6 ( .A(\input [0]), .Z(n1) );
  HS65_LS_AND3X9 U7 ( .A(\input [1]), .B(\input [0]), .C(\input [2]), .Z(n5)
         );
endmodule


module crossbar_1 ( preset, .switch_sel({\switch_sel[4][4] , 
        \switch_sel[4][3] , \switch_sel[4][2] , \switch_sel[4][1] , 
        \switch_sel[4][0] , \switch_sel[3][4] , \switch_sel[3][3] , 
        \switch_sel[3][2] , \switch_sel[3][1] , \switch_sel[3][0] , 
        \switch_sel[2][4] , \switch_sel[2][3] , \switch_sel[2][2] , 
        \switch_sel[2][1] , \switch_sel[2][0] , \switch_sel[1][4] , 
        \switch_sel[1][3] , \switch_sel[1][2] , \switch_sel[1][1] , 
        \switch_sel[1][0] , \switch_sel[0][4] , \switch_sel[0][3] , 
        \switch_sel[0][2] , \switch_sel[0][1] , \switch_sel[0][0] }), 
    .chs_in_f({\chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] , 
        \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] , 
        \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] , 
        \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] , 
        \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] , 
        \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] , 
        \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] , 
        \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] , 
        \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] , 
        \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] , 
        \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] , 
        \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] , 
        \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] , 
        \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] , \chs_in_f[4][DATA][7] , 
        \chs_in_f[4][DATA][6] , \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] , 
        \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] , \chs_in_f[4][DATA][1] , 
        \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] , \chs_in_f[3][DATA][34] , 
        \chs_in_f[3][DATA][33] , \chs_in_f[3][DATA][32] , 
        \chs_in_f[3][DATA][31] , \chs_in_f[3][DATA][30] , 
        \chs_in_f[3][DATA][29] , \chs_in_f[3][DATA][28] , 
        \chs_in_f[3][DATA][27] , \chs_in_f[3][DATA][26] , 
        \chs_in_f[3][DATA][25] , \chs_in_f[3][DATA][24] , 
        \chs_in_f[3][DATA][23] , \chs_in_f[3][DATA][22] , 
        \chs_in_f[3][DATA][21] , \chs_in_f[3][DATA][20] , 
        \chs_in_f[3][DATA][19] , \chs_in_f[3][DATA][18] , 
        \chs_in_f[3][DATA][17] , \chs_in_f[3][DATA][16] , 
        \chs_in_f[3][DATA][15] , \chs_in_f[3][DATA][14] , 
        \chs_in_f[3][DATA][13] , \chs_in_f[3][DATA][12] , 
        \chs_in_f[3][DATA][11] , \chs_in_f[3][DATA][10] , 
        \chs_in_f[3][DATA][9] , \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] , 
        \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] , \chs_in_f[3][DATA][4] , 
        \chs_in_f[3][DATA][3] , \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] , 
        \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] , 
        \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] , 
        \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] , 
        \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] , 
        \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] , 
        \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] , 
        \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] , 
        \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] , 
        \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] , 
        \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] , 
        \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] , 
        \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] , 
        \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] , 
        \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] , \chs_in_f[2][DATA][7] , 
        \chs_in_f[2][DATA][6] , \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] , 
        \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] , \chs_in_f[2][DATA][1] , 
        \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] , \chs_in_f[1][DATA][34] , 
        \chs_in_f[1][DATA][33] , \chs_in_f[1][DATA][32] , 
        \chs_in_f[1][DATA][31] , \chs_in_f[1][DATA][30] , 
        \chs_in_f[1][DATA][29] , \chs_in_f[1][DATA][28] , 
        \chs_in_f[1][DATA][27] , \chs_in_f[1][DATA][26] , 
        \chs_in_f[1][DATA][25] , \chs_in_f[1][DATA][24] , 
        \chs_in_f[1][DATA][23] , \chs_in_f[1][DATA][22] , 
        \chs_in_f[1][DATA][21] , \chs_in_f[1][DATA][20] , 
        \chs_in_f[1][DATA][19] , \chs_in_f[1][DATA][18] , 
        \chs_in_f[1][DATA][17] , \chs_in_f[1][DATA][16] , 
        \chs_in_f[1][DATA][15] , \chs_in_f[1][DATA][14] , 
        \chs_in_f[1][DATA][13] , \chs_in_f[1][DATA][12] , 
        \chs_in_f[1][DATA][11] , \chs_in_f[1][DATA][10] , 
        \chs_in_f[1][DATA][9] , \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] , 
        \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] , \chs_in_f[1][DATA][4] , 
        \chs_in_f[1][DATA][3] , \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] , 
        \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] , 
        \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] , 
        \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] , 
        \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] , 
        \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] , 
        \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] , 
        \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] , 
        \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] , 
        \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] , 
        \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] , 
        \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] , 
        \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] , 
        \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] , 
        \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] , \chs_in_f[0][DATA][7] , 
        \chs_in_f[0][DATA][6] , \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] , 
        \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] , \chs_in_f[0][DATA][1] , 
        \chs_in_f[0][DATA][0] }), .chs_in_b({\chs_in_b[4][ACK] , 
        \chs_in_b[3][ACK] , \chs_in_b[2][ACK] , \chs_in_b[1][ACK] , 
        \chs_in_b[0][ACK] }), .chs_out_f({\chs_out_f[4][REQ] , 
        \chs_out_f[4][DATA][34] , \chs_out_f[4][DATA][33] , 
        \chs_out_f[4][DATA][32] , \chs_out_f[4][DATA][31] , 
        \chs_out_f[4][DATA][30] , \chs_out_f[4][DATA][29] , 
        \chs_out_f[4][DATA][28] , \chs_out_f[4][DATA][27] , 
        \chs_out_f[4][DATA][26] , \chs_out_f[4][DATA][25] , 
        \chs_out_f[4][DATA][24] , \chs_out_f[4][DATA][23] , 
        \chs_out_f[4][DATA][22] , \chs_out_f[4][DATA][21] , 
        \chs_out_f[4][DATA][20] , \chs_out_f[4][DATA][19] , 
        \chs_out_f[4][DATA][18] , \chs_out_f[4][DATA][17] , 
        \chs_out_f[4][DATA][16] , \chs_out_f[4][DATA][15] , 
        \chs_out_f[4][DATA][14] , \chs_out_f[4][DATA][13] , 
        \chs_out_f[4][DATA][12] , \chs_out_f[4][DATA][11] , 
        \chs_out_f[4][DATA][10] , \chs_out_f[4][DATA][9] , 
        \chs_out_f[4][DATA][8] , \chs_out_f[4][DATA][7] , 
        \chs_out_f[4][DATA][6] , \chs_out_f[4][DATA][5] , 
        \chs_out_f[4][DATA][4] , \chs_out_f[4][DATA][3] , 
        \chs_out_f[4][DATA][2] , \chs_out_f[4][DATA][1] , 
        \chs_out_f[4][DATA][0] , \chs_out_f[3][REQ] , \chs_out_f[3][DATA][34] , 
        \chs_out_f[3][DATA][33] , \chs_out_f[3][DATA][32] , 
        \chs_out_f[3][DATA][31] , \chs_out_f[3][DATA][30] , 
        \chs_out_f[3][DATA][29] , \chs_out_f[3][DATA][28] , 
        \chs_out_f[3][DATA][27] , \chs_out_f[3][DATA][26] , 
        \chs_out_f[3][DATA][25] , \chs_out_f[3][DATA][24] , 
        \chs_out_f[3][DATA][23] , \chs_out_f[3][DATA][22] , 
        \chs_out_f[3][DATA][21] , \chs_out_f[3][DATA][20] , 
        \chs_out_f[3][DATA][19] , \chs_out_f[3][DATA][18] , 
        \chs_out_f[3][DATA][17] , \chs_out_f[3][DATA][16] , 
        \chs_out_f[3][DATA][15] , \chs_out_f[3][DATA][14] , 
        \chs_out_f[3][DATA][13] , \chs_out_f[3][DATA][12] , 
        \chs_out_f[3][DATA][11] , \chs_out_f[3][DATA][10] , 
        \chs_out_f[3][DATA][9] , \chs_out_f[3][DATA][8] , 
        \chs_out_f[3][DATA][7] , \chs_out_f[3][DATA][6] , 
        \chs_out_f[3][DATA][5] , \chs_out_f[3][DATA][4] , 
        \chs_out_f[3][DATA][3] , \chs_out_f[3][DATA][2] , 
        \chs_out_f[3][DATA][1] , \chs_out_f[3][DATA][0] , \chs_out_f[2][REQ] , 
        \chs_out_f[2][DATA][34] , \chs_out_f[2][DATA][33] , 
        \chs_out_f[2][DATA][32] , \chs_out_f[2][DATA][31] , 
        \chs_out_f[2][DATA][30] , \chs_out_f[2][DATA][29] , 
        \chs_out_f[2][DATA][28] , \chs_out_f[2][DATA][27] , 
        \chs_out_f[2][DATA][26] , \chs_out_f[2][DATA][25] , 
        \chs_out_f[2][DATA][24] , \chs_out_f[2][DATA][23] , 
        \chs_out_f[2][DATA][22] , \chs_out_f[2][DATA][21] , 
        \chs_out_f[2][DATA][20] , \chs_out_f[2][DATA][19] , 
        \chs_out_f[2][DATA][18] , \chs_out_f[2][DATA][17] , 
        \chs_out_f[2][DATA][16] , \chs_out_f[2][DATA][15] , 
        \chs_out_f[2][DATA][14] , \chs_out_f[2][DATA][13] , 
        \chs_out_f[2][DATA][12] , \chs_out_f[2][DATA][11] , 
        \chs_out_f[2][DATA][10] , \chs_out_f[2][DATA][9] , 
        \chs_out_f[2][DATA][8] , \chs_out_f[2][DATA][7] , 
        \chs_out_f[2][DATA][6] , \chs_out_f[2][DATA][5] , 
        \chs_out_f[2][DATA][4] , \chs_out_f[2][DATA][3] , 
        \chs_out_f[2][DATA][2] , \chs_out_f[2][DATA][1] , 
        \chs_out_f[2][DATA][0] , \chs_out_f[1][REQ] , \chs_out_f[1][DATA][34] , 
        \chs_out_f[1][DATA][33] , \chs_out_f[1][DATA][32] , 
        \chs_out_f[1][DATA][31] , \chs_out_f[1][DATA][30] , 
        \chs_out_f[1][DATA][29] , \chs_out_f[1][DATA][28] , 
        \chs_out_f[1][DATA][27] , \chs_out_f[1][DATA][26] , 
        \chs_out_f[1][DATA][25] , \chs_out_f[1][DATA][24] , 
        \chs_out_f[1][DATA][23] , \chs_out_f[1][DATA][22] , 
        \chs_out_f[1][DATA][21] , \chs_out_f[1][DATA][20] , 
        \chs_out_f[1][DATA][19] , \chs_out_f[1][DATA][18] , 
        \chs_out_f[1][DATA][17] , \chs_out_f[1][DATA][16] , 
        \chs_out_f[1][DATA][15] , \chs_out_f[1][DATA][14] , 
        \chs_out_f[1][DATA][13] , \chs_out_f[1][DATA][12] , 
        \chs_out_f[1][DATA][11] , \chs_out_f[1][DATA][10] , 
        \chs_out_f[1][DATA][9] , \chs_out_f[1][DATA][8] , 
        \chs_out_f[1][DATA][7] , \chs_out_f[1][DATA][6] , 
        \chs_out_f[1][DATA][5] , \chs_out_f[1][DATA][4] , 
        \chs_out_f[1][DATA][3] , \chs_out_f[1][DATA][2] , 
        \chs_out_f[1][DATA][1] , \chs_out_f[1][DATA][0] , \chs_out_f[0][REQ] , 
        \chs_out_f[0][DATA][34] , \chs_out_f[0][DATA][33] , 
        \chs_out_f[0][DATA][32] , \chs_out_f[0][DATA][31] , 
        \chs_out_f[0][DATA][30] , \chs_out_f[0][DATA][29] , 
        \chs_out_f[0][DATA][28] , \chs_out_f[0][DATA][27] , 
        \chs_out_f[0][DATA][26] , \chs_out_f[0][DATA][25] , 
        \chs_out_f[0][DATA][24] , \chs_out_f[0][DATA][23] , 
        \chs_out_f[0][DATA][22] , \chs_out_f[0][DATA][21] , 
        \chs_out_f[0][DATA][20] , \chs_out_f[0][DATA][19] , 
        \chs_out_f[0][DATA][18] , \chs_out_f[0][DATA][17] , 
        \chs_out_f[0][DATA][16] , \chs_out_f[0][DATA][15] , 
        \chs_out_f[0][DATA][14] , \chs_out_f[0][DATA][13] , 
        \chs_out_f[0][DATA][12] , \chs_out_f[0][DATA][11] , 
        \chs_out_f[0][DATA][10] , \chs_out_f[0][DATA][9] , 
        \chs_out_f[0][DATA][8] , \chs_out_f[0][DATA][7] , 
        \chs_out_f[0][DATA][6] , \chs_out_f[0][DATA][5] , 
        \chs_out_f[0][DATA][4] , \chs_out_f[0][DATA][3] , 
        \chs_out_f[0][DATA][2] , \chs_out_f[0][DATA][1] , 
        \chs_out_f[0][DATA][0] }), .chs_out_b({\chs_out_b[4][ACK] , 
        \chs_out_b[3][ACK] , \chs_out_b[2][ACK] , \chs_out_b[1][ACK] , 
        \chs_out_b[0][ACK] }) );
  input preset, \switch_sel[4][4] , \switch_sel[4][3] , \switch_sel[4][2] ,
         \switch_sel[4][1] , \switch_sel[4][0] , \switch_sel[3][4] ,
         \switch_sel[3][3] , \switch_sel[3][2] , \switch_sel[3][1] ,
         \switch_sel[3][0] , \switch_sel[2][4] , \switch_sel[2][3] ,
         \switch_sel[2][2] , \switch_sel[2][1] , \switch_sel[2][0] ,
         \switch_sel[1][4] , \switch_sel[1][3] , \switch_sel[1][2] ,
         \switch_sel[1][1] , \switch_sel[1][0] , \switch_sel[0][4] ,
         \switch_sel[0][3] , \switch_sel[0][2] , \switch_sel[0][1] ,
         \switch_sel[0][0] , \chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] ,
         \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] ,
         \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] ,
         \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] ,
         \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] ,
         \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] ,
         \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] ,
         \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] ,
         \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] ,
         \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] ,
         \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] ,
         \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] ,
         \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] ,
         \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] ,
         \chs_in_f[4][DATA][7] , \chs_in_f[4][DATA][6] ,
         \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] ,
         \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] ,
         \chs_in_f[4][DATA][1] , \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] ,
         \chs_in_f[3][DATA][34] , \chs_in_f[3][DATA][33] ,
         \chs_in_f[3][DATA][32] , \chs_in_f[3][DATA][31] ,
         \chs_in_f[3][DATA][30] , \chs_in_f[3][DATA][29] ,
         \chs_in_f[3][DATA][28] , \chs_in_f[3][DATA][27] ,
         \chs_in_f[3][DATA][26] , \chs_in_f[3][DATA][25] ,
         \chs_in_f[3][DATA][24] , \chs_in_f[3][DATA][23] ,
         \chs_in_f[3][DATA][22] , \chs_in_f[3][DATA][21] ,
         \chs_in_f[3][DATA][20] , \chs_in_f[3][DATA][19] ,
         \chs_in_f[3][DATA][18] , \chs_in_f[3][DATA][17] ,
         \chs_in_f[3][DATA][16] , \chs_in_f[3][DATA][15] ,
         \chs_in_f[3][DATA][14] , \chs_in_f[3][DATA][13] ,
         \chs_in_f[3][DATA][12] , \chs_in_f[3][DATA][11] ,
         \chs_in_f[3][DATA][10] , \chs_in_f[3][DATA][9] ,
         \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] ,
         \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] ,
         \chs_in_f[3][DATA][4] , \chs_in_f[3][DATA][3] ,
         \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] ,
         \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] ,
         \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] ,
         \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] ,
         \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] ,
         \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] ,
         \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] ,
         \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] ,
         \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] ,
         \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] ,
         \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] ,
         \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] ,
         \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] ,
         \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] ,
         \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] ,
         \chs_in_f[2][DATA][7] , \chs_in_f[2][DATA][6] ,
         \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] ,
         \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] ,
         \chs_in_f[2][DATA][1] , \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] ,
         \chs_in_f[1][DATA][34] , \chs_in_f[1][DATA][33] ,
         \chs_in_f[1][DATA][32] , \chs_in_f[1][DATA][31] ,
         \chs_in_f[1][DATA][30] , \chs_in_f[1][DATA][29] ,
         \chs_in_f[1][DATA][28] , \chs_in_f[1][DATA][27] ,
         \chs_in_f[1][DATA][26] , \chs_in_f[1][DATA][25] ,
         \chs_in_f[1][DATA][24] , \chs_in_f[1][DATA][23] ,
         \chs_in_f[1][DATA][22] , \chs_in_f[1][DATA][21] ,
         \chs_in_f[1][DATA][20] , \chs_in_f[1][DATA][19] ,
         \chs_in_f[1][DATA][18] , \chs_in_f[1][DATA][17] ,
         \chs_in_f[1][DATA][16] , \chs_in_f[1][DATA][15] ,
         \chs_in_f[1][DATA][14] , \chs_in_f[1][DATA][13] ,
         \chs_in_f[1][DATA][12] , \chs_in_f[1][DATA][11] ,
         \chs_in_f[1][DATA][10] , \chs_in_f[1][DATA][9] ,
         \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] ,
         \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] ,
         \chs_in_f[1][DATA][4] , \chs_in_f[1][DATA][3] ,
         \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] ,
         \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] ,
         \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] ,
         \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] ,
         \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] ,
         \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] ,
         \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] ,
         \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] ,
         \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] ,
         \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] ,
         \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] ,
         \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] ,
         \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] ,
         \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] ,
         \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] ,
         \chs_in_f[0][DATA][7] , \chs_in_f[0][DATA][6] ,
         \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] ,
         \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] ,
         \chs_in_f[0][DATA][1] , \chs_in_f[0][DATA][0] , \chs_out_b[4][ACK] ,
         \chs_out_b[3][ACK] , \chs_out_b[2][ACK] , \chs_out_b[1][ACK] ,
         \chs_out_b[0][ACK] ;
  output \chs_in_b[4][ACK] , \chs_in_b[3][ACK] , \chs_in_b[2][ACK] ,
         \chs_in_b[1][ACK] , \chs_in_b[0][ACK] , \chs_out_f[4][REQ] ,
         \chs_out_f[4][DATA][34] , \chs_out_f[4][DATA][33] ,
         \chs_out_f[4][DATA][32] , \chs_out_f[4][DATA][31] ,
         \chs_out_f[4][DATA][30] , \chs_out_f[4][DATA][29] ,
         \chs_out_f[4][DATA][28] , \chs_out_f[4][DATA][27] ,
         \chs_out_f[4][DATA][26] , \chs_out_f[4][DATA][25] ,
         \chs_out_f[4][DATA][24] , \chs_out_f[4][DATA][23] ,
         \chs_out_f[4][DATA][22] , \chs_out_f[4][DATA][21] ,
         \chs_out_f[4][DATA][20] , \chs_out_f[4][DATA][19] ,
         \chs_out_f[4][DATA][18] , \chs_out_f[4][DATA][17] ,
         \chs_out_f[4][DATA][16] , \chs_out_f[4][DATA][15] ,
         \chs_out_f[4][DATA][14] , \chs_out_f[4][DATA][13] ,
         \chs_out_f[4][DATA][12] , \chs_out_f[4][DATA][11] ,
         \chs_out_f[4][DATA][10] , \chs_out_f[4][DATA][9] ,
         \chs_out_f[4][DATA][8] , \chs_out_f[4][DATA][7] ,
         \chs_out_f[4][DATA][6] , \chs_out_f[4][DATA][5] ,
         \chs_out_f[4][DATA][4] , \chs_out_f[4][DATA][3] ,
         \chs_out_f[4][DATA][2] , \chs_out_f[4][DATA][1] ,
         \chs_out_f[4][DATA][0] , \chs_out_f[3][REQ] ,
         \chs_out_f[3][DATA][34] , \chs_out_f[3][DATA][33] ,
         \chs_out_f[3][DATA][32] , \chs_out_f[3][DATA][31] ,
         \chs_out_f[3][DATA][30] , \chs_out_f[3][DATA][29] ,
         \chs_out_f[3][DATA][28] , \chs_out_f[3][DATA][27] ,
         \chs_out_f[3][DATA][26] , \chs_out_f[3][DATA][25] ,
         \chs_out_f[3][DATA][24] , \chs_out_f[3][DATA][23] ,
         \chs_out_f[3][DATA][22] , \chs_out_f[3][DATA][21] ,
         \chs_out_f[3][DATA][20] , \chs_out_f[3][DATA][19] ,
         \chs_out_f[3][DATA][18] , \chs_out_f[3][DATA][17] ,
         \chs_out_f[3][DATA][16] , \chs_out_f[3][DATA][15] ,
         \chs_out_f[3][DATA][14] , \chs_out_f[3][DATA][13] ,
         \chs_out_f[3][DATA][12] , \chs_out_f[3][DATA][11] ,
         \chs_out_f[3][DATA][10] , \chs_out_f[3][DATA][9] ,
         \chs_out_f[3][DATA][8] , \chs_out_f[3][DATA][7] ,
         \chs_out_f[3][DATA][6] , \chs_out_f[3][DATA][5] ,
         \chs_out_f[3][DATA][4] , \chs_out_f[3][DATA][3] ,
         \chs_out_f[3][DATA][2] , \chs_out_f[3][DATA][1] ,
         \chs_out_f[3][DATA][0] , \chs_out_f[2][REQ] ,
         \chs_out_f[2][DATA][34] , \chs_out_f[2][DATA][33] ,
         \chs_out_f[2][DATA][32] , \chs_out_f[2][DATA][31] ,
         \chs_out_f[2][DATA][30] , \chs_out_f[2][DATA][29] ,
         \chs_out_f[2][DATA][28] , \chs_out_f[2][DATA][27] ,
         \chs_out_f[2][DATA][26] , \chs_out_f[2][DATA][25] ,
         \chs_out_f[2][DATA][24] , \chs_out_f[2][DATA][23] ,
         \chs_out_f[2][DATA][22] , \chs_out_f[2][DATA][21] ,
         \chs_out_f[2][DATA][20] , \chs_out_f[2][DATA][19] ,
         \chs_out_f[2][DATA][18] , \chs_out_f[2][DATA][17] ,
         \chs_out_f[2][DATA][16] , \chs_out_f[2][DATA][15] ,
         \chs_out_f[2][DATA][14] , \chs_out_f[2][DATA][13] ,
         \chs_out_f[2][DATA][12] , \chs_out_f[2][DATA][11] ,
         \chs_out_f[2][DATA][10] , \chs_out_f[2][DATA][9] ,
         \chs_out_f[2][DATA][8] , \chs_out_f[2][DATA][7] ,
         \chs_out_f[2][DATA][6] , \chs_out_f[2][DATA][5] ,
         \chs_out_f[2][DATA][4] , \chs_out_f[2][DATA][3] ,
         \chs_out_f[2][DATA][2] , \chs_out_f[2][DATA][1] ,
         \chs_out_f[2][DATA][0] , \chs_out_f[1][REQ] ,
         \chs_out_f[1][DATA][34] , \chs_out_f[1][DATA][33] ,
         \chs_out_f[1][DATA][32] , \chs_out_f[1][DATA][31] ,
         \chs_out_f[1][DATA][30] , \chs_out_f[1][DATA][29] ,
         \chs_out_f[1][DATA][28] , \chs_out_f[1][DATA][27] ,
         \chs_out_f[1][DATA][26] , \chs_out_f[1][DATA][25] ,
         \chs_out_f[1][DATA][24] , \chs_out_f[1][DATA][23] ,
         \chs_out_f[1][DATA][22] , \chs_out_f[1][DATA][21] ,
         \chs_out_f[1][DATA][20] , \chs_out_f[1][DATA][19] ,
         \chs_out_f[1][DATA][18] , \chs_out_f[1][DATA][17] ,
         \chs_out_f[1][DATA][16] , \chs_out_f[1][DATA][15] ,
         \chs_out_f[1][DATA][14] , \chs_out_f[1][DATA][13] ,
         \chs_out_f[1][DATA][12] , \chs_out_f[1][DATA][11] ,
         \chs_out_f[1][DATA][10] , \chs_out_f[1][DATA][9] ,
         \chs_out_f[1][DATA][8] , \chs_out_f[1][DATA][7] ,
         \chs_out_f[1][DATA][6] , \chs_out_f[1][DATA][5] ,
         \chs_out_f[1][DATA][4] , \chs_out_f[1][DATA][3] ,
         \chs_out_f[1][DATA][2] , \chs_out_f[1][DATA][1] ,
         \chs_out_f[1][DATA][0] , \chs_out_f[0][REQ] ,
         \chs_out_f[0][DATA][34] , \chs_out_f[0][DATA][33] ,
         \chs_out_f[0][DATA][32] , \chs_out_f[0][DATA][31] ,
         \chs_out_f[0][DATA][30] , \chs_out_f[0][DATA][29] ,
         \chs_out_f[0][DATA][28] , \chs_out_f[0][DATA][27] ,
         \chs_out_f[0][DATA][26] , \chs_out_f[0][DATA][25] ,
         \chs_out_f[0][DATA][24] , \chs_out_f[0][DATA][23] ,
         \chs_out_f[0][DATA][22] , \chs_out_f[0][DATA][21] ,
         \chs_out_f[0][DATA][20] , \chs_out_f[0][DATA][19] ,
         \chs_out_f[0][DATA][18] , \chs_out_f[0][DATA][17] ,
         \chs_out_f[0][DATA][16] , \chs_out_f[0][DATA][15] ,
         \chs_out_f[0][DATA][14] , \chs_out_f[0][DATA][13] ,
         \chs_out_f[0][DATA][12] , \chs_out_f[0][DATA][11] ,
         \chs_out_f[0][DATA][10] , \chs_out_f[0][DATA][9] ,
         \chs_out_f[0][DATA][8] , \chs_out_f[0][DATA][7] ,
         \chs_out_f[0][DATA][6] , \chs_out_f[0][DATA][5] ,
         \chs_out_f[0][DATA][4] , \chs_out_f[0][DATA][3] ,
         \chs_out_f[0][DATA][2] , \chs_out_f[0][DATA][1] ,
         \chs_out_f[0][DATA][0] ;
  wire   \chs_in_b[4][ACK] , \chs_out_f[4][REQ] , synced_req, del, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510;
  assign \chs_in_b[0][ACK]  = \chs_in_b[4][ACK] ;
  assign \chs_in_b[1][ACK]  = \chs_in_b[4][ACK] ;
  assign \chs_in_b[2][ACK]  = \chs_in_b[4][ACK] ;
  assign \chs_in_b[3][ACK]  = \chs_in_b[4][ACK] ;
  assign \chs_out_f[0][REQ]  = \chs_out_f[4][REQ] ;
  assign \chs_out_f[1][REQ]  = \chs_out_f[4][REQ] ;
  assign \chs_out_f[2][REQ]  = \chs_out_f[4][REQ] ;
  assign \chs_out_f[3][REQ]  = \chs_out_f[4][REQ] ;

  c_gate_generic_1_5_2 c_sync_req ( .preset(preset), .\input ({
        \chs_in_f[4][REQ] , \chs_in_f[3][REQ] , \chs_in_f[2][REQ] , 
        \chs_in_f[1][REQ] , \chs_in_f[0][REQ] }), .\output (synced_req) );
  c_gate_generic_1_5_1 c_sync_ack ( .preset(preset), .\input ({
        \chs_out_b[4][ACK] , \chs_out_b[3][ACK] , \chs_out_b[2][ACK] , 
        \chs_out_b[1][ACK] , \chs_out_b[0][ACK] }), .\output (
        \chs_in_b[4][ACK] ) );
  HS65_LS_IVX9 I_1 ( .A(n1), .Z(\chs_out_f[4][REQ] ) );
  HS65_LH_IVX2 I_0 ( .A(synced_req), .Z(del) );
  HS65_LS_IVX9 U2 ( .A(\switch_sel[3][4] ), .Z(n261) );
  HS65_LS_IVX9 U3 ( .A(\switch_sel[3][2] ), .Z(n262) );
  HS65_LS_IVX9 U4 ( .A(\switch_sel[3][1] ), .Z(n263) );
  HS65_LS_IVX9 U5 ( .A(\switch_sel[3][0] ), .Z(n264) );
  HS65_LS_BFX9 U6 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U7 ( .A(del), .Z(n2) );
  HS65_LS_BFX9 U8 ( .A(n258), .Z(n10) );
  HS65_LS_BFX9 U9 ( .A(n257), .Z(n8) );
  HS65_LS_BFX9 U10 ( .A(n256), .Z(n5) );
  HS65_LS_BFX7 U11 ( .A(n259), .Z(n12) );
  HS65_LS_BFX7 U12 ( .A(n259), .Z(n13) );
  HS65_LS_BFX9 U13 ( .A(\switch_sel[0][4] ), .Z(n45) );
  HS65_LS_BFX9 U14 ( .A(\switch_sel[1][4] ), .Z(n61) );
  HS65_LS_BFX9 U15 ( .A(\switch_sel[0][3] ), .Z(n41) );
  HS65_LS_BFX9 U16 ( .A(\switch_sel[1][3] ), .Z(n57) );
  HS65_LS_BFX9 U17 ( .A(\switch_sel[1][2] ), .Z(n53) );
  HS65_LS_BFX9 U18 ( .A(\switch_sel[0][1] ), .Z(n33) );
  HS65_LS_BFX9 U19 ( .A(\switch_sel[1][0] ), .Z(n49) );
  HS65_LS_BFX9 U20 ( .A(n261), .Z(n18) );
  HS65_LS_BFX9 U21 ( .A(n261), .Z(n19) );
  HS65_LS_BFX9 U22 ( .A(n61), .Z(n62) );
  HS65_LS_BFX9 U23 ( .A(n61), .Z(n63) );
  HS65_LS_BFX9 U24 ( .A(n77), .Z(n78) );
  HS65_LS_BFX9 U25 ( .A(n77), .Z(n79) );
  HS65_LS_BFX9 U26 ( .A(n45), .Z(n46) );
  HS65_LS_BFX9 U27 ( .A(n45), .Z(n47) );
  HS65_LS_BFX9 U28 ( .A(n262), .Z(n21) );
  HS65_LS_BFX9 U29 ( .A(n262), .Z(n22) );
  HS65_LS_BFX9 U30 ( .A(n263), .Z(n24) );
  HS65_LS_BFX9 U31 ( .A(n263), .Z(n25) );
  HS65_LS_BFX9 U32 ( .A(n264), .Z(n27) );
  HS65_LS_BFX9 U33 ( .A(n264), .Z(n28) );
  HS65_LS_BFX9 U34 ( .A(n57), .Z(n58) );
  HS65_LS_BFX9 U35 ( .A(n57), .Z(n59) );
  HS65_LS_BFX9 U36 ( .A(n53), .Z(n54) );
  HS65_LS_BFX9 U37 ( .A(n53), .Z(n55) );
  HS65_LS_BFX9 U38 ( .A(n49), .Z(n50) );
  HS65_LS_BFX9 U39 ( .A(n49), .Z(n51) );
  HS65_LS_BFX9 U40 ( .A(n73), .Z(n74) );
  HS65_LS_BFX9 U41 ( .A(n73), .Z(n75) );
  HS65_LS_BFX9 U42 ( .A(n69), .Z(n70) );
  HS65_LS_BFX9 U43 ( .A(n69), .Z(n71) );
  HS65_LS_BFX9 U44 ( .A(n65), .Z(n66) );
  HS65_LS_BFX9 U45 ( .A(n65), .Z(n67) );
  HS65_LS_BFX9 U46 ( .A(n261), .Z(n20) );
  HS65_LS_BFX9 U47 ( .A(n41), .Z(n42) );
  HS65_LS_BFX9 U48 ( .A(n41), .Z(n43) );
  HS65_LS_BFX9 U49 ( .A(n37), .Z(n38) );
  HS65_LS_BFX9 U50 ( .A(n37), .Z(n39) );
  HS65_LS_BFX9 U51 ( .A(n33), .Z(n34) );
  HS65_LS_BFX9 U52 ( .A(n33), .Z(n35) );
  HS65_LS_BFX9 U53 ( .A(n45), .Z(n48) );
  HS65_LS_BFX9 U54 ( .A(n256), .Z(n3) );
  HS65_LS_BFX9 U55 ( .A(n256), .Z(n4) );
  HS65_LS_BFX9 U56 ( .A(n257), .Z(n6) );
  HS65_LS_BFX9 U57 ( .A(n257), .Z(n7) );
  HS65_LS_BFX9 U58 ( .A(n258), .Z(n9) );
  HS65_LS_BFX9 U59 ( .A(n57), .Z(n60) );
  HS65_LS_BFX9 U60 ( .A(n53), .Z(n56) );
  HS65_LS_BFX9 U61 ( .A(n49), .Z(n52) );
  HS65_LS_BFX9 U62 ( .A(n73), .Z(n76) );
  HS65_LS_BFX9 U63 ( .A(n69), .Z(n72) );
  HS65_LS_BFX9 U64 ( .A(n65), .Z(n68) );
  HS65_LS_BFX9 U65 ( .A(n41), .Z(n44) );
  HS65_LS_BFX9 U66 ( .A(n37), .Z(n40) );
  HS65_LS_BFX9 U67 ( .A(n33), .Z(n36) );
  HS65_LS_BFX9 U68 ( .A(n258), .Z(n11) );
  HS65_LS_BFX9 U69 ( .A(n259), .Z(n14) );
  HS65_LS_BFX9 U70 ( .A(n262), .Z(n23) );
  HS65_LS_BFX9 U71 ( .A(n263), .Z(n26) );
  HS65_LS_BFX9 U72 ( .A(n264), .Z(n29) );
  HS65_LS_BFX9 U73 ( .A(n61), .Z(n64) );
  HS65_LS_BFX9 U74 ( .A(n77), .Z(n80) );
  HS65_LS_BFX9 U75 ( .A(n260), .Z(n15) );
  HS65_LS_BFX9 U76 ( .A(n260), .Z(n16) );
  HS65_LS_BFX9 U77 ( .A(n265), .Z(n30) );
  HS65_LS_BFX9 U78 ( .A(n265), .Z(n31) );
  HS65_LS_BFX9 U79 ( .A(n260), .Z(n17) );
  HS65_LS_BFX9 U80 ( .A(n265), .Z(n32) );
  HS65_LS_IVX9 U81 ( .A(\switch_sel[4][0] ), .Z(n259) );
  HS65_LS_IVX9 U82 ( .A(\switch_sel[4][2] ), .Z(n257) );
  HS65_LS_IVX9 U83 ( .A(\switch_sel[4][1] ), .Z(n258) );
  HS65_LS_IVX9 U84 ( .A(\switch_sel[4][3] ), .Z(n256) );
  HS65_LS_AOI222X2 U85 ( .A(\chs_in_f[2][DATA][34] ), .B(n78), .C(
        \chs_in_f[0][DATA][34] ), .D(n48), .E(\chs_in_f[1][DATA][34] ), .F(n62), .Z(n503) );
  HS65_LS_OAI212X5 U86 ( .A(n291), .B(n20), .C(n326), .D(n17), .E(n510), .Z(
        \chs_out_f[4][DATA][9] ) );
  HS65_LS_AOI222X2 U87 ( .A(n78), .B(\chs_in_f[2][DATA][9] ), .C(n48), .D(
        \chs_in_f[0][DATA][9] ), .E(n62), .F(\chs_in_f[1][DATA][9] ), .Z(n510)
         );
  HS65_LS_AOI222X2 U88 ( .A(n76), .B(\chs_in_f[2][DATA][34] ), .C(n44), .D(
        \chs_in_f[0][DATA][34] ), .E(n60), .F(\chs_in_f[1][DATA][34] ), .Z(
        n468) );
  HS65_LS_AOI222X2 U89 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][34] ), 
        .C(n40), .D(\chs_in_f[0][DATA][34] ), .E(n56), .F(
        \chs_in_f[1][DATA][34] ), .Z(n433) );
  HS65_LS_AOI222X2 U90 ( .A(n72), .B(\chs_in_f[2][DATA][34] ), .C(n36), .D(
        \chs_in_f[0][DATA][34] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][34] ), .Z(n398) );
  HS65_LS_AOI222X2 U91 ( .A(n68), .B(\chs_in_f[2][DATA][34] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][34] ), .E(n52), .F(
        \chs_in_f[1][DATA][34] ), .Z(n363) );
  HS65_LS_IVX9 U92 ( .A(\chs_in_f[3][DATA][9] ), .Z(n291) );
  HS65_LS_IVX9 U93 ( .A(\chs_in_f[3][DATA][34] ), .Z(n266) );
  HS65_LS_IVX9 U94 ( .A(\chs_in_f[3][DATA][0] ), .Z(n300) );
  HS65_LS_IVX9 U95 ( .A(\chs_in_f[3][DATA][1] ), .Z(n299) );
  HS65_LS_IVX9 U96 ( .A(\chs_in_f[3][DATA][2] ), .Z(n298) );
  HS65_LS_IVX9 U97 ( .A(\chs_in_f[3][DATA][3] ), .Z(n297) );
  HS65_LS_IVX9 U98 ( .A(\chs_in_f[3][DATA][4] ), .Z(n296) );
  HS65_LS_IVX9 U99 ( .A(\chs_in_f[3][DATA][5] ), .Z(n295) );
  HS65_LS_IVX9 U100 ( .A(\chs_in_f[3][DATA][6] ), .Z(n294) );
  HS65_LS_IVX9 U101 ( .A(\chs_in_f[3][DATA][7] ), .Z(n293) );
  HS65_LS_IVX9 U102 ( .A(\chs_in_f[3][DATA][8] ), .Z(n292) );
  HS65_LS_IVX9 U103 ( .A(\chs_in_f[3][DATA][10] ), .Z(n290) );
  HS65_LS_IVX9 U104 ( .A(\chs_in_f[3][DATA][11] ), .Z(n289) );
  HS65_LS_IVX9 U105 ( .A(\chs_in_f[3][DATA][12] ), .Z(n288) );
  HS65_LS_IVX9 U106 ( .A(\chs_in_f[3][DATA][13] ), .Z(n287) );
  HS65_LS_IVX9 U107 ( .A(\chs_in_f[3][DATA][14] ), .Z(n286) );
  HS65_LS_IVX9 U108 ( .A(\chs_in_f[3][DATA][15] ), .Z(n285) );
  HS65_LS_IVX9 U109 ( .A(\chs_in_f[3][DATA][16] ), .Z(n284) );
  HS65_LS_IVX9 U110 ( .A(\chs_in_f[3][DATA][17] ), .Z(n283) );
  HS65_LS_IVX9 U111 ( .A(\chs_in_f[3][DATA][18] ), .Z(n282) );
  HS65_LS_IVX9 U112 ( .A(\chs_in_f[3][DATA][19] ), .Z(n281) );
  HS65_LS_IVX9 U113 ( .A(\chs_in_f[3][DATA][20] ), .Z(n280) );
  HS65_LS_IVX9 U114 ( .A(\chs_in_f[3][DATA][21] ), .Z(n279) );
  HS65_LS_IVX9 U115 ( .A(\chs_in_f[3][DATA][22] ), .Z(n278) );
  HS65_LS_IVX9 U116 ( .A(\chs_in_f[3][DATA][23] ), .Z(n277) );
  HS65_LS_IVX9 U117 ( .A(\chs_in_f[3][DATA][24] ), .Z(n276) );
  HS65_LS_IVX9 U118 ( .A(\chs_in_f[3][DATA][25] ), .Z(n275) );
  HS65_LS_IVX9 U119 ( .A(\chs_in_f[3][DATA][26] ), .Z(n274) );
  HS65_LS_IVX9 U120 ( .A(\chs_in_f[3][DATA][27] ), .Z(n273) );
  HS65_LS_IVX9 U121 ( .A(\chs_in_f[3][DATA][28] ), .Z(n272) );
  HS65_LS_IVX9 U122 ( .A(\chs_in_f[3][DATA][29] ), .Z(n271) );
  HS65_LS_IVX9 U123 ( .A(\chs_in_f[3][DATA][30] ), .Z(n270) );
  HS65_LS_IVX9 U124 ( .A(\chs_in_f[3][DATA][31] ), .Z(n269) );
  HS65_LS_IVX9 U125 ( .A(\chs_in_f[3][DATA][32] ), .Z(n268) );
  HS65_LS_IVX9 U126 ( .A(\chs_in_f[3][DATA][33] ), .Z(n267) );
  HS65_LS_IVX9 U127 ( .A(\chs_in_f[4][DATA][9] ), .Z(n326) );
  HS65_LS_IVX9 U128 ( .A(\chs_in_f[4][DATA][34] ), .Z(n301) );
  HS65_LS_IVX9 U129 ( .A(\chs_in_f[4][DATA][0] ), .Z(n335) );
  HS65_LS_IVX9 U130 ( .A(\chs_in_f[4][DATA][1] ), .Z(n334) );
  HS65_LS_IVX9 U131 ( .A(\chs_in_f[4][DATA][2] ), .Z(n333) );
  HS65_LS_IVX9 U132 ( .A(\chs_in_f[4][DATA][3] ), .Z(n332) );
  HS65_LS_IVX9 U133 ( .A(\chs_in_f[4][DATA][4] ), .Z(n331) );
  HS65_LS_IVX9 U134 ( .A(\chs_in_f[4][DATA][5] ), .Z(n330) );
  HS65_LS_IVX9 U135 ( .A(\chs_in_f[4][DATA][6] ), .Z(n329) );
  HS65_LS_IVX9 U136 ( .A(\chs_in_f[4][DATA][7] ), .Z(n328) );
  HS65_LS_IVX9 U137 ( .A(\chs_in_f[4][DATA][8] ), .Z(n327) );
  HS65_LS_IVX9 U138 ( .A(\chs_in_f[4][DATA][10] ), .Z(n325) );
  HS65_LS_IVX9 U139 ( .A(\chs_in_f[4][DATA][11] ), .Z(n324) );
  HS65_LS_IVX9 U140 ( .A(\chs_in_f[4][DATA][12] ), .Z(n323) );
  HS65_LS_IVX9 U141 ( .A(\chs_in_f[4][DATA][13] ), .Z(n322) );
  HS65_LS_IVX9 U142 ( .A(\chs_in_f[4][DATA][14] ), .Z(n321) );
  HS65_LS_IVX9 U143 ( .A(\chs_in_f[4][DATA][15] ), .Z(n320) );
  HS65_LS_IVX9 U144 ( .A(\chs_in_f[4][DATA][16] ), .Z(n319) );
  HS65_LS_IVX9 U145 ( .A(\chs_in_f[4][DATA][17] ), .Z(n318) );
  HS65_LS_IVX9 U146 ( .A(\chs_in_f[4][DATA][18] ), .Z(n317) );
  HS65_LS_IVX9 U147 ( .A(\chs_in_f[4][DATA][19] ), .Z(n316) );
  HS65_LS_IVX9 U148 ( .A(\chs_in_f[4][DATA][20] ), .Z(n315) );
  HS65_LS_IVX9 U149 ( .A(\chs_in_f[4][DATA][21] ), .Z(n314) );
  HS65_LS_IVX9 U150 ( .A(\chs_in_f[4][DATA][22] ), .Z(n313) );
  HS65_LS_IVX9 U151 ( .A(\chs_in_f[4][DATA][23] ), .Z(n312) );
  HS65_LS_IVX9 U152 ( .A(\chs_in_f[4][DATA][24] ), .Z(n311) );
  HS65_LS_IVX9 U153 ( .A(\chs_in_f[4][DATA][25] ), .Z(n310) );
  HS65_LS_IVX9 U154 ( .A(\chs_in_f[4][DATA][26] ), .Z(n309) );
  HS65_LS_IVX9 U155 ( .A(\chs_in_f[4][DATA][27] ), .Z(n308) );
  HS65_LS_IVX9 U156 ( .A(\chs_in_f[4][DATA][28] ), .Z(n307) );
  HS65_LS_IVX9 U157 ( .A(\chs_in_f[4][DATA][29] ), .Z(n306) );
  HS65_LS_IVX9 U158 ( .A(\chs_in_f[4][DATA][30] ), .Z(n305) );
  HS65_LS_IVX9 U159 ( .A(\chs_in_f[4][DATA][31] ), .Z(n304) );
  HS65_LS_IVX9 U160 ( .A(\chs_in_f[4][DATA][32] ), .Z(n303) );
  HS65_LS_IVX9 U161 ( .A(\chs_in_f[4][DATA][33] ), .Z(n302) );
  HS65_LS_BFX18 U162 ( .A(\switch_sel[2][4] ), .Z(n77) );
  HS65_LS_BFX18 U163 ( .A(\switch_sel[2][3] ), .Z(n73) );
  HS65_LS_BFX18 U164 ( .A(\switch_sel[0][2] ), .Z(n37) );
  HS65_LS_BFX18 U165 ( .A(\switch_sel[2][1] ), .Z(n69) );
  HS65_LS_BFX18 U166 ( .A(\switch_sel[2][0] ), .Z(n65) );
  HS65_LS_OAI212X5 U167 ( .A(n18), .B(n300), .C(n15), .D(n335), .E(n476), .Z(
        \chs_out_f[4][DATA][0] ) );
  HS65_LS_AOI222X2 U168 ( .A(\chs_in_f[2][DATA][0] ), .B(n80), .C(
        \chs_in_f[0][DATA][0] ), .D(n46), .E(\chs_in_f[1][DATA][0] ), .F(n64), 
        .Z(n476) );
  HS65_LS_OAI212X5 U169 ( .A(n18), .B(n299), .C(n15), .D(n334), .E(n487), .Z(
        \chs_out_f[4][DATA][1] ) );
  HS65_LS_AOI222X2 U170 ( .A(\chs_in_f[2][DATA][1] ), .B(n79), .C(
        \chs_in_f[0][DATA][1] ), .D(n46), .E(\chs_in_f[1][DATA][1] ), .F(n63), 
        .Z(n487) );
  HS65_LS_OAI212X5 U171 ( .A(n19), .B(n298), .C(n16), .D(n333), .E(n498), .Z(
        \chs_out_f[4][DATA][2] ) );
  HS65_LS_AOI222X2 U172 ( .A(\chs_in_f[2][DATA][2] ), .B(n78), .C(
        \chs_in_f[0][DATA][2] ), .D(n47), .E(\chs_in_f[1][DATA][2] ), .F(n62), 
        .Z(n498) );
  HS65_LS_OAI212X5 U173 ( .A(n20), .B(n297), .C(n17), .D(n332), .E(n504), .Z(
        \chs_out_f[4][DATA][3] ) );
  HS65_LS_AOI222X2 U174 ( .A(\chs_in_f[2][DATA][3] ), .B(n78), .C(
        \chs_in_f[0][DATA][3] ), .D(n48), .E(\chs_in_f[1][DATA][3] ), .F(n62), 
        .Z(n504) );
  HS65_LS_OAI212X5 U175 ( .A(n20), .B(n296), .C(n17), .D(n331), .E(n505), .Z(
        \chs_out_f[4][DATA][4] ) );
  HS65_LS_AOI222X2 U176 ( .A(\chs_in_f[2][DATA][4] ), .B(n78), .C(
        \chs_in_f[0][DATA][4] ), .D(n48), .E(\chs_in_f[1][DATA][4] ), .F(n62), 
        .Z(n505) );
  HS65_LS_OAI212X5 U177 ( .A(n20), .B(n295), .C(n17), .D(n330), .E(n506), .Z(
        \chs_out_f[4][DATA][5] ) );
  HS65_LS_AOI222X2 U178 ( .A(\chs_in_f[2][DATA][5] ), .B(n78), .C(
        \chs_in_f[0][DATA][5] ), .D(n48), .E(\chs_in_f[1][DATA][5] ), .F(n62), 
        .Z(n506) );
  HS65_LS_OAI212X5 U179 ( .A(n20), .B(n294), .C(n17), .D(n329), .E(n507), .Z(
        \chs_out_f[4][DATA][6] ) );
  HS65_LS_AOI222X2 U180 ( .A(\chs_in_f[2][DATA][6] ), .B(n78), .C(
        \chs_in_f[0][DATA][6] ), .D(n48), .E(\chs_in_f[1][DATA][6] ), .F(n62), 
        .Z(n507) );
  HS65_LS_OAI212X5 U181 ( .A(n20), .B(n293), .C(n17), .D(n328), .E(n508), .Z(
        \chs_out_f[4][DATA][7] ) );
  HS65_LS_AOI222X2 U182 ( .A(\chs_in_f[2][DATA][7] ), .B(n78), .C(
        \chs_in_f[0][DATA][7] ), .D(n48), .E(\chs_in_f[1][DATA][7] ), .F(n62), 
        .Z(n508) );
  HS65_LS_OAI212X5 U183 ( .A(n20), .B(n292), .C(n17), .D(n327), .E(n509), .Z(
        \chs_out_f[4][DATA][8] ) );
  HS65_LS_AOI222X2 U184 ( .A(\chs_in_f[2][DATA][8] ), .B(n78), .C(
        \chs_in_f[0][DATA][8] ), .D(n48), .E(\chs_in_f[1][DATA][8] ), .F(n62), 
        .Z(n509) );
  HS65_LS_OAI212X5 U185 ( .A(n18), .B(n290), .C(n15), .D(n325), .E(n477), .Z(
        \chs_out_f[4][DATA][10] ) );
  HS65_LS_AOI222X2 U186 ( .A(\chs_in_f[2][DATA][10] ), .B(n80), .C(
        \chs_in_f[0][DATA][10] ), .D(n46), .E(\chs_in_f[1][DATA][10] ), .F(n64), .Z(n477) );
  HS65_LS_OAI212X5 U187 ( .A(n18), .B(n289), .C(n15), .D(n324), .E(n478), .Z(
        \chs_out_f[4][DATA][11] ) );
  HS65_LS_AOI222X2 U188 ( .A(\chs_in_f[2][DATA][11] ), .B(n80), .C(
        \chs_in_f[0][DATA][11] ), .D(n46), .E(\chs_in_f[1][DATA][11] ), .F(n64), .Z(n478) );
  HS65_LS_OAI212X5 U189 ( .A(n18), .B(n288), .C(n15), .D(n323), .E(n479), .Z(
        \chs_out_f[4][DATA][12] ) );
  HS65_LS_AOI222X2 U190 ( .A(\chs_in_f[2][DATA][12] ), .B(n80), .C(
        \chs_in_f[0][DATA][12] ), .D(n46), .E(\chs_in_f[1][DATA][12] ), .F(n64), .Z(n479) );
  HS65_LS_OAI212X5 U191 ( .A(n18), .B(n287), .C(n15), .D(n322), .E(n480), .Z(
        \chs_out_f[4][DATA][13] ) );
  HS65_LS_AOI222X2 U192 ( .A(\chs_in_f[2][DATA][13] ), .B(n80), .C(
        \chs_in_f[0][DATA][13] ), .D(n46), .E(\chs_in_f[1][DATA][13] ), .F(n64), .Z(n480) );
  HS65_LS_OAI212X5 U193 ( .A(n18), .B(n286), .C(n15), .D(n321), .E(n481), .Z(
        \chs_out_f[4][DATA][14] ) );
  HS65_LS_AOI222X2 U194 ( .A(\chs_in_f[2][DATA][14] ), .B(n80), .C(
        \chs_in_f[0][DATA][14] ), .D(n46), .E(\chs_in_f[1][DATA][14] ), .F(n64), .Z(n481) );
  HS65_LS_OAI212X5 U195 ( .A(n18), .B(n285), .C(n15), .D(n320), .E(n482), .Z(
        \chs_out_f[4][DATA][15] ) );
  HS65_LS_AOI222X2 U196 ( .A(\chs_in_f[2][DATA][15] ), .B(n80), .C(
        \chs_in_f[0][DATA][15] ), .D(n46), .E(\chs_in_f[1][DATA][15] ), .F(n64), .Z(n482) );
  HS65_LS_OAI212X5 U197 ( .A(n18), .B(n284), .C(n15), .D(n319), .E(n483), .Z(
        \chs_out_f[4][DATA][16] ) );
  HS65_LS_AOI222X2 U198 ( .A(\chs_in_f[2][DATA][16] ), .B(n80), .C(
        \chs_in_f[0][DATA][16] ), .D(n46), .E(\chs_in_f[1][DATA][16] ), .F(n64), .Z(n483) );
  HS65_LS_OAI212X5 U199 ( .A(n18), .B(n283), .C(n15), .D(n318), .E(n484), .Z(
        \chs_out_f[4][DATA][17] ) );
  HS65_LS_AOI222X2 U200 ( .A(\chs_in_f[2][DATA][17] ), .B(n80), .C(
        \chs_in_f[0][DATA][17] ), .D(n46), .E(\chs_in_f[1][DATA][17] ), .F(n64), .Z(n484) );
  HS65_LS_OAI212X5 U201 ( .A(n18), .B(n282), .C(n15), .D(n317), .E(n485), .Z(
        \chs_out_f[4][DATA][18] ) );
  HS65_LS_AOI222X2 U202 ( .A(\chs_in_f[2][DATA][18] ), .B(n79), .C(
        \chs_in_f[0][DATA][18] ), .D(n46), .E(\chs_in_f[1][DATA][18] ), .F(n63), .Z(n485) );
  HS65_LS_OAI212X5 U203 ( .A(n18), .B(n281), .C(n15), .D(n316), .E(n486), .Z(
        \chs_out_f[4][DATA][19] ) );
  HS65_LS_AOI222X2 U204 ( .A(\chs_in_f[2][DATA][19] ), .B(n79), .C(
        \chs_in_f[0][DATA][19] ), .D(n46), .E(\chs_in_f[1][DATA][19] ), .F(n63), .Z(n486) );
  HS65_LS_OAI212X5 U205 ( .A(n19), .B(n280), .C(n15), .D(n315), .E(n488), .Z(
        \chs_out_f[4][DATA][20] ) );
  HS65_LS_AOI222X2 U206 ( .A(\chs_in_f[2][DATA][20] ), .B(n79), .C(
        \chs_in_f[0][DATA][20] ), .D(n47), .E(\chs_in_f[1][DATA][20] ), .F(n63), .Z(n488) );
  HS65_LS_OAI212X5 U207 ( .A(n19), .B(n279), .C(n16), .D(n314), .E(n489), .Z(
        \chs_out_f[4][DATA][21] ) );
  HS65_LS_AOI222X2 U208 ( .A(\chs_in_f[2][DATA][21] ), .B(n79), .C(
        \chs_in_f[0][DATA][21] ), .D(n47), .E(\chs_in_f[1][DATA][21] ), .F(n63), .Z(n489) );
  HS65_LS_OAI212X5 U209 ( .A(n19), .B(n278), .C(n16), .D(n313), .E(n490), .Z(
        \chs_out_f[4][DATA][22] ) );
  HS65_LS_AOI222X2 U210 ( .A(\chs_in_f[2][DATA][22] ), .B(n79), .C(
        \chs_in_f[0][DATA][22] ), .D(n47), .E(\chs_in_f[1][DATA][22] ), .F(n63), .Z(n490) );
  HS65_LS_OAI212X5 U211 ( .A(n19), .B(n277), .C(n16), .D(n312), .E(n491), .Z(
        \chs_out_f[4][DATA][23] ) );
  HS65_LS_AOI222X2 U212 ( .A(\chs_in_f[2][DATA][23] ), .B(n79), .C(
        \chs_in_f[0][DATA][23] ), .D(n47), .E(\chs_in_f[1][DATA][23] ), .F(n63), .Z(n491) );
  HS65_LS_OAI212X5 U213 ( .A(n19), .B(n276), .C(n16), .D(n311), .E(n492), .Z(
        \chs_out_f[4][DATA][24] ) );
  HS65_LS_AOI222X2 U214 ( .A(\chs_in_f[2][DATA][24] ), .B(n79), .C(
        \chs_in_f[0][DATA][24] ), .D(n47), .E(\chs_in_f[1][DATA][24] ), .F(n63), .Z(n492) );
  HS65_LS_OAI212X5 U215 ( .A(n19), .B(n275), .C(n16), .D(n310), .E(n493), .Z(
        \chs_out_f[4][DATA][25] ) );
  HS65_LS_AOI222X2 U216 ( .A(\chs_in_f[2][DATA][25] ), .B(n79), .C(
        \chs_in_f[0][DATA][25] ), .D(n47), .E(\chs_in_f[1][DATA][25] ), .F(n63), .Z(n493) );
  HS65_LS_OAI212X5 U217 ( .A(n19), .B(n274), .C(n16), .D(n309), .E(n494), .Z(
        \chs_out_f[4][DATA][26] ) );
  HS65_LS_AOI222X2 U218 ( .A(\chs_in_f[2][DATA][26] ), .B(n79), .C(
        \chs_in_f[0][DATA][26] ), .D(n47), .E(\chs_in_f[1][DATA][26] ), .F(n63), .Z(n494) );
  HS65_LS_OAI212X5 U219 ( .A(n19), .B(n273), .C(n16), .D(n308), .E(n495), .Z(
        \chs_out_f[4][DATA][27] ) );
  HS65_LS_AOI222X2 U220 ( .A(\chs_in_f[2][DATA][27] ), .B(n79), .C(
        \chs_in_f[0][DATA][27] ), .D(n47), .E(\chs_in_f[1][DATA][27] ), .F(n63), .Z(n495) );
  HS65_LS_OAI212X5 U221 ( .A(n19), .B(n272), .C(n16), .D(n307), .E(n496), .Z(
        \chs_out_f[4][DATA][28] ) );
  HS65_LS_AOI222X2 U222 ( .A(\chs_in_f[2][DATA][28] ), .B(n79), .C(
        \chs_in_f[0][DATA][28] ), .D(n47), .E(\chs_in_f[1][DATA][28] ), .F(n63), .Z(n496) );
  HS65_LS_OAI212X5 U223 ( .A(n19), .B(n271), .C(n16), .D(n306), .E(n497), .Z(
        \chs_out_f[4][DATA][29] ) );
  HS65_LS_AOI222X2 U224 ( .A(\chs_in_f[2][DATA][29] ), .B(n79), .C(
        \chs_in_f[0][DATA][29] ), .D(n47), .E(\chs_in_f[1][DATA][29] ), .F(n63), .Z(n497) );
  HS65_LS_OAI212X5 U225 ( .A(n19), .B(n270), .C(n16), .D(n305), .E(n499), .Z(
        \chs_out_f[4][DATA][30] ) );
  HS65_LS_AOI222X2 U226 ( .A(\chs_in_f[2][DATA][30] ), .B(n78), .C(
        \chs_in_f[0][DATA][30] ), .D(n47), .E(\chs_in_f[1][DATA][30] ), .F(n62), .Z(n499) );
  HS65_LS_OAI212X5 U227 ( .A(n20), .B(n269), .C(n16), .D(n304), .E(n500), .Z(
        \chs_out_f[4][DATA][31] ) );
  HS65_LS_AOI222X2 U228 ( .A(\chs_in_f[2][DATA][31] ), .B(n78), .C(
        \chs_in_f[0][DATA][31] ), .D(n48), .E(\chs_in_f[1][DATA][31] ), .F(n62), .Z(n500) );
  HS65_LS_OAI212X5 U229 ( .A(n20), .B(n268), .C(n16), .D(n303), .E(n501), .Z(
        \chs_out_f[4][DATA][32] ) );
  HS65_LS_AOI222X2 U230 ( .A(\chs_in_f[2][DATA][32] ), .B(n78), .C(
        \chs_in_f[0][DATA][32] ), .D(n48), .E(\chs_in_f[1][DATA][32] ), .F(n62), .Z(n501) );
  HS65_LS_OAI212X5 U231 ( .A(n20), .B(n267), .C(n17), .D(n302), .E(n502), .Z(
        \chs_out_f[4][DATA][33] ) );
  HS65_LS_AOI222X2 U232 ( .A(\chs_in_f[2][DATA][33] ), .B(n78), .C(
        \chs_in_f[0][DATA][33] ), .D(n48), .E(\chs_in_f[1][DATA][33] ), .F(n62), .Z(n502) );
  HS65_LS_OAI212X5 U233 ( .A(n291), .B(n29), .C(n326), .D(n14), .E(n370), .Z(
        \chs_out_f[0][DATA][9] ) );
  HS65_LS_AOI222X2 U234 ( .A(n68), .B(\chs_in_f[2][DATA][9] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][9] ), .E(n52), .F(
        \chs_in_f[1][DATA][9] ), .Z(n370) );
  HS65_LS_OAI212X5 U235 ( .A(n291), .B(n23), .C(n326), .D(n8), .E(n440), .Z(
        \chs_out_f[2][DATA][9] ) );
  HS65_LS_AOI222X2 U236 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][9] ), 
        .C(n40), .D(\chs_in_f[0][DATA][9] ), .E(n56), .F(
        \chs_in_f[1][DATA][9] ), .Z(n440) );
  HS65_LS_OAI212X5 U237 ( .A(n291), .B(n26), .C(n326), .D(n11), .E(n405), .Z(
        \chs_out_f[1][DATA][9] ) );
  HS65_LS_AOI222X2 U238 ( .A(n72), .B(\chs_in_f[2][DATA][9] ), .C(n36), .D(
        \chs_in_f[0][DATA][9] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][9] ), .Z(n405) );
  HS65_LS_OAI212X5 U239 ( .A(n300), .B(n27), .C(n335), .D(n12), .E(n336), .Z(
        \chs_out_f[0][DATA][0] ) );
  HS65_LS_AOI222X2 U240 ( .A(n66), .B(\chs_in_f[2][DATA][0] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][0] ), .E(n50), .F(
        \chs_in_f[1][DATA][0] ), .Z(n336) );
  HS65_LS_OAI212X5 U241 ( .A(n299), .B(n27), .C(n334), .D(n12), .E(n347), .Z(
        \chs_out_f[0][DATA][1] ) );
  HS65_LS_AOI222X2 U242 ( .A(n66), .B(\chs_in_f[2][DATA][1] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][1] ), .E(n50), .F(
        \chs_in_f[1][DATA][1] ), .Z(n347) );
  HS65_LS_OAI212X5 U243 ( .A(n298), .B(n28), .C(n333), .D(n13), .E(n358), .Z(
        \chs_out_f[0][DATA][2] ) );
  HS65_LS_AOI222X2 U244 ( .A(n67), .B(\chs_in_f[2][DATA][2] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][2] ), .E(n51), .F(
        \chs_in_f[1][DATA][2] ), .Z(n358) );
  HS65_LS_OAI212X5 U245 ( .A(n290), .B(n27), .C(n325), .D(n12), .E(n337), .Z(
        \chs_out_f[0][DATA][10] ) );
  HS65_LS_AOI222X2 U246 ( .A(n66), .B(\chs_in_f[2][DATA][10] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][10] ), .E(n50), .F(
        \chs_in_f[1][DATA][10] ), .Z(n337) );
  HS65_LS_OAI212X5 U247 ( .A(n289), .B(n27), .C(n324), .D(n12), .E(n338), .Z(
        \chs_out_f[0][DATA][11] ) );
  HS65_LS_AOI222X2 U248 ( .A(n66), .B(\chs_in_f[2][DATA][11] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][11] ), .E(n50), .F(
        \chs_in_f[1][DATA][11] ), .Z(n338) );
  HS65_LS_OAI212X5 U249 ( .A(n288), .B(n27), .C(n323), .D(n12), .E(n339), .Z(
        \chs_out_f[0][DATA][12] ) );
  HS65_LS_AOI222X2 U250 ( .A(n66), .B(\chs_in_f[2][DATA][12] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][12] ), .E(n50), .F(
        \chs_in_f[1][DATA][12] ), .Z(n339) );
  HS65_LS_OAI212X5 U251 ( .A(n287), .B(n27), .C(n322), .D(n12), .E(n340), .Z(
        \chs_out_f[0][DATA][13] ) );
  HS65_LS_AOI222X2 U252 ( .A(n66), .B(\chs_in_f[2][DATA][13] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][13] ), .E(n50), .F(
        \chs_in_f[1][DATA][13] ), .Z(n340) );
  HS65_LS_OAI212X5 U253 ( .A(n286), .B(n27), .C(n321), .D(n12), .E(n341), .Z(
        \chs_out_f[0][DATA][14] ) );
  HS65_LS_AOI222X2 U254 ( .A(n66), .B(\chs_in_f[2][DATA][14] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][14] ), .E(n50), .F(
        \chs_in_f[1][DATA][14] ), .Z(n341) );
  HS65_LS_OAI212X5 U255 ( .A(n285), .B(n27), .C(n320), .D(n12), .E(n342), .Z(
        \chs_out_f[0][DATA][15] ) );
  HS65_LS_AOI222X2 U256 ( .A(n66), .B(\chs_in_f[2][DATA][15] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][15] ), .E(n50), .F(
        \chs_in_f[1][DATA][15] ), .Z(n342) );
  HS65_LS_OAI212X5 U257 ( .A(n284), .B(n27), .C(n319), .D(n12), .E(n343), .Z(
        \chs_out_f[0][DATA][16] ) );
  HS65_LS_AOI222X2 U258 ( .A(n66), .B(\chs_in_f[2][DATA][16] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][16] ), .E(n50), .F(
        \chs_in_f[1][DATA][16] ), .Z(n343) );
  HS65_LS_OAI212X5 U259 ( .A(n283), .B(n27), .C(n318), .D(n12), .E(n344), .Z(
        \chs_out_f[0][DATA][17] ) );
  HS65_LS_AOI222X2 U260 ( .A(n66), .B(\chs_in_f[2][DATA][17] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][17] ), .E(n50), .F(
        \chs_in_f[1][DATA][17] ), .Z(n344) );
  HS65_LS_OAI212X5 U261 ( .A(n282), .B(n27), .C(n317), .D(n12), .E(n345), .Z(
        \chs_out_f[0][DATA][18] ) );
  HS65_LS_AOI222X2 U262 ( .A(n66), .B(\chs_in_f[2][DATA][18] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][18] ), .E(n50), .F(
        \chs_in_f[1][DATA][18] ), .Z(n345) );
  HS65_LS_OAI212X5 U263 ( .A(n281), .B(n27), .C(n316), .D(n12), .E(n346), .Z(
        \chs_out_f[0][DATA][19] ) );
  HS65_LS_AOI222X2 U264 ( .A(n66), .B(\chs_in_f[2][DATA][19] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][19] ), .E(n50), .F(
        \chs_in_f[1][DATA][19] ), .Z(n346) );
  HS65_LS_OAI212X5 U265 ( .A(n280), .B(n27), .C(n315), .D(n13), .E(n348), .Z(
        \chs_out_f[0][DATA][20] ) );
  HS65_LS_AOI222X2 U266 ( .A(n67), .B(\chs_in_f[2][DATA][20] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][20] ), .E(n51), .F(
        \chs_in_f[1][DATA][20] ), .Z(n348) );
  HS65_LS_OAI212X5 U267 ( .A(n279), .B(n28), .C(n314), .D(n13), .E(n349), .Z(
        \chs_out_f[0][DATA][21] ) );
  HS65_LS_AOI222X2 U268 ( .A(n67), .B(\chs_in_f[2][DATA][21] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][21] ), .E(n51), .F(
        \chs_in_f[1][DATA][21] ), .Z(n349) );
  HS65_LS_OAI212X5 U269 ( .A(n278), .B(n28), .C(n313), .D(n13), .E(n350), .Z(
        \chs_out_f[0][DATA][22] ) );
  HS65_LS_AOI222X2 U270 ( .A(n67), .B(\chs_in_f[2][DATA][22] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][22] ), .E(n51), .F(
        \chs_in_f[1][DATA][22] ), .Z(n350) );
  HS65_LS_OAI212X5 U271 ( .A(n277), .B(n28), .C(n312), .D(n13), .E(n351), .Z(
        \chs_out_f[0][DATA][23] ) );
  HS65_LS_AOI222X2 U272 ( .A(n67), .B(\chs_in_f[2][DATA][23] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][23] ), .E(n51), .F(
        \chs_in_f[1][DATA][23] ), .Z(n351) );
  HS65_LS_OAI212X5 U273 ( .A(n276), .B(n28), .C(n311), .D(n13), .E(n352), .Z(
        \chs_out_f[0][DATA][24] ) );
  HS65_LS_AOI222X2 U274 ( .A(n67), .B(\chs_in_f[2][DATA][24] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][24] ), .E(n51), .F(
        \chs_in_f[1][DATA][24] ), .Z(n352) );
  HS65_LS_OAI212X5 U275 ( .A(n275), .B(n28), .C(n310), .D(n13), .E(n353), .Z(
        \chs_out_f[0][DATA][25] ) );
  HS65_LS_AOI222X2 U276 ( .A(n67), .B(\chs_in_f[2][DATA][25] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][25] ), .E(n51), .F(
        \chs_in_f[1][DATA][25] ), .Z(n353) );
  HS65_LS_OAI212X5 U277 ( .A(n274), .B(n28), .C(n309), .D(n13), .E(n354), .Z(
        \chs_out_f[0][DATA][26] ) );
  HS65_LS_AOI222X2 U278 ( .A(n67), .B(\chs_in_f[2][DATA][26] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][26] ), .E(n51), .F(
        \chs_in_f[1][DATA][26] ), .Z(n354) );
  HS65_LS_OAI212X5 U279 ( .A(n273), .B(n28), .C(n308), .D(n13), .E(n355), .Z(
        \chs_out_f[0][DATA][27] ) );
  HS65_LS_AOI222X2 U280 ( .A(n67), .B(\chs_in_f[2][DATA][27] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][27] ), .E(n51), .F(
        \chs_in_f[1][DATA][27] ), .Z(n355) );
  HS65_LS_OAI212X5 U281 ( .A(n272), .B(n28), .C(n307), .D(n13), .E(n356), .Z(
        \chs_out_f[0][DATA][28] ) );
  HS65_LS_AOI222X2 U282 ( .A(n67), .B(\chs_in_f[2][DATA][28] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][28] ), .E(n51), .F(
        \chs_in_f[1][DATA][28] ), .Z(n356) );
  HS65_LS_OAI212X5 U283 ( .A(n271), .B(n28), .C(n306), .D(n13), .E(n357), .Z(
        \chs_out_f[0][DATA][29] ) );
  HS65_LS_AOI222X2 U284 ( .A(n67), .B(\chs_in_f[2][DATA][29] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][29] ), .E(n51), .F(
        \chs_in_f[1][DATA][29] ), .Z(n357) );
  HS65_LS_OAI212X5 U285 ( .A(n270), .B(n28), .C(n305), .D(n13), .E(n359), .Z(
        \chs_out_f[0][DATA][30] ) );
  HS65_LS_AOI222X2 U286 ( .A(n67), .B(\chs_in_f[2][DATA][30] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][30] ), .E(n51), .F(
        \chs_in_f[1][DATA][30] ), .Z(n359) );
  HS65_LS_OAI212X5 U287 ( .A(n269), .B(n28), .C(n304), .D(n14), .E(n360), .Z(
        \chs_out_f[0][DATA][31] ) );
  HS65_LS_AOI222X2 U288 ( .A(n68), .B(\chs_in_f[2][DATA][31] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][31] ), .E(n52), .F(
        \chs_in_f[1][DATA][31] ), .Z(n360) );
  HS65_LS_OAI212X5 U289 ( .A(n268), .B(n28), .C(n303), .D(n14), .E(n361), .Z(
        \chs_out_f[0][DATA][32] ) );
  HS65_LS_AOI222X2 U290 ( .A(n68), .B(\chs_in_f[2][DATA][32] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][32] ), .E(n52), .F(
        \chs_in_f[1][DATA][32] ), .Z(n361) );
  HS65_LS_OAI212X5 U291 ( .A(n300), .B(n21), .C(n335), .D(n6), .E(n406), .Z(
        \chs_out_f[2][DATA][0] ) );
  HS65_LS_AOI222X2 U292 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][0] ), 
        .C(n38), .D(\chs_in_f[0][DATA][0] ), .E(n54), .F(
        \chs_in_f[1][DATA][0] ), .Z(n406) );
  HS65_LS_OAI212X5 U293 ( .A(n299), .B(n21), .C(n334), .D(n6), .E(n417), .Z(
        \chs_out_f[2][DATA][1] ) );
  HS65_LS_AOI222X2 U294 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][1] ), 
        .C(n38), .D(\chs_in_f[0][DATA][1] ), .E(n54), .F(
        \chs_in_f[1][DATA][1] ), .Z(n417) );
  HS65_LS_OAI212X5 U295 ( .A(n298), .B(n22), .C(n333), .D(n7), .E(n428), .Z(
        \chs_out_f[2][DATA][2] ) );
  HS65_LS_AOI222X2 U296 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][2] ), 
        .C(n39), .D(\chs_in_f[0][DATA][2] ), .E(n55), .F(
        \chs_in_f[1][DATA][2] ), .Z(n428) );
  HS65_LS_OAI212X5 U297 ( .A(n290), .B(n21), .C(n325), .D(n6), .E(n407), .Z(
        \chs_out_f[2][DATA][10] ) );
  HS65_LS_AOI222X2 U298 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][10] ), 
        .C(n38), .D(\chs_in_f[0][DATA][10] ), .E(n54), .F(
        \chs_in_f[1][DATA][10] ), .Z(n407) );
  HS65_LS_OAI212X5 U299 ( .A(n289), .B(n21), .C(n324), .D(n6), .E(n408), .Z(
        \chs_out_f[2][DATA][11] ) );
  HS65_LS_AOI222X2 U300 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][11] ), 
        .C(n38), .D(\chs_in_f[0][DATA][11] ), .E(n54), .F(
        \chs_in_f[1][DATA][11] ), .Z(n408) );
  HS65_LS_OAI212X5 U301 ( .A(n288), .B(n21), .C(n323), .D(n6), .E(n409), .Z(
        \chs_out_f[2][DATA][12] ) );
  HS65_LS_AOI222X2 U302 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][12] ), 
        .C(n38), .D(\chs_in_f[0][DATA][12] ), .E(n54), .F(
        \chs_in_f[1][DATA][12] ), .Z(n409) );
  HS65_LS_OAI212X5 U303 ( .A(n287), .B(n21), .C(n322), .D(n6), .E(n410), .Z(
        \chs_out_f[2][DATA][13] ) );
  HS65_LS_AOI222X2 U304 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][13] ), 
        .C(n38), .D(\chs_in_f[0][DATA][13] ), .E(n54), .F(
        \chs_in_f[1][DATA][13] ), .Z(n410) );
  HS65_LS_OAI212X5 U305 ( .A(n286), .B(n21), .C(n321), .D(n6), .E(n411), .Z(
        \chs_out_f[2][DATA][14] ) );
  HS65_LS_AOI222X2 U306 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][14] ), 
        .C(n38), .D(\chs_in_f[0][DATA][14] ), .E(n54), .F(
        \chs_in_f[1][DATA][14] ), .Z(n411) );
  HS65_LS_OAI212X5 U307 ( .A(n285), .B(n21), .C(n320), .D(n6), .E(n412), .Z(
        \chs_out_f[2][DATA][15] ) );
  HS65_LS_AOI222X2 U308 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][15] ), 
        .C(n38), .D(\chs_in_f[0][DATA][15] ), .E(n54), .F(
        \chs_in_f[1][DATA][15] ), .Z(n412) );
  HS65_LS_OAI212X5 U309 ( .A(n284), .B(n21), .C(n319), .D(n6), .E(n413), .Z(
        \chs_out_f[2][DATA][16] ) );
  HS65_LS_AOI222X2 U310 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][16] ), 
        .C(n38), .D(\chs_in_f[0][DATA][16] ), .E(n54), .F(
        \chs_in_f[1][DATA][16] ), .Z(n413) );
  HS65_LS_OAI212X5 U311 ( .A(n283), .B(n21), .C(n318), .D(n6), .E(n414), .Z(
        \chs_out_f[2][DATA][17] ) );
  HS65_LS_AOI222X2 U312 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][17] ), 
        .C(n38), .D(\chs_in_f[0][DATA][17] ), .E(n54), .F(
        \chs_in_f[1][DATA][17] ), .Z(n414) );
  HS65_LS_OAI212X5 U313 ( .A(n282), .B(n21), .C(n317), .D(n6), .E(n415), .Z(
        \chs_out_f[2][DATA][18] ) );
  HS65_LS_AOI222X2 U314 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][18] ), 
        .C(n38), .D(\chs_in_f[0][DATA][18] ), .E(n54), .F(
        \chs_in_f[1][DATA][18] ), .Z(n415) );
  HS65_LS_OAI212X5 U315 ( .A(n281), .B(n21), .C(n316), .D(n6), .E(n416), .Z(
        \chs_out_f[2][DATA][19] ) );
  HS65_LS_AOI222X2 U316 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][19] ), 
        .C(n38), .D(\chs_in_f[0][DATA][19] ), .E(n54), .F(
        \chs_in_f[1][DATA][19] ), .Z(n416) );
  HS65_LS_OAI212X5 U317 ( .A(n280), .B(n21), .C(n315), .D(n7), .E(n418), .Z(
        \chs_out_f[2][DATA][20] ) );
  HS65_LS_AOI222X2 U318 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][20] ), 
        .C(n39), .D(\chs_in_f[0][DATA][20] ), .E(n55), .F(
        \chs_in_f[1][DATA][20] ), .Z(n418) );
  HS65_LS_OAI212X5 U319 ( .A(n279), .B(n22), .C(n314), .D(n7), .E(n419), .Z(
        \chs_out_f[2][DATA][21] ) );
  HS65_LS_AOI222X2 U320 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][21] ), 
        .C(n39), .D(\chs_in_f[0][DATA][21] ), .E(n55), .F(
        \chs_in_f[1][DATA][21] ), .Z(n419) );
  HS65_LS_OAI212X5 U321 ( .A(n278), .B(n22), .C(n313), .D(n7), .E(n420), .Z(
        \chs_out_f[2][DATA][22] ) );
  HS65_LS_AOI222X2 U322 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][22] ), 
        .C(n39), .D(\chs_in_f[0][DATA][22] ), .E(n55), .F(
        \chs_in_f[1][DATA][22] ), .Z(n420) );
  HS65_LS_OAI212X5 U323 ( .A(n277), .B(n22), .C(n312), .D(n7), .E(n421), .Z(
        \chs_out_f[2][DATA][23] ) );
  HS65_LS_AOI222X2 U324 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][23] ), 
        .C(n39), .D(\chs_in_f[0][DATA][23] ), .E(n55), .F(
        \chs_in_f[1][DATA][23] ), .Z(n421) );
  HS65_LS_OAI212X5 U325 ( .A(n276), .B(n22), .C(n311), .D(n7), .E(n422), .Z(
        \chs_out_f[2][DATA][24] ) );
  HS65_LS_AOI222X2 U326 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][24] ), 
        .C(n39), .D(\chs_in_f[0][DATA][24] ), .E(n55), .F(
        \chs_in_f[1][DATA][24] ), .Z(n422) );
  HS65_LS_OAI212X5 U327 ( .A(n275), .B(n22), .C(n310), .D(n7), .E(n423), .Z(
        \chs_out_f[2][DATA][25] ) );
  HS65_LS_AOI222X2 U328 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][25] ), 
        .C(n39), .D(\chs_in_f[0][DATA][25] ), .E(n55), .F(
        \chs_in_f[1][DATA][25] ), .Z(n423) );
  HS65_LS_OAI212X5 U329 ( .A(n274), .B(n22), .C(n309), .D(n7), .E(n424), .Z(
        \chs_out_f[2][DATA][26] ) );
  HS65_LS_AOI222X2 U330 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][26] ), 
        .C(n39), .D(\chs_in_f[0][DATA][26] ), .E(n55), .F(
        \chs_in_f[1][DATA][26] ), .Z(n424) );
  HS65_LS_OAI212X5 U331 ( .A(n273), .B(n22), .C(n308), .D(n7), .E(n425), .Z(
        \chs_out_f[2][DATA][27] ) );
  HS65_LS_AOI222X2 U332 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][27] ), 
        .C(n39), .D(\chs_in_f[0][DATA][27] ), .E(n55), .F(
        \chs_in_f[1][DATA][27] ), .Z(n425) );
  HS65_LS_OAI212X5 U333 ( .A(n272), .B(n22), .C(n307), .D(n7), .E(n426), .Z(
        \chs_out_f[2][DATA][28] ) );
  HS65_LS_AOI222X2 U334 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][28] ), 
        .C(n39), .D(\chs_in_f[0][DATA][28] ), .E(n55), .F(
        \chs_in_f[1][DATA][28] ), .Z(n426) );
  HS65_LS_OAI212X5 U335 ( .A(n271), .B(n22), .C(n306), .D(n7), .E(n427), .Z(
        \chs_out_f[2][DATA][29] ) );
  HS65_LS_AOI222X2 U336 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][29] ), 
        .C(n39), .D(\chs_in_f[0][DATA][29] ), .E(n55), .F(
        \chs_in_f[1][DATA][29] ), .Z(n427) );
  HS65_LS_OAI212X5 U337 ( .A(n270), .B(n22), .C(n305), .D(n7), .E(n429), .Z(
        \chs_out_f[2][DATA][30] ) );
  HS65_LS_AOI222X2 U338 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][30] ), 
        .C(n39), .D(\chs_in_f[0][DATA][30] ), .E(n55), .F(
        \chs_in_f[1][DATA][30] ), .Z(n429) );
  HS65_LS_OAI212X5 U339 ( .A(n269), .B(n22), .C(n304), .D(n8), .E(n430), .Z(
        \chs_out_f[2][DATA][31] ) );
  HS65_LS_AOI222X2 U340 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][31] ), 
        .C(n40), .D(\chs_in_f[0][DATA][31] ), .E(n56), .F(
        \chs_in_f[1][DATA][31] ), .Z(n430) );
  HS65_LS_OAI212X5 U341 ( .A(n268), .B(n22), .C(n303), .D(n8), .E(n431), .Z(
        \chs_out_f[2][DATA][32] ) );
  HS65_LS_AOI222X2 U342 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][32] ), 
        .C(n40), .D(\chs_in_f[0][DATA][32] ), .E(n56), .F(
        \chs_in_f[1][DATA][32] ), .Z(n431) );
  HS65_LS_OAI212X5 U343 ( .A(n300), .B(n24), .C(n335), .D(n9), .E(n371), .Z(
        \chs_out_f[1][DATA][0] ) );
  HS65_LS_AOI222X2 U344 ( .A(n70), .B(\chs_in_f[2][DATA][0] ), .C(n34), .D(
        \chs_in_f[0][DATA][0] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][0] ), .Z(n371) );
  HS65_LS_OAI212X5 U345 ( .A(n299), .B(n24), .C(n334), .D(n9), .E(n382), .Z(
        \chs_out_f[1][DATA][1] ) );
  HS65_LS_AOI222X2 U346 ( .A(n70), .B(\chs_in_f[2][DATA][1] ), .C(n34), .D(
        \chs_in_f[0][DATA][1] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][1] ), .Z(n382) );
  HS65_LS_OAI212X5 U347 ( .A(n298), .B(n25), .C(n333), .D(n10), .E(n393), .Z(
        \chs_out_f[1][DATA][2] ) );
  HS65_LS_AOI222X2 U348 ( .A(n71), .B(\chs_in_f[2][DATA][2] ), .C(n35), .D(
        \chs_in_f[0][DATA][2] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][2] ), .Z(n393) );
  HS65_LS_OAI212X5 U349 ( .A(n290), .B(n24), .C(n325), .D(n9), .E(n372), .Z(
        \chs_out_f[1][DATA][10] ) );
  HS65_LS_AOI222X2 U350 ( .A(n70), .B(\chs_in_f[2][DATA][10] ), .C(n34), .D(
        \chs_in_f[0][DATA][10] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][10] ), .Z(n372) );
  HS65_LS_OAI212X5 U351 ( .A(n289), .B(n24), .C(n324), .D(n9), .E(n373), .Z(
        \chs_out_f[1][DATA][11] ) );
  HS65_LS_AOI222X2 U352 ( .A(n70), .B(\chs_in_f[2][DATA][11] ), .C(n34), .D(
        \chs_in_f[0][DATA][11] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][11] ), .Z(n373) );
  HS65_LS_OAI212X5 U353 ( .A(n288), .B(n24), .C(n323), .D(n9), .E(n374), .Z(
        \chs_out_f[1][DATA][12] ) );
  HS65_LS_AOI222X2 U354 ( .A(n70), .B(\chs_in_f[2][DATA][12] ), .C(n34), .D(
        \chs_in_f[0][DATA][12] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][12] ), .Z(n374) );
  HS65_LS_OAI212X5 U355 ( .A(n287), .B(n24), .C(n322), .D(n9), .E(n375), .Z(
        \chs_out_f[1][DATA][13] ) );
  HS65_LS_AOI222X2 U356 ( .A(n70), .B(\chs_in_f[2][DATA][13] ), .C(n34), .D(
        \chs_in_f[0][DATA][13] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][13] ), .Z(n375) );
  HS65_LS_OAI212X5 U357 ( .A(n286), .B(n24), .C(n321), .D(n9), .E(n376), .Z(
        \chs_out_f[1][DATA][14] ) );
  HS65_LS_AOI222X2 U358 ( .A(n70), .B(\chs_in_f[2][DATA][14] ), .C(n34), .D(
        \chs_in_f[0][DATA][14] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][14] ), .Z(n376) );
  HS65_LS_OAI212X5 U359 ( .A(n285), .B(n24), .C(n320), .D(n9), .E(n377), .Z(
        \chs_out_f[1][DATA][15] ) );
  HS65_LS_AOI222X2 U360 ( .A(n70), .B(\chs_in_f[2][DATA][15] ), .C(n34), .D(
        \chs_in_f[0][DATA][15] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][15] ), .Z(n377) );
  HS65_LS_OAI212X5 U361 ( .A(n284), .B(n24), .C(n319), .D(n9), .E(n378), .Z(
        \chs_out_f[1][DATA][16] ) );
  HS65_LS_AOI222X2 U362 ( .A(n70), .B(\chs_in_f[2][DATA][16] ), .C(n34), .D(
        \chs_in_f[0][DATA][16] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][16] ), .Z(n378) );
  HS65_LS_OAI212X5 U363 ( .A(n283), .B(n24), .C(n318), .D(n9), .E(n379), .Z(
        \chs_out_f[1][DATA][17] ) );
  HS65_LS_AOI222X2 U364 ( .A(n70), .B(\chs_in_f[2][DATA][17] ), .C(n34), .D(
        \chs_in_f[0][DATA][17] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][17] ), .Z(n379) );
  HS65_LS_OAI212X5 U365 ( .A(n282), .B(n24), .C(n317), .D(n9), .E(n380), .Z(
        \chs_out_f[1][DATA][18] ) );
  HS65_LS_AOI222X2 U366 ( .A(n70), .B(\chs_in_f[2][DATA][18] ), .C(n34), .D(
        \chs_in_f[0][DATA][18] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][18] ), .Z(n380) );
  HS65_LS_OAI212X5 U367 ( .A(n281), .B(n24), .C(n316), .D(n9), .E(n381), .Z(
        \chs_out_f[1][DATA][19] ) );
  HS65_LS_AOI222X2 U368 ( .A(n70), .B(\chs_in_f[2][DATA][19] ), .C(n34), .D(
        \chs_in_f[0][DATA][19] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][19] ), .Z(n381) );
  HS65_LS_OAI212X5 U369 ( .A(n280), .B(n24), .C(n315), .D(n10), .E(n383), .Z(
        \chs_out_f[1][DATA][20] ) );
  HS65_LS_AOI222X2 U370 ( .A(n71), .B(\chs_in_f[2][DATA][20] ), .C(n35), .D(
        \chs_in_f[0][DATA][20] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][20] ), .Z(n383) );
  HS65_LS_OAI212X5 U371 ( .A(n279), .B(n25), .C(n314), .D(n10), .E(n384), .Z(
        \chs_out_f[1][DATA][21] ) );
  HS65_LS_AOI222X2 U372 ( .A(n71), .B(\chs_in_f[2][DATA][21] ), .C(n35), .D(
        \chs_in_f[0][DATA][21] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][21] ), .Z(n384) );
  HS65_LS_OAI212X5 U373 ( .A(n278), .B(n25), .C(n313), .D(n10), .E(n385), .Z(
        \chs_out_f[1][DATA][22] ) );
  HS65_LS_AOI222X2 U374 ( .A(n71), .B(\chs_in_f[2][DATA][22] ), .C(n35), .D(
        \chs_in_f[0][DATA][22] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][22] ), .Z(n385) );
  HS65_LS_OAI212X5 U375 ( .A(n277), .B(n25), .C(n312), .D(n10), .E(n386), .Z(
        \chs_out_f[1][DATA][23] ) );
  HS65_LS_AOI222X2 U376 ( .A(n71), .B(\chs_in_f[2][DATA][23] ), .C(n35), .D(
        \chs_in_f[0][DATA][23] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][23] ), .Z(n386) );
  HS65_LS_OAI212X5 U377 ( .A(n276), .B(n25), .C(n311), .D(n10), .E(n387), .Z(
        \chs_out_f[1][DATA][24] ) );
  HS65_LS_AOI222X2 U378 ( .A(n71), .B(\chs_in_f[2][DATA][24] ), .C(n35), .D(
        \chs_in_f[0][DATA][24] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][24] ), .Z(n387) );
  HS65_LS_OAI212X5 U379 ( .A(n275), .B(n25), .C(n310), .D(n10), .E(n388), .Z(
        \chs_out_f[1][DATA][25] ) );
  HS65_LS_AOI222X2 U380 ( .A(n71), .B(\chs_in_f[2][DATA][25] ), .C(n35), .D(
        \chs_in_f[0][DATA][25] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][25] ), .Z(n388) );
  HS65_LS_OAI212X5 U381 ( .A(n274), .B(n25), .C(n309), .D(n10), .E(n389), .Z(
        \chs_out_f[1][DATA][26] ) );
  HS65_LS_AOI222X2 U382 ( .A(n71), .B(\chs_in_f[2][DATA][26] ), .C(n35), .D(
        \chs_in_f[0][DATA][26] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][26] ), .Z(n389) );
  HS65_LS_OAI212X5 U383 ( .A(n273), .B(n25), .C(n308), .D(n10), .E(n390), .Z(
        \chs_out_f[1][DATA][27] ) );
  HS65_LS_AOI222X2 U384 ( .A(n71), .B(\chs_in_f[2][DATA][27] ), .C(n35), .D(
        \chs_in_f[0][DATA][27] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][27] ), .Z(n390) );
  HS65_LS_OAI212X5 U385 ( .A(n272), .B(n25), .C(n307), .D(n10), .E(n391), .Z(
        \chs_out_f[1][DATA][28] ) );
  HS65_LS_AOI222X2 U386 ( .A(n71), .B(\chs_in_f[2][DATA][28] ), .C(n35), .D(
        \chs_in_f[0][DATA][28] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][28] ), .Z(n391) );
  HS65_LS_OAI212X5 U387 ( .A(n271), .B(n25), .C(n306), .D(n10), .E(n392), .Z(
        \chs_out_f[1][DATA][29] ) );
  HS65_LS_AOI222X2 U388 ( .A(n71), .B(\chs_in_f[2][DATA][29] ), .C(n35), .D(
        \chs_in_f[0][DATA][29] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][29] ), .Z(n392) );
  HS65_LS_OAI212X5 U389 ( .A(n270), .B(n25), .C(n305), .D(n10), .E(n394), .Z(
        \chs_out_f[1][DATA][30] ) );
  HS65_LS_AOI222X2 U390 ( .A(n71), .B(\chs_in_f[2][DATA][30] ), .C(n35), .D(
        \chs_in_f[0][DATA][30] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][30] ), .Z(n394) );
  HS65_LS_OAI212X5 U391 ( .A(n269), .B(n25), .C(n304), .D(n11), .E(n395), .Z(
        \chs_out_f[1][DATA][31] ) );
  HS65_LS_AOI222X2 U392 ( .A(n72), .B(\chs_in_f[2][DATA][31] ), .C(n36), .D(
        \chs_in_f[0][DATA][31] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][31] ), .Z(n395) );
  HS65_LS_OAI212X5 U393 ( .A(n268), .B(n25), .C(n303), .D(n11), .E(n396), .Z(
        \chs_out_f[1][DATA][32] ) );
  HS65_LS_AOI222X2 U394 ( .A(n72), .B(\chs_in_f[2][DATA][32] ), .C(n36), .D(
        \chs_in_f[0][DATA][32] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][32] ), .Z(n396) );
  HS65_LS_OAI212X5 U395 ( .A(n297), .B(n29), .C(n332), .D(n14), .E(n364), .Z(
        \chs_out_f[0][DATA][3] ) );
  HS65_LS_AOI222X2 U396 ( .A(n68), .B(\chs_in_f[2][DATA][3] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][3] ), .E(n52), .F(
        \chs_in_f[1][DATA][3] ), .Z(n364) );
  HS65_LS_OAI212X5 U397 ( .A(n296), .B(n29), .C(n331), .D(n14), .E(n365), .Z(
        \chs_out_f[0][DATA][4] ) );
  HS65_LS_AOI222X2 U398 ( .A(n68), .B(\chs_in_f[2][DATA][4] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][4] ), .E(n52), .F(
        \chs_in_f[1][DATA][4] ), .Z(n365) );
  HS65_LS_OAI212X5 U399 ( .A(n295), .B(n29), .C(n330), .D(n14), .E(n366), .Z(
        \chs_out_f[0][DATA][5] ) );
  HS65_LS_AOI222X2 U400 ( .A(n68), .B(\chs_in_f[2][DATA][5] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][5] ), .E(n52), .F(
        \chs_in_f[1][DATA][5] ), .Z(n366) );
  HS65_LS_OAI212X5 U401 ( .A(n294), .B(n29), .C(n329), .D(n14), .E(n367), .Z(
        \chs_out_f[0][DATA][6] ) );
  HS65_LS_AOI222X2 U402 ( .A(n68), .B(\chs_in_f[2][DATA][6] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][6] ), .E(n52), .F(
        \chs_in_f[1][DATA][6] ), .Z(n367) );
  HS65_LS_OAI212X5 U403 ( .A(n293), .B(n29), .C(n328), .D(n14), .E(n368), .Z(
        \chs_out_f[0][DATA][7] ) );
  HS65_LS_AOI222X2 U404 ( .A(n68), .B(\chs_in_f[2][DATA][7] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][7] ), .E(n52), .F(
        \chs_in_f[1][DATA][7] ), .Z(n368) );
  HS65_LS_OAI212X5 U405 ( .A(n292), .B(n29), .C(n327), .D(n14), .E(n369), .Z(
        \chs_out_f[0][DATA][8] ) );
  HS65_LS_AOI222X2 U406 ( .A(n68), .B(\chs_in_f[2][DATA][8] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][8] ), .E(n52), .F(
        \chs_in_f[1][DATA][8] ), .Z(n369) );
  HS65_LS_OAI212X5 U407 ( .A(n267), .B(n29), .C(n302), .D(n14), .E(n362), .Z(
        \chs_out_f[0][DATA][33] ) );
  HS65_LS_AOI222X2 U408 ( .A(n68), .B(\chs_in_f[2][DATA][33] ), .C(
        \switch_sel[0][0] ), .D(\chs_in_f[0][DATA][33] ), .E(n52), .F(
        \chs_in_f[1][DATA][33] ), .Z(n362) );
  HS65_LS_OAI212X5 U409 ( .A(n297), .B(n23), .C(n332), .D(n8), .E(n434), .Z(
        \chs_out_f[2][DATA][3] ) );
  HS65_LS_AOI222X2 U410 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][3] ), 
        .C(n40), .D(\chs_in_f[0][DATA][3] ), .E(n56), .F(
        \chs_in_f[1][DATA][3] ), .Z(n434) );
  HS65_LS_OAI212X5 U411 ( .A(n296), .B(n23), .C(n331), .D(n8), .E(n435), .Z(
        \chs_out_f[2][DATA][4] ) );
  HS65_LS_AOI222X2 U412 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][4] ), 
        .C(n40), .D(\chs_in_f[0][DATA][4] ), .E(n56), .F(
        \chs_in_f[1][DATA][4] ), .Z(n435) );
  HS65_LS_OAI212X5 U413 ( .A(n295), .B(n23), .C(n330), .D(n8), .E(n436), .Z(
        \chs_out_f[2][DATA][5] ) );
  HS65_LS_AOI222X2 U414 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][5] ), 
        .C(n40), .D(\chs_in_f[0][DATA][5] ), .E(n56), .F(
        \chs_in_f[1][DATA][5] ), .Z(n436) );
  HS65_LS_OAI212X5 U415 ( .A(n294), .B(n23), .C(n329), .D(n8), .E(n437), .Z(
        \chs_out_f[2][DATA][6] ) );
  HS65_LS_AOI222X2 U416 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][6] ), 
        .C(n40), .D(\chs_in_f[0][DATA][6] ), .E(n56), .F(
        \chs_in_f[1][DATA][6] ), .Z(n437) );
  HS65_LS_OAI212X5 U417 ( .A(n293), .B(n23), .C(n328), .D(n8), .E(n438), .Z(
        \chs_out_f[2][DATA][7] ) );
  HS65_LS_AOI222X2 U418 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][7] ), 
        .C(n40), .D(\chs_in_f[0][DATA][7] ), .E(n56), .F(
        \chs_in_f[1][DATA][7] ), .Z(n438) );
  HS65_LS_OAI212X5 U419 ( .A(n292), .B(n23), .C(n327), .D(n8), .E(n439), .Z(
        \chs_out_f[2][DATA][8] ) );
  HS65_LS_AOI222X2 U420 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][8] ), 
        .C(n40), .D(\chs_in_f[0][DATA][8] ), .E(n56), .F(
        \chs_in_f[1][DATA][8] ), .Z(n439) );
  HS65_LS_OAI212X5 U421 ( .A(n267), .B(n23), .C(n302), .D(n8), .E(n432), .Z(
        \chs_out_f[2][DATA][33] ) );
  HS65_LS_AOI222X2 U422 ( .A(\switch_sel[2][2] ), .B(\chs_in_f[2][DATA][33] ), 
        .C(n40), .D(\chs_in_f[0][DATA][33] ), .E(n56), .F(
        \chs_in_f[1][DATA][33] ), .Z(n432) );
  HS65_LS_OAI212X5 U423 ( .A(n297), .B(n26), .C(n332), .D(n11), .E(n399), .Z(
        \chs_out_f[1][DATA][3] ) );
  HS65_LS_AOI222X2 U424 ( .A(n72), .B(\chs_in_f[2][DATA][3] ), .C(n36), .D(
        \chs_in_f[0][DATA][3] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][3] ), .Z(n399) );
  HS65_LS_OAI212X5 U425 ( .A(n296), .B(n26), .C(n331), .D(n11), .E(n400), .Z(
        \chs_out_f[1][DATA][4] ) );
  HS65_LS_AOI222X2 U426 ( .A(n72), .B(\chs_in_f[2][DATA][4] ), .C(n36), .D(
        \chs_in_f[0][DATA][4] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][4] ), .Z(n400) );
  HS65_LS_OAI212X5 U427 ( .A(n295), .B(n26), .C(n330), .D(n11), .E(n401), .Z(
        \chs_out_f[1][DATA][5] ) );
  HS65_LS_AOI222X2 U428 ( .A(n72), .B(\chs_in_f[2][DATA][5] ), .C(n36), .D(
        \chs_in_f[0][DATA][5] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][5] ), .Z(n401) );
  HS65_LS_OAI212X5 U429 ( .A(n294), .B(n26), .C(n329), .D(n11), .E(n402), .Z(
        \chs_out_f[1][DATA][6] ) );
  HS65_LS_AOI222X2 U430 ( .A(n72), .B(\chs_in_f[2][DATA][6] ), .C(n36), .D(
        \chs_in_f[0][DATA][6] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][6] ), .Z(n402) );
  HS65_LS_OAI212X5 U431 ( .A(n293), .B(n26), .C(n328), .D(n11), .E(n403), .Z(
        \chs_out_f[1][DATA][7] ) );
  HS65_LS_AOI222X2 U432 ( .A(n72), .B(\chs_in_f[2][DATA][7] ), .C(n36), .D(
        \chs_in_f[0][DATA][7] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][7] ), .Z(n403) );
  HS65_LS_OAI212X5 U433 ( .A(n292), .B(n26), .C(n327), .D(n11), .E(n404), .Z(
        \chs_out_f[1][DATA][8] ) );
  HS65_LS_AOI222X2 U434 ( .A(n72), .B(\chs_in_f[2][DATA][8] ), .C(n36), .D(
        \chs_in_f[0][DATA][8] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][8] ), .Z(n404) );
  HS65_LS_OAI212X5 U435 ( .A(n267), .B(n26), .C(n302), .D(n11), .E(n397), .Z(
        \chs_out_f[1][DATA][33] ) );
  HS65_LS_AOI222X2 U436 ( .A(n72), .B(\chs_in_f[2][DATA][33] ), .C(n36), .D(
        \chs_in_f[0][DATA][33] ), .E(\switch_sel[1][1] ), .F(
        \chs_in_f[1][DATA][33] ), .Z(n397) );
  HS65_LS_OAI212X5 U437 ( .A(n291), .B(n32), .C(n326), .D(n5), .E(n475), .Z(
        \chs_out_f[3][DATA][9] ) );
  HS65_LS_AOI222X2 U438 ( .A(n76), .B(\chs_in_f[2][DATA][9] ), .C(n44), .D(
        \chs_in_f[0][DATA][9] ), .E(n60), .F(\chs_in_f[1][DATA][9] ), .Z(n475)
         );
  HS65_LS_OAI212X5 U439 ( .A(n300), .B(n30), .C(n335), .D(n3), .E(n441), .Z(
        \chs_out_f[3][DATA][0] ) );
  HS65_LS_AOI222X2 U440 ( .A(n74), .B(\chs_in_f[2][DATA][0] ), .C(n42), .D(
        \chs_in_f[0][DATA][0] ), .E(n58), .F(\chs_in_f[1][DATA][0] ), .Z(n441)
         );
  HS65_LS_OAI212X5 U441 ( .A(n299), .B(n30), .C(n334), .D(n3), .E(n452), .Z(
        \chs_out_f[3][DATA][1] ) );
  HS65_LS_AOI222X2 U442 ( .A(n74), .B(\chs_in_f[2][DATA][1] ), .C(n42), .D(
        \chs_in_f[0][DATA][1] ), .E(n58), .F(\chs_in_f[1][DATA][1] ), .Z(n452)
         );
  HS65_LS_OAI212X5 U443 ( .A(n298), .B(n31), .C(n333), .D(n4), .E(n463), .Z(
        \chs_out_f[3][DATA][2] ) );
  HS65_LS_AOI222X2 U444 ( .A(n75), .B(\chs_in_f[2][DATA][2] ), .C(n43), .D(
        \chs_in_f[0][DATA][2] ), .E(n59), .F(\chs_in_f[1][DATA][2] ), .Z(n463)
         );
  HS65_LS_OAI212X5 U445 ( .A(n297), .B(n32), .C(n332), .D(n5), .E(n469), .Z(
        \chs_out_f[3][DATA][3] ) );
  HS65_LS_AOI222X2 U446 ( .A(n76), .B(\chs_in_f[2][DATA][3] ), .C(n44), .D(
        \chs_in_f[0][DATA][3] ), .E(n60), .F(\chs_in_f[1][DATA][3] ), .Z(n469)
         );
  HS65_LS_OAI212X5 U447 ( .A(n296), .B(n32), .C(n331), .D(n5), .E(n470), .Z(
        \chs_out_f[3][DATA][4] ) );
  HS65_LS_AOI222X2 U448 ( .A(n76), .B(\chs_in_f[2][DATA][4] ), .C(n44), .D(
        \chs_in_f[0][DATA][4] ), .E(n60), .F(\chs_in_f[1][DATA][4] ), .Z(n470)
         );
  HS65_LS_OAI212X5 U449 ( .A(n295), .B(n32), .C(n330), .D(n5), .E(n471), .Z(
        \chs_out_f[3][DATA][5] ) );
  HS65_LS_AOI222X2 U450 ( .A(n76), .B(\chs_in_f[2][DATA][5] ), .C(n44), .D(
        \chs_in_f[0][DATA][5] ), .E(n60), .F(\chs_in_f[1][DATA][5] ), .Z(n471)
         );
  HS65_LS_OAI212X5 U451 ( .A(n294), .B(n32), .C(n329), .D(n5), .E(n472), .Z(
        \chs_out_f[3][DATA][6] ) );
  HS65_LS_AOI222X2 U452 ( .A(n76), .B(\chs_in_f[2][DATA][6] ), .C(n44), .D(
        \chs_in_f[0][DATA][6] ), .E(n60), .F(\chs_in_f[1][DATA][6] ), .Z(n472)
         );
  HS65_LS_OAI212X5 U453 ( .A(n293), .B(n32), .C(n328), .D(n5), .E(n473), .Z(
        \chs_out_f[3][DATA][7] ) );
  HS65_LS_AOI222X2 U454 ( .A(n76), .B(\chs_in_f[2][DATA][7] ), .C(n44), .D(
        \chs_in_f[0][DATA][7] ), .E(n60), .F(\chs_in_f[1][DATA][7] ), .Z(n473)
         );
  HS65_LS_OAI212X5 U455 ( .A(n292), .B(n32), .C(n327), .D(n5), .E(n474), .Z(
        \chs_out_f[3][DATA][8] ) );
  HS65_LS_AOI222X2 U456 ( .A(n76), .B(\chs_in_f[2][DATA][8] ), .C(n44), .D(
        \chs_in_f[0][DATA][8] ), .E(n60), .F(\chs_in_f[1][DATA][8] ), .Z(n474)
         );
  HS65_LS_OAI212X5 U457 ( .A(n290), .B(n30), .C(n325), .D(n3), .E(n442), .Z(
        \chs_out_f[3][DATA][10] ) );
  HS65_LS_AOI222X2 U458 ( .A(n74), .B(\chs_in_f[2][DATA][10] ), .C(n42), .D(
        \chs_in_f[0][DATA][10] ), .E(n58), .F(\chs_in_f[1][DATA][10] ), .Z(
        n442) );
  HS65_LS_OAI212X5 U459 ( .A(n289), .B(n30), .C(n324), .D(n3), .E(n443), .Z(
        \chs_out_f[3][DATA][11] ) );
  HS65_LS_AOI222X2 U460 ( .A(n74), .B(\chs_in_f[2][DATA][11] ), .C(n42), .D(
        \chs_in_f[0][DATA][11] ), .E(n58), .F(\chs_in_f[1][DATA][11] ), .Z(
        n443) );
  HS65_LS_OAI212X5 U461 ( .A(n288), .B(n30), .C(n323), .D(n3), .E(n444), .Z(
        \chs_out_f[3][DATA][12] ) );
  HS65_LS_AOI222X2 U462 ( .A(n74), .B(\chs_in_f[2][DATA][12] ), .C(n42), .D(
        \chs_in_f[0][DATA][12] ), .E(n58), .F(\chs_in_f[1][DATA][12] ), .Z(
        n444) );
  HS65_LS_OAI212X5 U463 ( .A(n287), .B(n30), .C(n322), .D(n3), .E(n445), .Z(
        \chs_out_f[3][DATA][13] ) );
  HS65_LS_AOI222X2 U464 ( .A(n74), .B(\chs_in_f[2][DATA][13] ), .C(n42), .D(
        \chs_in_f[0][DATA][13] ), .E(n58), .F(\chs_in_f[1][DATA][13] ), .Z(
        n445) );
  HS65_LS_OAI212X5 U465 ( .A(n286), .B(n30), .C(n321), .D(n3), .E(n446), .Z(
        \chs_out_f[3][DATA][14] ) );
  HS65_LS_AOI222X2 U466 ( .A(n74), .B(\chs_in_f[2][DATA][14] ), .C(n42), .D(
        \chs_in_f[0][DATA][14] ), .E(n58), .F(\chs_in_f[1][DATA][14] ), .Z(
        n446) );
  HS65_LS_OAI212X5 U467 ( .A(n285), .B(n30), .C(n320), .D(n3), .E(n447), .Z(
        \chs_out_f[3][DATA][15] ) );
  HS65_LS_AOI222X2 U468 ( .A(n74), .B(\chs_in_f[2][DATA][15] ), .C(n42), .D(
        \chs_in_f[0][DATA][15] ), .E(n58), .F(\chs_in_f[1][DATA][15] ), .Z(
        n447) );
  HS65_LS_OAI212X5 U469 ( .A(n284), .B(n30), .C(n319), .D(n3), .E(n448), .Z(
        \chs_out_f[3][DATA][16] ) );
  HS65_LS_AOI222X2 U470 ( .A(n74), .B(\chs_in_f[2][DATA][16] ), .C(n42), .D(
        \chs_in_f[0][DATA][16] ), .E(n58), .F(\chs_in_f[1][DATA][16] ), .Z(
        n448) );
  HS65_LS_OAI212X5 U471 ( .A(n283), .B(n30), .C(n318), .D(n3), .E(n449), .Z(
        \chs_out_f[3][DATA][17] ) );
  HS65_LS_AOI222X2 U472 ( .A(n74), .B(\chs_in_f[2][DATA][17] ), .C(n42), .D(
        \chs_in_f[0][DATA][17] ), .E(n58), .F(\chs_in_f[1][DATA][17] ), .Z(
        n449) );
  HS65_LS_OAI212X5 U473 ( .A(n282), .B(n30), .C(n317), .D(n3), .E(n450), .Z(
        \chs_out_f[3][DATA][18] ) );
  HS65_LS_AOI222X2 U474 ( .A(n74), .B(\chs_in_f[2][DATA][18] ), .C(n42), .D(
        \chs_in_f[0][DATA][18] ), .E(n58), .F(\chs_in_f[1][DATA][18] ), .Z(
        n450) );
  HS65_LS_OAI212X5 U475 ( .A(n281), .B(n30), .C(n316), .D(n3), .E(n451), .Z(
        \chs_out_f[3][DATA][19] ) );
  HS65_LS_AOI222X2 U476 ( .A(n74), .B(\chs_in_f[2][DATA][19] ), .C(n42), .D(
        \chs_in_f[0][DATA][19] ), .E(n58), .F(\chs_in_f[1][DATA][19] ), .Z(
        n451) );
  HS65_LS_OAI212X5 U477 ( .A(n280), .B(n30), .C(n315), .D(n4), .E(n453), .Z(
        \chs_out_f[3][DATA][20] ) );
  HS65_LS_AOI222X2 U478 ( .A(n75), .B(\chs_in_f[2][DATA][20] ), .C(n43), .D(
        \chs_in_f[0][DATA][20] ), .E(n59), .F(\chs_in_f[1][DATA][20] ), .Z(
        n453) );
  HS65_LS_OAI212X5 U479 ( .A(n279), .B(n31), .C(n314), .D(n4), .E(n454), .Z(
        \chs_out_f[3][DATA][21] ) );
  HS65_LS_AOI222X2 U480 ( .A(n75), .B(\chs_in_f[2][DATA][21] ), .C(n43), .D(
        \chs_in_f[0][DATA][21] ), .E(n59), .F(\chs_in_f[1][DATA][21] ), .Z(
        n454) );
  HS65_LS_OAI212X5 U481 ( .A(n278), .B(n31), .C(n313), .D(n4), .E(n455), .Z(
        \chs_out_f[3][DATA][22] ) );
  HS65_LS_AOI222X2 U482 ( .A(n75), .B(\chs_in_f[2][DATA][22] ), .C(n43), .D(
        \chs_in_f[0][DATA][22] ), .E(n59), .F(\chs_in_f[1][DATA][22] ), .Z(
        n455) );
  HS65_LS_OAI212X5 U483 ( .A(n277), .B(n31), .C(n312), .D(n4), .E(n456), .Z(
        \chs_out_f[3][DATA][23] ) );
  HS65_LS_AOI222X2 U484 ( .A(n75), .B(\chs_in_f[2][DATA][23] ), .C(n43), .D(
        \chs_in_f[0][DATA][23] ), .E(n59), .F(\chs_in_f[1][DATA][23] ), .Z(
        n456) );
  HS65_LS_OAI212X5 U485 ( .A(n276), .B(n31), .C(n311), .D(n4), .E(n457), .Z(
        \chs_out_f[3][DATA][24] ) );
  HS65_LS_AOI222X2 U486 ( .A(n75), .B(\chs_in_f[2][DATA][24] ), .C(n43), .D(
        \chs_in_f[0][DATA][24] ), .E(n59), .F(\chs_in_f[1][DATA][24] ), .Z(
        n457) );
  HS65_LS_OAI212X5 U487 ( .A(n275), .B(n31), .C(n310), .D(n4), .E(n458), .Z(
        \chs_out_f[3][DATA][25] ) );
  HS65_LS_AOI222X2 U488 ( .A(n75), .B(\chs_in_f[2][DATA][25] ), .C(n43), .D(
        \chs_in_f[0][DATA][25] ), .E(n59), .F(\chs_in_f[1][DATA][25] ), .Z(
        n458) );
  HS65_LS_OAI212X5 U489 ( .A(n274), .B(n31), .C(n309), .D(n4), .E(n459), .Z(
        \chs_out_f[3][DATA][26] ) );
  HS65_LS_AOI222X2 U490 ( .A(n75), .B(\chs_in_f[2][DATA][26] ), .C(n43), .D(
        \chs_in_f[0][DATA][26] ), .E(n59), .F(\chs_in_f[1][DATA][26] ), .Z(
        n459) );
  HS65_LS_OAI212X5 U491 ( .A(n273), .B(n31), .C(n308), .D(n4), .E(n460), .Z(
        \chs_out_f[3][DATA][27] ) );
  HS65_LS_AOI222X2 U492 ( .A(n75), .B(\chs_in_f[2][DATA][27] ), .C(n43), .D(
        \chs_in_f[0][DATA][27] ), .E(n59), .F(\chs_in_f[1][DATA][27] ), .Z(
        n460) );
  HS65_LS_OAI212X5 U493 ( .A(n272), .B(n31), .C(n307), .D(n4), .E(n461), .Z(
        \chs_out_f[3][DATA][28] ) );
  HS65_LS_AOI222X2 U494 ( .A(n75), .B(\chs_in_f[2][DATA][28] ), .C(n43), .D(
        \chs_in_f[0][DATA][28] ), .E(n59), .F(\chs_in_f[1][DATA][28] ), .Z(
        n461) );
  HS65_LS_OAI212X5 U495 ( .A(n271), .B(n31), .C(n306), .D(n4), .E(n462), .Z(
        \chs_out_f[3][DATA][29] ) );
  HS65_LS_AOI222X2 U496 ( .A(n75), .B(\chs_in_f[2][DATA][29] ), .C(n43), .D(
        \chs_in_f[0][DATA][29] ), .E(n59), .F(\chs_in_f[1][DATA][29] ), .Z(
        n462) );
  HS65_LS_OAI212X5 U497 ( .A(n270), .B(n31), .C(n305), .D(n4), .E(n464), .Z(
        \chs_out_f[3][DATA][30] ) );
  HS65_LS_AOI222X2 U498 ( .A(n75), .B(\chs_in_f[2][DATA][30] ), .C(n43), .D(
        \chs_in_f[0][DATA][30] ), .E(n59), .F(\chs_in_f[1][DATA][30] ), .Z(
        n464) );
  HS65_LS_OAI212X5 U499 ( .A(n269), .B(n31), .C(n304), .D(n5), .E(n465), .Z(
        \chs_out_f[3][DATA][31] ) );
  HS65_LS_AOI222X2 U500 ( .A(n76), .B(\chs_in_f[2][DATA][31] ), .C(n44), .D(
        \chs_in_f[0][DATA][31] ), .E(n60), .F(\chs_in_f[1][DATA][31] ), .Z(
        n465) );
  HS65_LS_OAI212X5 U501 ( .A(n268), .B(n31), .C(n303), .D(n5), .E(n466), .Z(
        \chs_out_f[3][DATA][32] ) );
  HS65_LS_AOI222X2 U502 ( .A(n76), .B(\chs_in_f[2][DATA][32] ), .C(n44), .D(
        \chs_in_f[0][DATA][32] ), .E(n60), .F(\chs_in_f[1][DATA][32] ), .Z(
        n466) );
  HS65_LS_OAI212X5 U503 ( .A(n267), .B(n32), .C(n302), .D(n5), .E(n467), .Z(
        \chs_out_f[3][DATA][33] ) );
  HS65_LS_AOI222X2 U504 ( .A(n76), .B(\chs_in_f[2][DATA][33] ), .C(n44), .D(
        \chs_in_f[0][DATA][33] ), .E(n60), .F(\chs_in_f[1][DATA][33] ), .Z(
        n467) );
  HS65_LS_OAI212X5 U505 ( .A(n266), .B(n32), .C(n301), .D(n5), .E(n468), .Z(
        \chs_out_f[3][DATA][34] ) );
  HS65_LS_OAI212X5 U506 ( .A(n20), .B(n266), .C(n17), .D(n301), .E(n503), .Z(
        \chs_out_f[4][DATA][34] ) );
  HS65_LS_OAI212X5 U507 ( .A(n266), .B(n23), .C(n301), .D(n8), .E(n433), .Z(
        \chs_out_f[2][DATA][34] ) );
  HS65_LS_OAI212X5 U508 ( .A(n266), .B(n26), .C(n301), .D(n11), .E(n398), .Z(
        \chs_out_f[1][DATA][34] ) );
  HS65_LS_OAI212X5 U509 ( .A(n266), .B(n29), .C(n301), .D(n14), .E(n363), .Z(
        \chs_out_f[0][DATA][34] ) );
  HS65_LS_IVX9 U510 ( .A(\switch_sel[4][4] ), .Z(n260) );
  HS65_LS_IVX9 U511 ( .A(\switch_sel[3][3] ), .Z(n265) );
endmodule


module latch_controller_0_5 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_0_000000000_5 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, n3, n5, n6, n7, n8, n9, n10;
  assign N0 = preset;

  latch_controller_0_5 controller ( .preset(n6), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLQX9 type_out_reg ( .D(N4), .GN(n8), .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U8 ( .A(\left_in[DATA][34] ), .B(n3), .Z(n9) );
  HS65_LS_AND2X4 U7 ( .A(1'b0), .B(n7), .Z(n10) );
  HS65_LS_OR2X9 U9 ( .A(n10), .B(n9), .Z(N4) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(N39), .Q(\right_out[DATA][33] )
         );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(N38), .Q(\right_out[DATA][32] )
         );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(N37), .Q(\right_out[DATA][31] )
         );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(N36), .Q(\right_out[DATA][30] )
         );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(N35), .Q(\right_out[DATA][29] )
         );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(N34), .Q(\right_out[DATA][28] )
         );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(N33), .Q(\right_out[DATA][27] )
         );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(N32), .Q(\right_out[DATA][26] )
         );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(N31), .Q(\right_out[DATA][25] )
         );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(N30), .Q(\right_out[DATA][24] )
         );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(N29), .Q(\right_out[DATA][23] )
         );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(N28), .Q(\right_out[DATA][22] )
         );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(N27), .Q(\right_out[DATA][21] )
         );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(N26), .Q(\right_out[DATA][20] )
         );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(N25), .Q(\right_out[DATA][19] )
         );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(N24), .Q(\right_out[DATA][18] )
         );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(N23), .Q(\right_out[DATA][17] )
         );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(N22), .Q(\right_out[DATA][16] )
         );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(N21), .Q(\right_out[DATA][15] )
         );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(N20), .Q(\right_out[DATA][14] )
         );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(N19), .Q(\right_out[DATA][13] )
         );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(N18), .Q(\right_out[DATA][12] )
         );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(N17), .Q(\right_out[DATA][11] )
         );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(N16), .Q(\right_out[DATA][10] )
         );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(N15), .Q(\right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(N14), .Q(\right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(N13), .Q(\right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(N12), .Q(\right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(N11), .Q(\right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(N10), .Q(\right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(N9), .Q(\right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(N8), .Q(\right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(N7), .Q(\right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(N6), .Q(\right_out[DATA][0] ) );
  HS65_LS_BFX9 U3 ( .A(N0), .Z(n6) );
  HS65_LS_IVX9 U4 ( .A(n6), .Z(n3) );
  HS65_LS_IVX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_NOR2X6 U6 ( .A(lt_enable), .B(n7), .Z(n8) );
  HS65_LS_AND2X4 U10 ( .A(\left_in[DATA][9] ), .B(n3), .Z(N15) );
  HS65_LS_AND2X4 U11 ( .A(\left_in[DATA][0] ), .B(n3), .Z(N6) );
  HS65_LS_AND2X4 U12 ( .A(\left_in[DATA][1] ), .B(n5), .Z(N7) );
  HS65_LS_AND2X4 U13 ( .A(\left_in[DATA][2] ), .B(n3), .Z(N8) );
  HS65_LS_AND2X4 U14 ( .A(\left_in[DATA][3] ), .B(n5), .Z(N9) );
  HS65_LS_AND2X4 U15 ( .A(\left_in[DATA][4] ), .B(n3), .Z(N10) );
  HS65_LS_AND2X4 U16 ( .A(\left_in[DATA][5] ), .B(n3), .Z(N11) );
  HS65_LS_AND2X4 U17 ( .A(\left_in[DATA][6] ), .B(n3), .Z(N12) );
  HS65_LS_AND2X4 U18 ( .A(\left_in[DATA][7] ), .B(n3), .Z(N13) );
  HS65_LS_AND2X4 U19 ( .A(\left_in[DATA][8] ), .B(n3), .Z(N14) );
  HS65_LS_AND2X4 U20 ( .A(\left_in[DATA][10] ), .B(n3), .Z(N16) );
  HS65_LS_AND2X4 U21 ( .A(\left_in[DATA][11] ), .B(n3), .Z(N17) );
  HS65_LS_AND2X4 U22 ( .A(\left_in[DATA][12] ), .B(n3), .Z(N18) );
  HS65_LS_AND2X4 U23 ( .A(\left_in[DATA][13] ), .B(n3), .Z(N19) );
  HS65_LS_AND2X4 U24 ( .A(\left_in[DATA][14] ), .B(n3), .Z(N20) );
  HS65_LS_AND2X4 U25 ( .A(\left_in[DATA][15] ), .B(n3), .Z(N21) );
  HS65_LS_AND2X4 U26 ( .A(\left_in[DATA][16] ), .B(n3), .Z(N22) );
  HS65_LS_AND2X4 U27 ( .A(\left_in[DATA][17] ), .B(n5), .Z(N23) );
  HS65_LS_AND2X4 U28 ( .A(\left_in[DATA][18] ), .B(n5), .Z(N24) );
  HS65_LS_AND2X4 U29 ( .A(\left_in[DATA][19] ), .B(n5), .Z(N25) );
  HS65_LS_AND2X4 U30 ( .A(\left_in[DATA][20] ), .B(n5), .Z(N26) );
  HS65_LS_AND2X4 U31 ( .A(\left_in[DATA][21] ), .B(n5), .Z(N27) );
  HS65_LS_AND2X4 U32 ( .A(\left_in[DATA][22] ), .B(n5), .Z(N28) );
  HS65_LS_AND2X4 U33 ( .A(\left_in[DATA][23] ), .B(n5), .Z(N29) );
  HS65_LS_AND2X4 U34 ( .A(\left_in[DATA][24] ), .B(n5), .Z(N30) );
  HS65_LS_AND2X4 U35 ( .A(\left_in[DATA][25] ), .B(n5), .Z(N31) );
  HS65_LS_AND2X4 U36 ( .A(\left_in[DATA][26] ), .B(n5), .Z(N32) );
  HS65_LS_AND2X4 U37 ( .A(\left_in[DATA][27] ), .B(n5), .Z(N33) );
  HS65_LS_AND2X4 U38 ( .A(\left_in[DATA][28] ), .B(n5), .Z(N34) );
  HS65_LS_AND2X4 U39 ( .A(\left_in[DATA][29] ), .B(n5), .Z(N35) );
  HS65_LS_AND2X4 U40 ( .A(\left_in[DATA][30] ), .B(n3), .Z(N36) );
  HS65_LS_AND2X4 U41 ( .A(\left_in[DATA][31] ), .B(n5), .Z(N37) );
  HS65_LS_AND2X4 U42 ( .A(\left_in[DATA][32] ), .B(n3), .Z(N38) );
  HS65_LS_AND2X4 U43 ( .A(\left_in[DATA][33] ), .B(n5), .Z(N39) );
  HS65_LS_BFX9 U44 ( .A(N0), .Z(n7) );
  HS65_LS_NAND2X7 U45 ( .A(\right_out[DATA][34] ), .B(n8), .Z(N5) );
endmodule


module latch_controller_0_4 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_0_000000000_4 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, n3, n5, n6, n7, n8, n9, n10;
  assign N0 = preset;

  latch_controller_0_4 controller ( .preset(n6), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLQX9 type_out_reg ( .D(N4), .GN(n8), .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U7 ( .A(1'b0), .B(n7), .Z(n10) );
  HS65_LS_OR2X9 U9 ( .A(n10), .B(n9), .Z(N4) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(N39), .Q(\right_out[DATA][33] )
         );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(N38), .Q(\right_out[DATA][32] )
         );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(N37), .Q(\right_out[DATA][31] )
         );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(N36), .Q(\right_out[DATA][30] )
         );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(N35), .Q(\right_out[DATA][29] )
         );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(N34), .Q(\right_out[DATA][28] )
         );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(N33), .Q(\right_out[DATA][27] )
         );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(N32), .Q(\right_out[DATA][26] )
         );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(N31), .Q(\right_out[DATA][25] )
         );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(N30), .Q(\right_out[DATA][24] )
         );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(N29), .Q(\right_out[DATA][23] )
         );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(N28), .Q(\right_out[DATA][22] )
         );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(N27), .Q(\right_out[DATA][21] )
         );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(N26), .Q(\right_out[DATA][20] )
         );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(N25), .Q(\right_out[DATA][19] )
         );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(N24), .Q(\right_out[DATA][18] )
         );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(N23), .Q(\right_out[DATA][17] )
         );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(N22), .Q(\right_out[DATA][16] )
         );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(N21), .Q(\right_out[DATA][15] )
         );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(N20), .Q(\right_out[DATA][14] )
         );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(N19), .Q(\right_out[DATA][13] )
         );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(N18), .Q(\right_out[DATA][12] )
         );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(N17), .Q(\right_out[DATA][11] )
         );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(N16), .Q(\right_out[DATA][10] )
         );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(N15), .Q(\right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(N14), .Q(\right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(N13), .Q(\right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(N12), .Q(\right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(N11), .Q(\right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(N10), .Q(\right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(N9), .Q(\right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(N8), .Q(\right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(N7), .Q(\right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(N6), .Q(\right_out[DATA][0] ) );
  HS65_LS_AND2X4 U8 ( .A(\left_in[DATA][34] ), .B(n3), .Z(n9) );
  HS65_LS_BFX9 U3 ( .A(N0), .Z(n6) );
  HS65_LS_IVX9 U4 ( .A(n6), .Z(n3) );
  HS65_LS_IVX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_NOR2X6 U6 ( .A(lt_enable), .B(n7), .Z(n8) );
  HS65_LS_AND2X4 U10 ( .A(\left_in[DATA][9] ), .B(n3), .Z(N15) );
  HS65_LS_AND2X4 U11 ( .A(\left_in[DATA][0] ), .B(n5), .Z(N6) );
  HS65_LS_AND2X4 U12 ( .A(\left_in[DATA][1] ), .B(n3), .Z(N7) );
  HS65_LS_AND2X4 U13 ( .A(\left_in[DATA][2] ), .B(n5), .Z(N8) );
  HS65_LS_AND2X4 U14 ( .A(\left_in[DATA][3] ), .B(n3), .Z(N9) );
  HS65_LS_AND2X4 U15 ( .A(\left_in[DATA][4] ), .B(n3), .Z(N10) );
  HS65_LS_AND2X4 U16 ( .A(\left_in[DATA][5] ), .B(n3), .Z(N11) );
  HS65_LS_AND2X4 U17 ( .A(\left_in[DATA][6] ), .B(n3), .Z(N12) );
  HS65_LS_AND2X4 U18 ( .A(\left_in[DATA][7] ), .B(n3), .Z(N13) );
  HS65_LS_AND2X4 U19 ( .A(\left_in[DATA][8] ), .B(n3), .Z(N14) );
  HS65_LS_AND2X4 U20 ( .A(\left_in[DATA][10] ), .B(n3), .Z(N16) );
  HS65_LS_AND2X4 U21 ( .A(\left_in[DATA][11] ), .B(n3), .Z(N17) );
  HS65_LS_AND2X4 U22 ( .A(\left_in[DATA][12] ), .B(n3), .Z(N18) );
  HS65_LS_AND2X4 U23 ( .A(\left_in[DATA][13] ), .B(n3), .Z(N19) );
  HS65_LS_AND2X4 U24 ( .A(\left_in[DATA][14] ), .B(n3), .Z(N20) );
  HS65_LS_AND2X4 U25 ( .A(\left_in[DATA][15] ), .B(n3), .Z(N21) );
  HS65_LS_AND2X4 U26 ( .A(\left_in[DATA][16] ), .B(n3), .Z(N22) );
  HS65_LS_AND2X4 U27 ( .A(\left_in[DATA][17] ), .B(n5), .Z(N23) );
  HS65_LS_AND2X4 U28 ( .A(\left_in[DATA][18] ), .B(n5), .Z(N24) );
  HS65_LS_AND2X4 U29 ( .A(\left_in[DATA][19] ), .B(n5), .Z(N25) );
  HS65_LS_AND2X4 U30 ( .A(\left_in[DATA][20] ), .B(n5), .Z(N26) );
  HS65_LS_AND2X4 U31 ( .A(\left_in[DATA][21] ), .B(n5), .Z(N27) );
  HS65_LS_AND2X4 U32 ( .A(\left_in[DATA][22] ), .B(n5), .Z(N28) );
  HS65_LS_AND2X4 U33 ( .A(\left_in[DATA][23] ), .B(n5), .Z(N29) );
  HS65_LS_AND2X4 U34 ( .A(\left_in[DATA][24] ), .B(n5), .Z(N30) );
  HS65_LS_AND2X4 U35 ( .A(\left_in[DATA][25] ), .B(n5), .Z(N31) );
  HS65_LS_AND2X4 U36 ( .A(\left_in[DATA][26] ), .B(n5), .Z(N32) );
  HS65_LS_AND2X4 U37 ( .A(\left_in[DATA][27] ), .B(n5), .Z(N33) );
  HS65_LS_AND2X4 U38 ( .A(\left_in[DATA][28] ), .B(n5), .Z(N34) );
  HS65_LS_AND2X4 U39 ( .A(\left_in[DATA][29] ), .B(n5), .Z(N35) );
  HS65_LS_AND2X4 U40 ( .A(\left_in[DATA][30] ), .B(n5), .Z(N36) );
  HS65_LS_AND2X4 U41 ( .A(\left_in[DATA][31] ), .B(n3), .Z(N37) );
  HS65_LS_AND2X4 U42 ( .A(\left_in[DATA][32] ), .B(n5), .Z(N38) );
  HS65_LS_AND2X4 U43 ( .A(\left_in[DATA][33] ), .B(n3), .Z(N39) );
  HS65_LS_BFX9 U44 ( .A(N0), .Z(n7) );
  HS65_LS_NAND2X7 U45 ( .A(\right_out[DATA][34] ), .B(n8), .Z(N5) );
endmodule


module latch_controller_0_3 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_0_000000000_3 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, n3, n5, n6, n7, n8, n9, n10;
  assign N0 = preset;

  latch_controller_0_3 controller ( .preset(n6), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLQX9 type_out_reg ( .D(N4), .GN(n8), .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U8 ( .A(\left_in[DATA][34] ), .B(n3), .Z(n9) );
  HS65_LS_AND2X4 U7 ( .A(1'b0), .B(n7), .Z(n10) );
  HS65_LS_OR2X9 U9 ( .A(n10), .B(n9), .Z(N4) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(N39), .Q(\right_out[DATA][33] )
         );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(N38), .Q(\right_out[DATA][32] )
         );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(N37), .Q(\right_out[DATA][31] )
         );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(N36), .Q(\right_out[DATA][30] )
         );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(N35), .Q(\right_out[DATA][29] )
         );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(N34), .Q(\right_out[DATA][28] )
         );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(N33), .Q(\right_out[DATA][27] )
         );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(N32), .Q(\right_out[DATA][26] )
         );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(N31), .Q(\right_out[DATA][25] )
         );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(N30), .Q(\right_out[DATA][24] )
         );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(N29), .Q(\right_out[DATA][23] )
         );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(N28), .Q(\right_out[DATA][22] )
         );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(N27), .Q(\right_out[DATA][21] )
         );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(N26), .Q(\right_out[DATA][20] )
         );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(N25), .Q(\right_out[DATA][19] )
         );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(N24), .Q(\right_out[DATA][18] )
         );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(N23), .Q(\right_out[DATA][17] )
         );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(N22), .Q(\right_out[DATA][16] )
         );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(N21), .Q(\right_out[DATA][15] )
         );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(N20), .Q(\right_out[DATA][14] )
         );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(N19), .Q(\right_out[DATA][13] )
         );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(N18), .Q(\right_out[DATA][12] )
         );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(N17), .Q(\right_out[DATA][11] )
         );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(N16), .Q(\right_out[DATA][10] )
         );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(N15), .Q(\right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(N14), .Q(\right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(N13), .Q(\right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(N12), .Q(\right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(N11), .Q(\right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(N10), .Q(\right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(N9), .Q(\right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(N8), .Q(\right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(N7), .Q(\right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(N6), .Q(\right_out[DATA][0] ) );
  HS65_LS_BFX9 U3 ( .A(N0), .Z(n6) );
  HS65_LS_IVX9 U4 ( .A(n6), .Z(n3) );
  HS65_LS_IVX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_NOR2X6 U6 ( .A(lt_enable), .B(n7), .Z(n8) );
  HS65_LS_AND2X4 U10 ( .A(\left_in[DATA][9] ), .B(n3), .Z(N15) );
  HS65_LS_AND2X4 U11 ( .A(\left_in[DATA][0] ), .B(n3), .Z(N6) );
  HS65_LS_AND2X4 U12 ( .A(\left_in[DATA][1] ), .B(n5), .Z(N7) );
  HS65_LS_AND2X4 U13 ( .A(\left_in[DATA][2] ), .B(n3), .Z(N8) );
  HS65_LS_AND2X4 U14 ( .A(\left_in[DATA][10] ), .B(n3), .Z(N16) );
  HS65_LS_AND2X4 U15 ( .A(\left_in[DATA][11] ), .B(n3), .Z(N17) );
  HS65_LS_AND2X4 U16 ( .A(\left_in[DATA][12] ), .B(n3), .Z(N18) );
  HS65_LS_AND2X4 U17 ( .A(\left_in[DATA][13] ), .B(n3), .Z(N19) );
  HS65_LS_AND2X4 U18 ( .A(\left_in[DATA][14] ), .B(n3), .Z(N20) );
  HS65_LS_AND2X4 U19 ( .A(\left_in[DATA][15] ), .B(n3), .Z(N21) );
  HS65_LS_AND2X4 U20 ( .A(\left_in[DATA][16] ), .B(n3), .Z(N22) );
  HS65_LS_AND2X4 U21 ( .A(\left_in[DATA][17] ), .B(n5), .Z(N23) );
  HS65_LS_AND2X4 U22 ( .A(\left_in[DATA][18] ), .B(n5), .Z(N24) );
  HS65_LS_AND2X4 U23 ( .A(\left_in[DATA][19] ), .B(n5), .Z(N25) );
  HS65_LS_AND2X4 U24 ( .A(\left_in[DATA][20] ), .B(n5), .Z(N26) );
  HS65_LS_AND2X4 U25 ( .A(\left_in[DATA][21] ), .B(n5), .Z(N27) );
  HS65_LS_AND2X4 U26 ( .A(\left_in[DATA][22] ), .B(n5), .Z(N28) );
  HS65_LS_AND2X4 U27 ( .A(\left_in[DATA][23] ), .B(n5), .Z(N29) );
  HS65_LS_AND2X4 U28 ( .A(\left_in[DATA][24] ), .B(n5), .Z(N30) );
  HS65_LS_AND2X4 U29 ( .A(\left_in[DATA][25] ), .B(n5), .Z(N31) );
  HS65_LS_AND2X4 U30 ( .A(\left_in[DATA][26] ), .B(n5), .Z(N32) );
  HS65_LS_AND2X4 U31 ( .A(\left_in[DATA][27] ), .B(n5), .Z(N33) );
  HS65_LS_AND2X4 U32 ( .A(\left_in[DATA][28] ), .B(n5), .Z(N34) );
  HS65_LS_AND2X4 U33 ( .A(\left_in[DATA][29] ), .B(n5), .Z(N35) );
  HS65_LS_AND2X4 U34 ( .A(\left_in[DATA][30] ), .B(n5), .Z(N36) );
  HS65_LS_AND2X4 U35 ( .A(\left_in[DATA][31] ), .B(n3), .Z(N37) );
  HS65_LS_AND2X4 U36 ( .A(\left_in[DATA][32] ), .B(n5), .Z(N38) );
  HS65_LS_AND2X4 U37 ( .A(\left_in[DATA][3] ), .B(n3), .Z(N9) );
  HS65_LS_AND2X4 U38 ( .A(\left_in[DATA][4] ), .B(n3), .Z(N10) );
  HS65_LS_AND2X4 U39 ( .A(\left_in[DATA][5] ), .B(n3), .Z(N11) );
  HS65_LS_AND2X4 U40 ( .A(\left_in[DATA][6] ), .B(n3), .Z(N12) );
  HS65_LS_AND2X4 U41 ( .A(\left_in[DATA][7] ), .B(n3), .Z(N13) );
  HS65_LS_AND2X4 U42 ( .A(\left_in[DATA][8] ), .B(n3), .Z(N14) );
  HS65_LS_AND2X4 U43 ( .A(\left_in[DATA][33] ), .B(n5), .Z(N39) );
  HS65_LS_BFX9 U44 ( .A(N0), .Z(n7) );
  HS65_LS_NAND2X7 U45 ( .A(\right_out[DATA][34] ), .B(n8), .Z(N5) );
endmodule


module latch_controller_0_2 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_0_000000000_2 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, n3, n5, n6, n7, n8, n9, n10;
  assign N0 = preset;

  latch_controller_0_2 controller ( .preset(n6), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLQX9 type_out_reg ( .D(N4), .GN(n8), .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U8 ( .A(\left_in[DATA][34] ), .B(n3), .Z(n9) );
  HS65_LS_AND2X4 U7 ( .A(1'b0), .B(n7), .Z(n10) );
  HS65_LS_OR2X9 U9 ( .A(n10), .B(n9), .Z(N4) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(N39), .Q(\right_out[DATA][33] )
         );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(N38), .Q(\right_out[DATA][32] )
         );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(N37), .Q(\right_out[DATA][31] )
         );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(N36), .Q(\right_out[DATA][30] )
         );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(N35), .Q(\right_out[DATA][29] )
         );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(N34), .Q(\right_out[DATA][28] )
         );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(N33), .Q(\right_out[DATA][27] )
         );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(N32), .Q(\right_out[DATA][26] )
         );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(N31), .Q(\right_out[DATA][25] )
         );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(N30), .Q(\right_out[DATA][24] )
         );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(N29), .Q(\right_out[DATA][23] )
         );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(N28), .Q(\right_out[DATA][22] )
         );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(N27), .Q(\right_out[DATA][21] )
         );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(N26), .Q(\right_out[DATA][20] )
         );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(N25), .Q(\right_out[DATA][19] )
         );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(N24), .Q(\right_out[DATA][18] )
         );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(N23), .Q(\right_out[DATA][17] )
         );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(N22), .Q(\right_out[DATA][16] )
         );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(N21), .Q(\right_out[DATA][15] )
         );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(N20), .Q(\right_out[DATA][14] )
         );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(N19), .Q(\right_out[DATA][13] )
         );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(N18), .Q(\right_out[DATA][12] )
         );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(N17), .Q(\right_out[DATA][11] )
         );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(N16), .Q(\right_out[DATA][10] )
         );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(N15), .Q(\right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(N14), .Q(\right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(N13), .Q(\right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(N12), .Q(\right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(N11), .Q(\right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(N10), .Q(\right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(N9), .Q(\right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(N8), .Q(\right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(N7), .Q(\right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(N6), .Q(\right_out[DATA][0] ) );
  HS65_LS_BFX9 U3 ( .A(N0), .Z(n6) );
  HS65_LS_IVX9 U4 ( .A(n6), .Z(n3) );
  HS65_LS_IVX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_NOR2X6 U6 ( .A(lt_enable), .B(n7), .Z(n8) );
  HS65_LS_AND2X4 U10 ( .A(\left_in[DATA][9] ), .B(n3), .Z(N15) );
  HS65_LS_AND2X4 U11 ( .A(\left_in[DATA][0] ), .B(n3), .Z(N6) );
  HS65_LS_AND2X4 U12 ( .A(\left_in[DATA][1] ), .B(n5), .Z(N7) );
  HS65_LS_AND2X4 U13 ( .A(\left_in[DATA][2] ), .B(n3), .Z(N8) );
  HS65_LS_AND2X4 U14 ( .A(\left_in[DATA][10] ), .B(n3), .Z(N16) );
  HS65_LS_AND2X4 U15 ( .A(\left_in[DATA][11] ), .B(n3), .Z(N17) );
  HS65_LS_AND2X4 U16 ( .A(\left_in[DATA][12] ), .B(n3), .Z(N18) );
  HS65_LS_AND2X4 U17 ( .A(\left_in[DATA][13] ), .B(n3), .Z(N19) );
  HS65_LS_AND2X4 U18 ( .A(\left_in[DATA][14] ), .B(n3), .Z(N20) );
  HS65_LS_AND2X4 U19 ( .A(\left_in[DATA][15] ), .B(n3), .Z(N21) );
  HS65_LS_AND2X4 U20 ( .A(\left_in[DATA][16] ), .B(n3), .Z(N22) );
  HS65_LS_AND2X4 U21 ( .A(\left_in[DATA][17] ), .B(n5), .Z(N23) );
  HS65_LS_AND2X4 U22 ( .A(\left_in[DATA][18] ), .B(n5), .Z(N24) );
  HS65_LS_AND2X4 U23 ( .A(\left_in[DATA][19] ), .B(n5), .Z(N25) );
  HS65_LS_AND2X4 U24 ( .A(\left_in[DATA][20] ), .B(n5), .Z(N26) );
  HS65_LS_AND2X4 U25 ( .A(\left_in[DATA][21] ), .B(n5), .Z(N27) );
  HS65_LS_AND2X4 U26 ( .A(\left_in[DATA][22] ), .B(n5), .Z(N28) );
  HS65_LS_AND2X4 U27 ( .A(\left_in[DATA][23] ), .B(n5), .Z(N29) );
  HS65_LS_AND2X4 U28 ( .A(\left_in[DATA][24] ), .B(n5), .Z(N30) );
  HS65_LS_AND2X4 U29 ( .A(\left_in[DATA][25] ), .B(n5), .Z(N31) );
  HS65_LS_AND2X4 U30 ( .A(\left_in[DATA][26] ), .B(n5), .Z(N32) );
  HS65_LS_AND2X4 U31 ( .A(\left_in[DATA][27] ), .B(n5), .Z(N33) );
  HS65_LS_AND2X4 U32 ( .A(\left_in[DATA][28] ), .B(n5), .Z(N34) );
  HS65_LS_AND2X4 U33 ( .A(\left_in[DATA][29] ), .B(n5), .Z(N35) );
  HS65_LS_AND2X4 U34 ( .A(\left_in[DATA][30] ), .B(n5), .Z(N36) );
  HS65_LS_AND2X4 U35 ( .A(\left_in[DATA][31] ), .B(n3), .Z(N37) );
  HS65_LS_AND2X4 U36 ( .A(\left_in[DATA][32] ), .B(n5), .Z(N38) );
  HS65_LS_AND2X4 U37 ( .A(\left_in[DATA][3] ), .B(n3), .Z(N9) );
  HS65_LS_AND2X4 U38 ( .A(\left_in[DATA][4] ), .B(n3), .Z(N10) );
  HS65_LS_AND2X4 U39 ( .A(\left_in[DATA][5] ), .B(n3), .Z(N11) );
  HS65_LS_AND2X4 U40 ( .A(\left_in[DATA][6] ), .B(n3), .Z(N12) );
  HS65_LS_AND2X4 U41 ( .A(\left_in[DATA][7] ), .B(n3), .Z(N13) );
  HS65_LS_AND2X4 U42 ( .A(\left_in[DATA][8] ), .B(n3), .Z(N14) );
  HS65_LS_AND2X4 U43 ( .A(\left_in[DATA][33] ), .B(n5), .Z(N39) );
  HS65_LS_BFX9 U44 ( .A(N0), .Z(n7) );
  HS65_LS_NAND2X7 U45 ( .A(\right_out[DATA][34] ), .B(n8), .Z(N5) );
endmodule


module latch_controller_0_1 ( preset, Rin, Ain, Rout, Aout, lt_en );
  input preset, Rin, Aout;
  output Ain, Rout, lt_en;
  wire   N2, Ain, N4, N5;
  assign Rout = Ain;

  HS65_LS_LDHQX9 r_next_reg ( .G(N4), .D(N5), .Q(Ain) );
  HS65_LS_IVX9 I_0 ( .A(N2), .Z(lt_en) );
  HS65_LS_OR2X9 U3 ( .A(Rin), .B(preset), .Z(N5) );
  HS65_LS_OR2X9 U4 ( .A(lt_en), .B(preset), .Z(N4) );
  HS65_LSS_XOR2X6 U5 ( .A(Ain), .B(Aout), .Z(N2) );
endmodule


module channel_latch_0_000000000_1 ( preset, .left_in({\left_in[REQ] , 
        \left_in[DATA][34] , \left_in[DATA][33] , \left_in[DATA][32] , 
        \left_in[DATA][31] , \left_in[DATA][30] , \left_in[DATA][29] , 
        \left_in[DATA][28] , \left_in[DATA][27] , \left_in[DATA][26] , 
        \left_in[DATA][25] , \left_in[DATA][24] , \left_in[DATA][23] , 
        \left_in[DATA][22] , \left_in[DATA][21] , \left_in[DATA][20] , 
        \left_in[DATA][19] , \left_in[DATA][18] , \left_in[DATA][17] , 
        \left_in[DATA][16] , \left_in[DATA][15] , \left_in[DATA][14] , 
        \left_in[DATA][13] , \left_in[DATA][12] , \left_in[DATA][11] , 
        \left_in[DATA][10] , \left_in[DATA][9] , \left_in[DATA][8] , 
        \left_in[DATA][7] , \left_in[DATA][6] , \left_in[DATA][5] , 
        \left_in[DATA][4] , \left_in[DATA][3] , \left_in[DATA][2] , 
        \left_in[DATA][1] , \left_in[DATA][0] }), .left_out(\left_out[ACK] ), 
    .right_out({\right_out[REQ] , \right_out[DATA][34] , \right_out[DATA][33] , 
        \right_out[DATA][32] , \right_out[DATA][31] , \right_out[DATA][30] , 
        \right_out[DATA][29] , \right_out[DATA][28] , \right_out[DATA][27] , 
        \right_out[DATA][26] , \right_out[DATA][25] , \right_out[DATA][24] , 
        \right_out[DATA][23] , \right_out[DATA][22] , \right_out[DATA][21] , 
        \right_out[DATA][20] , \right_out[DATA][19] , \right_out[DATA][18] , 
        \right_out[DATA][17] , \right_out[DATA][16] , \right_out[DATA][15] , 
        \right_out[DATA][14] , \right_out[DATA][13] , \right_out[DATA][12] , 
        \right_out[DATA][11] , \right_out[DATA][10] , \right_out[DATA][9] , 
        \right_out[DATA][8] , \right_out[DATA][7] , \right_out[DATA][6] , 
        \right_out[DATA][5] , \right_out[DATA][4] , \right_out[DATA][3] , 
        \right_out[DATA][2] , \right_out[DATA][1] , \right_out[DATA][0] }), 
    .right_in(\right_in[ACK] ), lt_enable );
  input preset, \left_in[REQ] , \left_in[DATA][34] , \left_in[DATA][33] ,
         \left_in[DATA][32] , \left_in[DATA][31] , \left_in[DATA][30] ,
         \left_in[DATA][29] , \left_in[DATA][28] , \left_in[DATA][27] ,
         \left_in[DATA][26] , \left_in[DATA][25] , \left_in[DATA][24] ,
         \left_in[DATA][23] , \left_in[DATA][22] , \left_in[DATA][21] ,
         \left_in[DATA][20] , \left_in[DATA][19] , \left_in[DATA][18] ,
         \left_in[DATA][17] , \left_in[DATA][16] , \left_in[DATA][15] ,
         \left_in[DATA][14] , \left_in[DATA][13] , \left_in[DATA][12] ,
         \left_in[DATA][11] , \left_in[DATA][10] , \left_in[DATA][9] ,
         \left_in[DATA][8] , \left_in[DATA][7] , \left_in[DATA][6] ,
         \left_in[DATA][5] , \left_in[DATA][4] , \left_in[DATA][3] ,
         \left_in[DATA][2] , \left_in[DATA][1] , \left_in[DATA][0] ,
         \right_in[ACK] ;
  output \left_out[ACK] , \right_out[REQ] , \right_out[DATA][34] ,
         \right_out[DATA][33] , \right_out[DATA][32] , \right_out[DATA][31] ,
         \right_out[DATA][30] , \right_out[DATA][29] , \right_out[DATA][28] ,
         \right_out[DATA][27] , \right_out[DATA][26] , \right_out[DATA][25] ,
         \right_out[DATA][24] , \right_out[DATA][23] , \right_out[DATA][22] ,
         \right_out[DATA][21] , \right_out[DATA][20] , \right_out[DATA][19] ,
         \right_out[DATA][18] , \right_out[DATA][17] , \right_out[DATA][16] ,
         \right_out[DATA][15] , \right_out[DATA][14] , \right_out[DATA][13] ,
         \right_out[DATA][12] , \right_out[DATA][11] , \right_out[DATA][10] ,
         \right_out[DATA][9] , \right_out[DATA][8] , \right_out[DATA][7] ,
         \right_out[DATA][6] , \right_out[DATA][5] , \right_out[DATA][4] ,
         \right_out[DATA][3] , \right_out[DATA][2] , \right_out[DATA][1] ,
         \right_out[DATA][0] , lt_enable;
  wire   N0, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, n3, n5, n6, n7, n8, n9, n10;
  assign N0 = preset;

  latch_controller_0_1 controller ( .preset(n6), .Rin(\left_in[REQ] ), .Ain(
        \left_out[ACK] ), .Rout(\right_out[REQ] ), .Aout(\right_in[ACK] ), 
        .lt_en(lt_enable) );
  HS65_LS_LDLQX9 type_out_reg ( .D(N4), .GN(n8), .Q(\right_out[DATA][34] ) );
  HS65_LS_AND2X4 U8 ( .A(\left_in[DATA][34] ), .B(n3), .Z(n9) );
  HS65_LS_AND2X4 U7 ( .A(1'b0), .B(n7), .Z(n10) );
  HS65_LS_OR2X9 U9 ( .A(n10), .B(n9), .Z(N4) );
  HS65_LS_LDHQX9 \data_reg[33]  ( .G(N5), .D(N39), .Q(\right_out[DATA][33] )
         );
  HS65_LS_LDHQX9 \data_reg[32]  ( .G(N5), .D(N38), .Q(\right_out[DATA][32] )
         );
  HS65_LS_LDHQX9 \data_reg[31]  ( .G(N5), .D(N37), .Q(\right_out[DATA][31] )
         );
  HS65_LS_LDHQX9 \data_reg[30]  ( .G(N5), .D(N36), .Q(\right_out[DATA][30] )
         );
  HS65_LS_LDHQX9 \data_reg[29]  ( .G(N5), .D(N35), .Q(\right_out[DATA][29] )
         );
  HS65_LS_LDHQX9 \data_reg[28]  ( .G(N5), .D(N34), .Q(\right_out[DATA][28] )
         );
  HS65_LS_LDHQX9 \data_reg[27]  ( .G(N5), .D(N33), .Q(\right_out[DATA][27] )
         );
  HS65_LS_LDHQX9 \data_reg[26]  ( .G(N5), .D(N32), .Q(\right_out[DATA][26] )
         );
  HS65_LS_LDHQX9 \data_reg[25]  ( .G(N5), .D(N31), .Q(\right_out[DATA][25] )
         );
  HS65_LS_LDHQX9 \data_reg[24]  ( .G(N5), .D(N30), .Q(\right_out[DATA][24] )
         );
  HS65_LS_LDHQX9 \data_reg[23]  ( .G(N5), .D(N29), .Q(\right_out[DATA][23] )
         );
  HS65_LS_LDHQX9 \data_reg[22]  ( .G(N5), .D(N28), .Q(\right_out[DATA][22] )
         );
  HS65_LS_LDHQX9 \data_reg[21]  ( .G(N5), .D(N27), .Q(\right_out[DATA][21] )
         );
  HS65_LS_LDHQX9 \data_reg[20]  ( .G(N5), .D(N26), .Q(\right_out[DATA][20] )
         );
  HS65_LS_LDHQX9 \data_reg[19]  ( .G(N5), .D(N25), .Q(\right_out[DATA][19] )
         );
  HS65_LS_LDHQX9 \data_reg[18]  ( .G(N5), .D(N24), .Q(\right_out[DATA][18] )
         );
  HS65_LS_LDHQX9 \data_reg[17]  ( .G(N5), .D(N23), .Q(\right_out[DATA][17] )
         );
  HS65_LS_LDHQX9 \data_reg[16]  ( .G(N5), .D(N22), .Q(\right_out[DATA][16] )
         );
  HS65_LS_LDHQX9 \data_reg[15]  ( .G(N5), .D(N21), .Q(\right_out[DATA][15] )
         );
  HS65_LS_LDHQX9 \data_reg[14]  ( .G(N5), .D(N20), .Q(\right_out[DATA][14] )
         );
  HS65_LS_LDHQX9 \data_reg[13]  ( .G(N5), .D(N19), .Q(\right_out[DATA][13] )
         );
  HS65_LS_LDHQX9 \data_reg[12]  ( .G(N5), .D(N18), .Q(\right_out[DATA][12] )
         );
  HS65_LS_LDHQX9 \data_reg[11]  ( .G(N5), .D(N17), .Q(\right_out[DATA][11] )
         );
  HS65_LS_LDHQX9 \data_reg[10]  ( .G(N5), .D(N16), .Q(\right_out[DATA][10] )
         );
  HS65_LS_LDHQX9 \data_reg[9]  ( .G(N5), .D(N15), .Q(\right_out[DATA][9] ) );
  HS65_LS_LDHQX9 \data_reg[8]  ( .G(N5), .D(N14), .Q(\right_out[DATA][8] ) );
  HS65_LS_LDHQX9 \data_reg[7]  ( .G(N5), .D(N13), .Q(\right_out[DATA][7] ) );
  HS65_LS_LDHQX9 \data_reg[6]  ( .G(N5), .D(N12), .Q(\right_out[DATA][6] ) );
  HS65_LS_LDHQX9 \data_reg[5]  ( .G(N5), .D(N11), .Q(\right_out[DATA][5] ) );
  HS65_LS_LDHQX9 \data_reg[4]  ( .G(N5), .D(N10), .Q(\right_out[DATA][4] ) );
  HS65_LS_LDHQX9 \data_reg[3]  ( .G(N5), .D(N9), .Q(\right_out[DATA][3] ) );
  HS65_LS_LDHQX9 \data_reg[2]  ( .G(N5), .D(N8), .Q(\right_out[DATA][2] ) );
  HS65_LS_LDHQX9 \data_reg[1]  ( .G(N5), .D(N7), .Q(\right_out[DATA][1] ) );
  HS65_LS_LDHQX9 \data_reg[0]  ( .G(N5), .D(N6), .Q(\right_out[DATA][0] ) );
  HS65_LS_AND2X4 U3 ( .A(\left_in[DATA][16] ), .B(n3), .Z(N22) );
  HS65_LS_AND2X4 U4 ( .A(\left_in[DATA][4] ), .B(n3), .Z(N10) );
  HS65_LS_AND2X4 U5 ( .A(\left_in[DATA][5] ), .B(n3), .Z(N11) );
  HS65_LS_AND2X4 U6 ( .A(\left_in[DATA][6] ), .B(n3), .Z(N12) );
  HS65_LS_AND2X4 U10 ( .A(\left_in[DATA][7] ), .B(n3), .Z(N13) );
  HS65_LS_AND2X4 U11 ( .A(\left_in[DATA][8] ), .B(n3), .Z(N14) );
  HS65_LS_AND2X4 U12 ( .A(\left_in[DATA][10] ), .B(n3), .Z(N16) );
  HS65_LS_AND2X4 U13 ( .A(\left_in[DATA][11] ), .B(n3), .Z(N17) );
  HS65_LS_AND2X4 U14 ( .A(\left_in[DATA][12] ), .B(n3), .Z(N18) );
  HS65_LS_AND2X4 U15 ( .A(\left_in[DATA][13] ), .B(n3), .Z(N19) );
  HS65_LS_AND2X4 U16 ( .A(\left_in[DATA][14] ), .B(n3), .Z(N20) );
  HS65_LS_AND2X4 U17 ( .A(\left_in[DATA][15] ), .B(n3), .Z(N21) );
  HS65_LS_AND2X4 U18 ( .A(\left_in[DATA][17] ), .B(n5), .Z(N23) );
  HS65_LS_AND2X4 U19 ( .A(\left_in[DATA][18] ), .B(n5), .Z(N24) );
  HS65_LS_AND2X4 U20 ( .A(\left_in[DATA][19] ), .B(n5), .Z(N25) );
  HS65_LS_AND2X4 U21 ( .A(\left_in[DATA][24] ), .B(n5), .Z(N30) );
  HS65_LS_AND2X4 U22 ( .A(\left_in[DATA][25] ), .B(n5), .Z(N31) );
  HS65_LS_AND2X4 U23 ( .A(\left_in[DATA][26] ), .B(n5), .Z(N32) );
  HS65_LS_AND2X4 U24 ( .A(\left_in[DATA][27] ), .B(n5), .Z(N33) );
  HS65_LS_AND2X4 U25 ( .A(\left_in[DATA][28] ), .B(n5), .Z(N34) );
  HS65_LS_AND2X4 U26 ( .A(\left_in[DATA][29] ), .B(n5), .Z(N35) );
  HS65_LS_AND2X4 U27 ( .A(\left_in[DATA][30] ), .B(n3), .Z(N36) );
  HS65_LS_AND2X4 U28 ( .A(\left_in[DATA][0] ), .B(n5), .Z(N6) );
  HS65_LS_AND2X4 U29 ( .A(\left_in[DATA][1] ), .B(n3), .Z(N7) );
  HS65_LS_AND2X4 U30 ( .A(\left_in[DATA][2] ), .B(n5), .Z(N8) );
  HS65_LS_BFX9 U31 ( .A(N0), .Z(n6) );
  HS65_LS_IVX9 U32 ( .A(n6), .Z(n3) );
  HS65_LS_IVX9 U33 ( .A(n6), .Z(n5) );
  HS65_LS_NOR2X6 U34 ( .A(lt_enable), .B(n7), .Z(n8) );
  HS65_LS_AND2X4 U35 ( .A(\left_in[DATA][9] ), .B(n3), .Z(N15) );
  HS65_LS_AND2X4 U36 ( .A(\left_in[DATA][20] ), .B(n5), .Z(N26) );
  HS65_LS_AND2X4 U37 ( .A(\left_in[DATA][21] ), .B(n5), .Z(N27) );
  HS65_LS_AND2X4 U38 ( .A(\left_in[DATA][22] ), .B(n5), .Z(N28) );
  HS65_LS_AND2X4 U39 ( .A(\left_in[DATA][23] ), .B(n5), .Z(N29) );
  HS65_LS_AND2X4 U40 ( .A(\left_in[DATA][31] ), .B(n3), .Z(N37) );
  HS65_LS_AND2X4 U41 ( .A(\left_in[DATA][32] ), .B(n5), .Z(N38) );
  HS65_LS_AND2X4 U42 ( .A(\left_in[DATA][3] ), .B(n3), .Z(N9) );
  HS65_LS_AND2X4 U43 ( .A(\left_in[DATA][33] ), .B(n5), .Z(N39) );
  HS65_LS_BFX9 U44 ( .A(N0), .Z(n7) );
  HS65_LS_NAND2X7 U45 ( .A(\right_out[DATA][34] ), .B(n8), .Z(N5) );
endmodule


module crossbar_stage_1 ( preset, .switch_sel({\switch_sel[4][4] , 
        \switch_sel[4][3] , \switch_sel[4][2] , \switch_sel[4][1] , 
        \switch_sel[4][0] , \switch_sel[3][4] , \switch_sel[3][3] , 
        \switch_sel[3][2] , \switch_sel[3][1] , \switch_sel[3][0] , 
        \switch_sel[2][4] , \switch_sel[2][3] , \switch_sel[2][2] , 
        \switch_sel[2][1] , \switch_sel[2][0] , \switch_sel[1][4] , 
        \switch_sel[1][3] , \switch_sel[1][2] , \switch_sel[1][1] , 
        \switch_sel[1][0] , \switch_sel[0][4] , \switch_sel[0][3] , 
        \switch_sel[0][2] , \switch_sel[0][1] , \switch_sel[0][0] }), 
    .chs_in_f({\chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] , 
        \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] , 
        \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] , 
        \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] , 
        \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] , 
        \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] , 
        \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] , 
        \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] , 
        \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] , 
        \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] , 
        \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] , 
        \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] , 
        \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] , 
        \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] , \chs_in_f[4][DATA][7] , 
        \chs_in_f[4][DATA][6] , \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] , 
        \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] , \chs_in_f[4][DATA][1] , 
        \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] , \chs_in_f[3][DATA][34] , 
        \chs_in_f[3][DATA][33] , \chs_in_f[3][DATA][32] , 
        \chs_in_f[3][DATA][31] , \chs_in_f[3][DATA][30] , 
        \chs_in_f[3][DATA][29] , \chs_in_f[3][DATA][28] , 
        \chs_in_f[3][DATA][27] , \chs_in_f[3][DATA][26] , 
        \chs_in_f[3][DATA][25] , \chs_in_f[3][DATA][24] , 
        \chs_in_f[3][DATA][23] , \chs_in_f[3][DATA][22] , 
        \chs_in_f[3][DATA][21] , \chs_in_f[3][DATA][20] , 
        \chs_in_f[3][DATA][19] , \chs_in_f[3][DATA][18] , 
        \chs_in_f[3][DATA][17] , \chs_in_f[3][DATA][16] , 
        \chs_in_f[3][DATA][15] , \chs_in_f[3][DATA][14] , 
        \chs_in_f[3][DATA][13] , \chs_in_f[3][DATA][12] , 
        \chs_in_f[3][DATA][11] , \chs_in_f[3][DATA][10] , 
        \chs_in_f[3][DATA][9] , \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] , 
        \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] , \chs_in_f[3][DATA][4] , 
        \chs_in_f[3][DATA][3] , \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] , 
        \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] , 
        \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] , 
        \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] , 
        \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] , 
        \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] , 
        \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] , 
        \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] , 
        \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] , 
        \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] , 
        \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] , 
        \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] , 
        \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] , 
        \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] , 
        \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] , \chs_in_f[2][DATA][7] , 
        \chs_in_f[2][DATA][6] , \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] , 
        \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] , \chs_in_f[2][DATA][1] , 
        \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] , \chs_in_f[1][DATA][34] , 
        \chs_in_f[1][DATA][33] , \chs_in_f[1][DATA][32] , 
        \chs_in_f[1][DATA][31] , \chs_in_f[1][DATA][30] , 
        \chs_in_f[1][DATA][29] , \chs_in_f[1][DATA][28] , 
        \chs_in_f[1][DATA][27] , \chs_in_f[1][DATA][26] , 
        \chs_in_f[1][DATA][25] , \chs_in_f[1][DATA][24] , 
        \chs_in_f[1][DATA][23] , \chs_in_f[1][DATA][22] , 
        \chs_in_f[1][DATA][21] , \chs_in_f[1][DATA][20] , 
        \chs_in_f[1][DATA][19] , \chs_in_f[1][DATA][18] , 
        \chs_in_f[1][DATA][17] , \chs_in_f[1][DATA][16] , 
        \chs_in_f[1][DATA][15] , \chs_in_f[1][DATA][14] , 
        \chs_in_f[1][DATA][13] , \chs_in_f[1][DATA][12] , 
        \chs_in_f[1][DATA][11] , \chs_in_f[1][DATA][10] , 
        \chs_in_f[1][DATA][9] , \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] , 
        \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] , \chs_in_f[1][DATA][4] , 
        \chs_in_f[1][DATA][3] , \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] , 
        \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] , 
        \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] , 
        \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] , 
        \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] , 
        \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] , 
        \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] , 
        \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] , 
        \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] , 
        \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] , 
        \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] , 
        \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] , 
        \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] , 
        \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] , 
        \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] , \chs_in_f[0][DATA][7] , 
        \chs_in_f[0][DATA][6] , \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] , 
        \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] , \chs_in_f[0][DATA][1] , 
        \chs_in_f[0][DATA][0] }), .chs_in_b({\chs_in_b[4][ACK] , 
        \chs_in_b[3][ACK] , \chs_in_b[2][ACK] , \chs_in_b[1][ACK] , 
        \chs_in_b[0][ACK] }), .latches_out_f({\latches_out_f[4][REQ] , 
        \latches_out_f[4][DATA][34] , \latches_out_f[4][DATA][33] , 
        \latches_out_f[4][DATA][32] , \latches_out_f[4][DATA][31] , 
        \latches_out_f[4][DATA][30] , \latches_out_f[4][DATA][29] , 
        \latches_out_f[4][DATA][28] , \latches_out_f[4][DATA][27] , 
        \latches_out_f[4][DATA][26] , \latches_out_f[4][DATA][25] , 
        \latches_out_f[4][DATA][24] , \latches_out_f[4][DATA][23] , 
        \latches_out_f[4][DATA][22] , \latches_out_f[4][DATA][21] , 
        \latches_out_f[4][DATA][20] , \latches_out_f[4][DATA][19] , 
        \latches_out_f[4][DATA][18] , \latches_out_f[4][DATA][17] , 
        \latches_out_f[4][DATA][16] , \latches_out_f[4][DATA][15] , 
        \latches_out_f[4][DATA][14] , \latches_out_f[4][DATA][13] , 
        \latches_out_f[4][DATA][12] , \latches_out_f[4][DATA][11] , 
        \latches_out_f[4][DATA][10] , \latches_out_f[4][DATA][9] , 
        \latches_out_f[4][DATA][8] , \latches_out_f[4][DATA][7] , 
        \latches_out_f[4][DATA][6] , \latches_out_f[4][DATA][5] , 
        \latches_out_f[4][DATA][4] , \latches_out_f[4][DATA][3] , 
        \latches_out_f[4][DATA][2] , \latches_out_f[4][DATA][1] , 
        \latches_out_f[4][DATA][0] , \latches_out_f[3][REQ] , 
        \latches_out_f[3][DATA][34] , \latches_out_f[3][DATA][33] , 
        \latches_out_f[3][DATA][32] , \latches_out_f[3][DATA][31] , 
        \latches_out_f[3][DATA][30] , \latches_out_f[3][DATA][29] , 
        \latches_out_f[3][DATA][28] , \latches_out_f[3][DATA][27] , 
        \latches_out_f[3][DATA][26] , \latches_out_f[3][DATA][25] , 
        \latches_out_f[3][DATA][24] , \latches_out_f[3][DATA][23] , 
        \latches_out_f[3][DATA][22] , \latches_out_f[3][DATA][21] , 
        \latches_out_f[3][DATA][20] , \latches_out_f[3][DATA][19] , 
        \latches_out_f[3][DATA][18] , \latches_out_f[3][DATA][17] , 
        \latches_out_f[3][DATA][16] , \latches_out_f[3][DATA][15] , 
        \latches_out_f[3][DATA][14] , \latches_out_f[3][DATA][13] , 
        \latches_out_f[3][DATA][12] , \latches_out_f[3][DATA][11] , 
        \latches_out_f[3][DATA][10] , \latches_out_f[3][DATA][9] , 
        \latches_out_f[3][DATA][8] , \latches_out_f[3][DATA][7] , 
        \latches_out_f[3][DATA][6] , \latches_out_f[3][DATA][5] , 
        \latches_out_f[3][DATA][4] , \latches_out_f[3][DATA][3] , 
        \latches_out_f[3][DATA][2] , \latches_out_f[3][DATA][1] , 
        \latches_out_f[3][DATA][0] , \latches_out_f[2][REQ] , 
        \latches_out_f[2][DATA][34] , \latches_out_f[2][DATA][33] , 
        \latches_out_f[2][DATA][32] , \latches_out_f[2][DATA][31] , 
        \latches_out_f[2][DATA][30] , \latches_out_f[2][DATA][29] , 
        \latches_out_f[2][DATA][28] , \latches_out_f[2][DATA][27] , 
        \latches_out_f[2][DATA][26] , \latches_out_f[2][DATA][25] , 
        \latches_out_f[2][DATA][24] , \latches_out_f[2][DATA][23] , 
        \latches_out_f[2][DATA][22] , \latches_out_f[2][DATA][21] , 
        \latches_out_f[2][DATA][20] , \latches_out_f[2][DATA][19] , 
        \latches_out_f[2][DATA][18] , \latches_out_f[2][DATA][17] , 
        \latches_out_f[2][DATA][16] , \latches_out_f[2][DATA][15] , 
        \latches_out_f[2][DATA][14] , \latches_out_f[2][DATA][13] , 
        \latches_out_f[2][DATA][12] , \latches_out_f[2][DATA][11] , 
        \latches_out_f[2][DATA][10] , \latches_out_f[2][DATA][9] , 
        \latches_out_f[2][DATA][8] , \latches_out_f[2][DATA][7] , 
        \latches_out_f[2][DATA][6] , \latches_out_f[2][DATA][5] , 
        \latches_out_f[2][DATA][4] , \latches_out_f[2][DATA][3] , 
        \latches_out_f[2][DATA][2] , \latches_out_f[2][DATA][1] , 
        \latches_out_f[2][DATA][0] , \latches_out_f[1][REQ] , 
        \latches_out_f[1][DATA][34] , \latches_out_f[1][DATA][33] , 
        \latches_out_f[1][DATA][32] , \latches_out_f[1][DATA][31] , 
        \latches_out_f[1][DATA][30] , \latches_out_f[1][DATA][29] , 
        \latches_out_f[1][DATA][28] , \latches_out_f[1][DATA][27] , 
        \latches_out_f[1][DATA][26] , \latches_out_f[1][DATA][25] , 
        \latches_out_f[1][DATA][24] , \latches_out_f[1][DATA][23] , 
        \latches_out_f[1][DATA][22] , \latches_out_f[1][DATA][21] , 
        \latches_out_f[1][DATA][20] , \latches_out_f[1][DATA][19] , 
        \latches_out_f[1][DATA][18] , \latches_out_f[1][DATA][17] , 
        \latches_out_f[1][DATA][16] , \latches_out_f[1][DATA][15] , 
        \latches_out_f[1][DATA][14] , \latches_out_f[1][DATA][13] , 
        \latches_out_f[1][DATA][12] , \latches_out_f[1][DATA][11] , 
        \latches_out_f[1][DATA][10] , \latches_out_f[1][DATA][9] , 
        \latches_out_f[1][DATA][8] , \latches_out_f[1][DATA][7] , 
        \latches_out_f[1][DATA][6] , \latches_out_f[1][DATA][5] , 
        \latches_out_f[1][DATA][4] , \latches_out_f[1][DATA][3] , 
        \latches_out_f[1][DATA][2] , \latches_out_f[1][DATA][1] , 
        \latches_out_f[1][DATA][0] , \latches_out_f[0][REQ] , 
        \latches_out_f[0][DATA][34] , \latches_out_f[0][DATA][33] , 
        \latches_out_f[0][DATA][32] , \latches_out_f[0][DATA][31] , 
        \latches_out_f[0][DATA][30] , \latches_out_f[0][DATA][29] , 
        \latches_out_f[0][DATA][28] , \latches_out_f[0][DATA][27] , 
        \latches_out_f[0][DATA][26] , \latches_out_f[0][DATA][25] , 
        \latches_out_f[0][DATA][24] , \latches_out_f[0][DATA][23] , 
        \latches_out_f[0][DATA][22] , \latches_out_f[0][DATA][21] , 
        \latches_out_f[0][DATA][20] , \latches_out_f[0][DATA][19] , 
        \latches_out_f[0][DATA][18] , \latches_out_f[0][DATA][17] , 
        \latches_out_f[0][DATA][16] , \latches_out_f[0][DATA][15] , 
        \latches_out_f[0][DATA][14] , \latches_out_f[0][DATA][13] , 
        \latches_out_f[0][DATA][12] , \latches_out_f[0][DATA][11] , 
        \latches_out_f[0][DATA][10] , \latches_out_f[0][DATA][9] , 
        \latches_out_f[0][DATA][8] , \latches_out_f[0][DATA][7] , 
        \latches_out_f[0][DATA][6] , \latches_out_f[0][DATA][5] , 
        \latches_out_f[0][DATA][4] , \latches_out_f[0][DATA][3] , 
        \latches_out_f[0][DATA][2] , \latches_out_f[0][DATA][1] , 
        \latches_out_f[0][DATA][0] }), .latches_out_b({\latches_out_b[4][ACK] , 
        \latches_out_b[3][ACK] , \latches_out_b[2][ACK] , 
        \latches_out_b[1][ACK] , \latches_out_b[0][ACK] }) );
  input preset, \switch_sel[4][4] , \switch_sel[4][3] , \switch_sel[4][2] ,
         \switch_sel[4][1] , \switch_sel[4][0] , \switch_sel[3][4] ,
         \switch_sel[3][3] , \switch_sel[3][2] , \switch_sel[3][1] ,
         \switch_sel[3][0] , \switch_sel[2][4] , \switch_sel[2][3] ,
         \switch_sel[2][2] , \switch_sel[2][1] , \switch_sel[2][0] ,
         \switch_sel[1][4] , \switch_sel[1][3] , \switch_sel[1][2] ,
         \switch_sel[1][1] , \switch_sel[1][0] , \switch_sel[0][4] ,
         \switch_sel[0][3] , \switch_sel[0][2] , \switch_sel[0][1] ,
         \switch_sel[0][0] , \chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] ,
         \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] ,
         \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] ,
         \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] ,
         \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] ,
         \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] ,
         \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] ,
         \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] ,
         \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] ,
         \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] ,
         \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] ,
         \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] ,
         \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] ,
         \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] ,
         \chs_in_f[4][DATA][7] , \chs_in_f[4][DATA][6] ,
         \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] ,
         \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] ,
         \chs_in_f[4][DATA][1] , \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] ,
         \chs_in_f[3][DATA][34] , \chs_in_f[3][DATA][33] ,
         \chs_in_f[3][DATA][32] , \chs_in_f[3][DATA][31] ,
         \chs_in_f[3][DATA][30] , \chs_in_f[3][DATA][29] ,
         \chs_in_f[3][DATA][28] , \chs_in_f[3][DATA][27] ,
         \chs_in_f[3][DATA][26] , \chs_in_f[3][DATA][25] ,
         \chs_in_f[3][DATA][24] , \chs_in_f[3][DATA][23] ,
         \chs_in_f[3][DATA][22] , \chs_in_f[3][DATA][21] ,
         \chs_in_f[3][DATA][20] , \chs_in_f[3][DATA][19] ,
         \chs_in_f[3][DATA][18] , \chs_in_f[3][DATA][17] ,
         \chs_in_f[3][DATA][16] , \chs_in_f[3][DATA][15] ,
         \chs_in_f[3][DATA][14] , \chs_in_f[3][DATA][13] ,
         \chs_in_f[3][DATA][12] , \chs_in_f[3][DATA][11] ,
         \chs_in_f[3][DATA][10] , \chs_in_f[3][DATA][9] ,
         \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] ,
         \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] ,
         \chs_in_f[3][DATA][4] , \chs_in_f[3][DATA][3] ,
         \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] ,
         \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] ,
         \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] ,
         \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] ,
         \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] ,
         \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] ,
         \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] ,
         \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] ,
         \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] ,
         \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] ,
         \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] ,
         \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] ,
         \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] ,
         \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] ,
         \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] ,
         \chs_in_f[2][DATA][7] , \chs_in_f[2][DATA][6] ,
         \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] ,
         \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] ,
         \chs_in_f[2][DATA][1] , \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] ,
         \chs_in_f[1][DATA][34] , \chs_in_f[1][DATA][33] ,
         \chs_in_f[1][DATA][32] , \chs_in_f[1][DATA][31] ,
         \chs_in_f[1][DATA][30] , \chs_in_f[1][DATA][29] ,
         \chs_in_f[1][DATA][28] , \chs_in_f[1][DATA][27] ,
         \chs_in_f[1][DATA][26] , \chs_in_f[1][DATA][25] ,
         \chs_in_f[1][DATA][24] , \chs_in_f[1][DATA][23] ,
         \chs_in_f[1][DATA][22] , \chs_in_f[1][DATA][21] ,
         \chs_in_f[1][DATA][20] , \chs_in_f[1][DATA][19] ,
         \chs_in_f[1][DATA][18] , \chs_in_f[1][DATA][17] ,
         \chs_in_f[1][DATA][16] , \chs_in_f[1][DATA][15] ,
         \chs_in_f[1][DATA][14] , \chs_in_f[1][DATA][13] ,
         \chs_in_f[1][DATA][12] , \chs_in_f[1][DATA][11] ,
         \chs_in_f[1][DATA][10] , \chs_in_f[1][DATA][9] ,
         \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] ,
         \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] ,
         \chs_in_f[1][DATA][4] , \chs_in_f[1][DATA][3] ,
         \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] ,
         \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] ,
         \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] ,
         \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] ,
         \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] ,
         \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] ,
         \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] ,
         \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] ,
         \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] ,
         \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] ,
         \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] ,
         \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] ,
         \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] ,
         \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] ,
         \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] ,
         \chs_in_f[0][DATA][7] , \chs_in_f[0][DATA][6] ,
         \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] ,
         \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] ,
         \chs_in_f[0][DATA][1] , \chs_in_f[0][DATA][0] ,
         \latches_out_b[4][ACK] , \latches_out_b[3][ACK] ,
         \latches_out_b[2][ACK] , \latches_out_b[1][ACK] ,
         \latches_out_b[0][ACK] ;
  output \chs_in_b[4][ACK] , \chs_in_b[3][ACK] , \chs_in_b[2][ACK] ,
         \chs_in_b[1][ACK] , \chs_in_b[0][ACK] , \latches_out_f[4][REQ] ,
         \latches_out_f[4][DATA][34] , \latches_out_f[4][DATA][33] ,
         \latches_out_f[4][DATA][32] , \latches_out_f[4][DATA][31] ,
         \latches_out_f[4][DATA][30] , \latches_out_f[4][DATA][29] ,
         \latches_out_f[4][DATA][28] , \latches_out_f[4][DATA][27] ,
         \latches_out_f[4][DATA][26] , \latches_out_f[4][DATA][25] ,
         \latches_out_f[4][DATA][24] , \latches_out_f[4][DATA][23] ,
         \latches_out_f[4][DATA][22] , \latches_out_f[4][DATA][21] ,
         \latches_out_f[4][DATA][20] , \latches_out_f[4][DATA][19] ,
         \latches_out_f[4][DATA][18] , \latches_out_f[4][DATA][17] ,
         \latches_out_f[4][DATA][16] , \latches_out_f[4][DATA][15] ,
         \latches_out_f[4][DATA][14] , \latches_out_f[4][DATA][13] ,
         \latches_out_f[4][DATA][12] , \latches_out_f[4][DATA][11] ,
         \latches_out_f[4][DATA][10] , \latches_out_f[4][DATA][9] ,
         \latches_out_f[4][DATA][8] , \latches_out_f[4][DATA][7] ,
         \latches_out_f[4][DATA][6] , \latches_out_f[4][DATA][5] ,
         \latches_out_f[4][DATA][4] , \latches_out_f[4][DATA][3] ,
         \latches_out_f[4][DATA][2] , \latches_out_f[4][DATA][1] ,
         \latches_out_f[4][DATA][0] , \latches_out_f[3][REQ] ,
         \latches_out_f[3][DATA][34] , \latches_out_f[3][DATA][33] ,
         \latches_out_f[3][DATA][32] , \latches_out_f[3][DATA][31] ,
         \latches_out_f[3][DATA][30] , \latches_out_f[3][DATA][29] ,
         \latches_out_f[3][DATA][28] , \latches_out_f[3][DATA][27] ,
         \latches_out_f[3][DATA][26] , \latches_out_f[3][DATA][25] ,
         \latches_out_f[3][DATA][24] , \latches_out_f[3][DATA][23] ,
         \latches_out_f[3][DATA][22] , \latches_out_f[3][DATA][21] ,
         \latches_out_f[3][DATA][20] , \latches_out_f[3][DATA][19] ,
         \latches_out_f[3][DATA][18] , \latches_out_f[3][DATA][17] ,
         \latches_out_f[3][DATA][16] , \latches_out_f[3][DATA][15] ,
         \latches_out_f[3][DATA][14] , \latches_out_f[3][DATA][13] ,
         \latches_out_f[3][DATA][12] , \latches_out_f[3][DATA][11] ,
         \latches_out_f[3][DATA][10] , \latches_out_f[3][DATA][9] ,
         \latches_out_f[3][DATA][8] , \latches_out_f[3][DATA][7] ,
         \latches_out_f[3][DATA][6] , \latches_out_f[3][DATA][5] ,
         \latches_out_f[3][DATA][4] , \latches_out_f[3][DATA][3] ,
         \latches_out_f[3][DATA][2] , \latches_out_f[3][DATA][1] ,
         \latches_out_f[3][DATA][0] , \latches_out_f[2][REQ] ,
         \latches_out_f[2][DATA][34] , \latches_out_f[2][DATA][33] ,
         \latches_out_f[2][DATA][32] , \latches_out_f[2][DATA][31] ,
         \latches_out_f[2][DATA][30] , \latches_out_f[2][DATA][29] ,
         \latches_out_f[2][DATA][28] , \latches_out_f[2][DATA][27] ,
         \latches_out_f[2][DATA][26] , \latches_out_f[2][DATA][25] ,
         \latches_out_f[2][DATA][24] , \latches_out_f[2][DATA][23] ,
         \latches_out_f[2][DATA][22] , \latches_out_f[2][DATA][21] ,
         \latches_out_f[2][DATA][20] , \latches_out_f[2][DATA][19] ,
         \latches_out_f[2][DATA][18] , \latches_out_f[2][DATA][17] ,
         \latches_out_f[2][DATA][16] , \latches_out_f[2][DATA][15] ,
         \latches_out_f[2][DATA][14] , \latches_out_f[2][DATA][13] ,
         \latches_out_f[2][DATA][12] , \latches_out_f[2][DATA][11] ,
         \latches_out_f[2][DATA][10] , \latches_out_f[2][DATA][9] ,
         \latches_out_f[2][DATA][8] , \latches_out_f[2][DATA][7] ,
         \latches_out_f[2][DATA][6] , \latches_out_f[2][DATA][5] ,
         \latches_out_f[2][DATA][4] , \latches_out_f[2][DATA][3] ,
         \latches_out_f[2][DATA][2] , \latches_out_f[2][DATA][1] ,
         \latches_out_f[2][DATA][0] , \latches_out_f[1][REQ] ,
         \latches_out_f[1][DATA][34] , \latches_out_f[1][DATA][33] ,
         \latches_out_f[1][DATA][32] , \latches_out_f[1][DATA][31] ,
         \latches_out_f[1][DATA][30] , \latches_out_f[1][DATA][29] ,
         \latches_out_f[1][DATA][28] , \latches_out_f[1][DATA][27] ,
         \latches_out_f[1][DATA][26] , \latches_out_f[1][DATA][25] ,
         \latches_out_f[1][DATA][24] , \latches_out_f[1][DATA][23] ,
         \latches_out_f[1][DATA][22] , \latches_out_f[1][DATA][21] ,
         \latches_out_f[1][DATA][20] , \latches_out_f[1][DATA][19] ,
         \latches_out_f[1][DATA][18] , \latches_out_f[1][DATA][17] ,
         \latches_out_f[1][DATA][16] , \latches_out_f[1][DATA][15] ,
         \latches_out_f[1][DATA][14] , \latches_out_f[1][DATA][13] ,
         \latches_out_f[1][DATA][12] , \latches_out_f[1][DATA][11] ,
         \latches_out_f[1][DATA][10] , \latches_out_f[1][DATA][9] ,
         \latches_out_f[1][DATA][8] , \latches_out_f[1][DATA][7] ,
         \latches_out_f[1][DATA][6] , \latches_out_f[1][DATA][5] ,
         \latches_out_f[1][DATA][4] , \latches_out_f[1][DATA][3] ,
         \latches_out_f[1][DATA][2] , \latches_out_f[1][DATA][1] ,
         \latches_out_f[1][DATA][0] , \latches_out_f[0][REQ] ,
         \latches_out_f[0][DATA][34] , \latches_out_f[0][DATA][33] ,
         \latches_out_f[0][DATA][32] , \latches_out_f[0][DATA][31] ,
         \latches_out_f[0][DATA][30] , \latches_out_f[0][DATA][29] ,
         \latches_out_f[0][DATA][28] , \latches_out_f[0][DATA][27] ,
         \latches_out_f[0][DATA][26] , \latches_out_f[0][DATA][25] ,
         \latches_out_f[0][DATA][24] , \latches_out_f[0][DATA][23] ,
         \latches_out_f[0][DATA][22] , \latches_out_f[0][DATA][21] ,
         \latches_out_f[0][DATA][20] , \latches_out_f[0][DATA][19] ,
         \latches_out_f[0][DATA][18] , \latches_out_f[0][DATA][17] ,
         \latches_out_f[0][DATA][16] , \latches_out_f[0][DATA][15] ,
         \latches_out_f[0][DATA][14] , \latches_out_f[0][DATA][13] ,
         \latches_out_f[0][DATA][12] , \latches_out_f[0][DATA][11] ,
         \latches_out_f[0][DATA][10] , \latches_out_f[0][DATA][9] ,
         \latches_out_f[0][DATA][8] , \latches_out_f[0][DATA][7] ,
         \latches_out_f[0][DATA][6] , \latches_out_f[0][DATA][5] ,
         \latches_out_f[0][DATA][4] , \latches_out_f[0][DATA][3] ,
         \latches_out_f[0][DATA][2] , \latches_out_f[0][DATA][1] ,
         \latches_out_f[0][DATA][0] ;
  wire   \latches_in_f[4][REQ] , \latches_in_f[4][DATA][34] ,
         \latches_in_f[4][DATA][33] , \latches_in_f[4][DATA][32] ,
         \latches_in_f[4][DATA][31] , \latches_in_f[4][DATA][30] ,
         \latches_in_f[4][DATA][29] , \latches_in_f[4][DATA][28] ,
         \latches_in_f[4][DATA][27] , \latches_in_f[4][DATA][26] ,
         \latches_in_f[4][DATA][25] , \latches_in_f[4][DATA][24] ,
         \latches_in_f[4][DATA][23] , \latches_in_f[4][DATA][22] ,
         \latches_in_f[4][DATA][21] , \latches_in_f[4][DATA][20] ,
         \latches_in_f[4][DATA][19] , \latches_in_f[4][DATA][18] ,
         \latches_in_f[4][DATA][17] , \latches_in_f[4][DATA][16] ,
         \latches_in_f[4][DATA][15] , \latches_in_f[4][DATA][14] ,
         \latches_in_f[4][DATA][13] , \latches_in_f[4][DATA][12] ,
         \latches_in_f[4][DATA][11] , \latches_in_f[4][DATA][10] ,
         \latches_in_f[4][DATA][9] , \latches_in_f[4][DATA][8] ,
         \latches_in_f[4][DATA][7] , \latches_in_f[4][DATA][6] ,
         \latches_in_f[4][DATA][5] , \latches_in_f[4][DATA][4] ,
         \latches_in_f[4][DATA][3] , \latches_in_f[4][DATA][2] ,
         \latches_in_f[4][DATA][1] , \latches_in_f[4][DATA][0] ,
         \latches_in_f[3][REQ] , \latches_in_f[3][DATA][34] ,
         \latches_in_f[3][DATA][33] , \latches_in_f[3][DATA][32] ,
         \latches_in_f[3][DATA][31] , \latches_in_f[3][DATA][30] ,
         \latches_in_f[3][DATA][29] , \latches_in_f[3][DATA][28] ,
         \latches_in_f[3][DATA][27] , \latches_in_f[3][DATA][26] ,
         \latches_in_f[3][DATA][25] , \latches_in_f[3][DATA][24] ,
         \latches_in_f[3][DATA][23] , \latches_in_f[3][DATA][22] ,
         \latches_in_f[3][DATA][21] , \latches_in_f[3][DATA][20] ,
         \latches_in_f[3][DATA][19] , \latches_in_f[3][DATA][18] ,
         \latches_in_f[3][DATA][17] , \latches_in_f[3][DATA][16] ,
         \latches_in_f[3][DATA][15] , \latches_in_f[3][DATA][14] ,
         \latches_in_f[3][DATA][13] , \latches_in_f[3][DATA][12] ,
         \latches_in_f[3][DATA][11] , \latches_in_f[3][DATA][10] ,
         \latches_in_f[3][DATA][9] , \latches_in_f[3][DATA][8] ,
         \latches_in_f[3][DATA][7] , \latches_in_f[3][DATA][6] ,
         \latches_in_f[3][DATA][5] , \latches_in_f[3][DATA][4] ,
         \latches_in_f[3][DATA][3] , \latches_in_f[3][DATA][2] ,
         \latches_in_f[3][DATA][1] , \latches_in_f[3][DATA][0] ,
         \latches_in_f[2][REQ] , \latches_in_f[2][DATA][34] ,
         \latches_in_f[2][DATA][33] , \latches_in_f[2][DATA][32] ,
         \latches_in_f[2][DATA][31] , \latches_in_f[2][DATA][30] ,
         \latches_in_f[2][DATA][29] , \latches_in_f[2][DATA][28] ,
         \latches_in_f[2][DATA][27] , \latches_in_f[2][DATA][26] ,
         \latches_in_f[2][DATA][25] , \latches_in_f[2][DATA][24] ,
         \latches_in_f[2][DATA][23] , \latches_in_f[2][DATA][22] ,
         \latches_in_f[2][DATA][21] , \latches_in_f[2][DATA][20] ,
         \latches_in_f[2][DATA][19] , \latches_in_f[2][DATA][18] ,
         \latches_in_f[2][DATA][17] , \latches_in_f[2][DATA][16] ,
         \latches_in_f[2][DATA][15] , \latches_in_f[2][DATA][14] ,
         \latches_in_f[2][DATA][13] , \latches_in_f[2][DATA][12] ,
         \latches_in_f[2][DATA][11] , \latches_in_f[2][DATA][10] ,
         \latches_in_f[2][DATA][9] , \latches_in_f[2][DATA][8] ,
         \latches_in_f[2][DATA][7] , \latches_in_f[2][DATA][6] ,
         \latches_in_f[2][DATA][5] , \latches_in_f[2][DATA][4] ,
         \latches_in_f[2][DATA][3] , \latches_in_f[2][DATA][2] ,
         \latches_in_f[2][DATA][1] , \latches_in_f[2][DATA][0] ,
         \latches_in_f[1][REQ] , \latches_in_f[1][DATA][34] ,
         \latches_in_f[1][DATA][33] , \latches_in_f[1][DATA][32] ,
         \latches_in_f[1][DATA][31] , \latches_in_f[1][DATA][30] ,
         \latches_in_f[1][DATA][29] , \latches_in_f[1][DATA][28] ,
         \latches_in_f[1][DATA][27] , \latches_in_f[1][DATA][26] ,
         \latches_in_f[1][DATA][25] , \latches_in_f[1][DATA][24] ,
         \latches_in_f[1][DATA][23] , \latches_in_f[1][DATA][22] ,
         \latches_in_f[1][DATA][21] , \latches_in_f[1][DATA][20] ,
         \latches_in_f[1][DATA][19] , \latches_in_f[1][DATA][18] ,
         \latches_in_f[1][DATA][17] , \latches_in_f[1][DATA][16] ,
         \latches_in_f[1][DATA][15] , \latches_in_f[1][DATA][14] ,
         \latches_in_f[1][DATA][13] , \latches_in_f[1][DATA][12] ,
         \latches_in_f[1][DATA][11] , \latches_in_f[1][DATA][10] ,
         \latches_in_f[1][DATA][9] , \latches_in_f[1][DATA][8] ,
         \latches_in_f[1][DATA][7] , \latches_in_f[1][DATA][6] ,
         \latches_in_f[1][DATA][5] , \latches_in_f[1][DATA][4] ,
         \latches_in_f[1][DATA][3] , \latches_in_f[1][DATA][2] ,
         \latches_in_f[1][DATA][1] , \latches_in_f[1][DATA][0] ,
         \latches_in_f[0][REQ] , \latches_in_f[0][DATA][34] ,
         \latches_in_f[0][DATA][33] , \latches_in_f[0][DATA][32] ,
         \latches_in_f[0][DATA][31] , \latches_in_f[0][DATA][30] ,
         \latches_in_f[0][DATA][29] , \latches_in_f[0][DATA][28] ,
         \latches_in_f[0][DATA][27] , \latches_in_f[0][DATA][26] ,
         \latches_in_f[0][DATA][25] , \latches_in_f[0][DATA][24] ,
         \latches_in_f[0][DATA][23] , \latches_in_f[0][DATA][22] ,
         \latches_in_f[0][DATA][21] , \latches_in_f[0][DATA][20] ,
         \latches_in_f[0][DATA][19] , \latches_in_f[0][DATA][18] ,
         \latches_in_f[0][DATA][17] , \latches_in_f[0][DATA][16] ,
         \latches_in_f[0][DATA][15] , \latches_in_f[0][DATA][14] ,
         \latches_in_f[0][DATA][13] , \latches_in_f[0][DATA][12] ,
         \latches_in_f[0][DATA][11] , \latches_in_f[0][DATA][10] ,
         \latches_in_f[0][DATA][9] , \latches_in_f[0][DATA][8] ,
         \latches_in_f[0][DATA][7] , \latches_in_f[0][DATA][6] ,
         \latches_in_f[0][DATA][5] , \latches_in_f[0][DATA][4] ,
         \latches_in_f[0][DATA][3] , \latches_in_f[0][DATA][2] ,
         \latches_in_f[0][DATA][1] , \latches_in_f[0][DATA][0] ,
         \latches_in_b[4][ACK] , \latches_in_b[3][ACK] ,
         \latches_in_b[2][ACK] , \latches_in_b[1][ACK] ,
         \latches_in_b[0][ACK] , n1;

  crossbar_1 crossbar ( .preset(n1), .switch_sel({\switch_sel[4][4] , 
        \switch_sel[4][3] , \switch_sel[4][2] , \switch_sel[4][1] , 
        \switch_sel[4][0] , \switch_sel[3][4] , \switch_sel[3][3] , 
        \switch_sel[3][2] , \switch_sel[3][1] , \switch_sel[3][0] , 
        \switch_sel[2][4] , \switch_sel[2][3] , \switch_sel[2][2] , 
        \switch_sel[2][1] , \switch_sel[2][0] , \switch_sel[1][4] , 
        \switch_sel[1][3] , \switch_sel[1][2] , \switch_sel[1][1] , 
        \switch_sel[1][0] , \switch_sel[0][4] , \switch_sel[0][3] , 
        \switch_sel[0][2] , \switch_sel[0][1] , \switch_sel[0][0] }), 
        .chs_in_f({\chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] , 
        \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] , 
        \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] , 
        \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] , 
        \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] , 
        \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] , 
        \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] , 
        \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] , 
        \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] , 
        \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] , 
        \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] , 
        \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] , 
        \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] , 
        \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] , \chs_in_f[4][DATA][7] , 
        \chs_in_f[4][DATA][6] , \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] , 
        \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] , \chs_in_f[4][DATA][1] , 
        \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] , \chs_in_f[3][DATA][34] , 
        \chs_in_f[3][DATA][33] , \chs_in_f[3][DATA][32] , 
        \chs_in_f[3][DATA][31] , \chs_in_f[3][DATA][30] , 
        \chs_in_f[3][DATA][29] , \chs_in_f[3][DATA][28] , 
        \chs_in_f[3][DATA][27] , \chs_in_f[3][DATA][26] , 
        \chs_in_f[3][DATA][25] , \chs_in_f[3][DATA][24] , 
        \chs_in_f[3][DATA][23] , \chs_in_f[3][DATA][22] , 
        \chs_in_f[3][DATA][21] , \chs_in_f[3][DATA][20] , 
        \chs_in_f[3][DATA][19] , \chs_in_f[3][DATA][18] , 
        \chs_in_f[3][DATA][17] , \chs_in_f[3][DATA][16] , 
        \chs_in_f[3][DATA][15] , \chs_in_f[3][DATA][14] , 
        \chs_in_f[3][DATA][13] , \chs_in_f[3][DATA][12] , 
        \chs_in_f[3][DATA][11] , \chs_in_f[3][DATA][10] , 
        \chs_in_f[3][DATA][9] , \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] , 
        \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] , \chs_in_f[3][DATA][4] , 
        \chs_in_f[3][DATA][3] , \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] , 
        \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] , 
        \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] , 
        \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] , 
        \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] , 
        \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] , 
        \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] , 
        \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] , 
        \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] , 
        \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] , 
        \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] , 
        \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] , 
        \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] , 
        \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] , 
        \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] , \chs_in_f[2][DATA][7] , 
        \chs_in_f[2][DATA][6] , \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] , 
        \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] , \chs_in_f[2][DATA][1] , 
        \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] , \chs_in_f[1][DATA][34] , 
        \chs_in_f[1][DATA][33] , \chs_in_f[1][DATA][32] , 
        \chs_in_f[1][DATA][31] , \chs_in_f[1][DATA][30] , 
        \chs_in_f[1][DATA][29] , \chs_in_f[1][DATA][28] , 
        \chs_in_f[1][DATA][27] , \chs_in_f[1][DATA][26] , 
        \chs_in_f[1][DATA][25] , \chs_in_f[1][DATA][24] , 
        \chs_in_f[1][DATA][23] , \chs_in_f[1][DATA][22] , 
        \chs_in_f[1][DATA][21] , \chs_in_f[1][DATA][20] , 
        \chs_in_f[1][DATA][19] , \chs_in_f[1][DATA][18] , 
        \chs_in_f[1][DATA][17] , \chs_in_f[1][DATA][16] , 
        \chs_in_f[1][DATA][15] , \chs_in_f[1][DATA][14] , 
        \chs_in_f[1][DATA][13] , \chs_in_f[1][DATA][12] , 
        \chs_in_f[1][DATA][11] , \chs_in_f[1][DATA][10] , 
        \chs_in_f[1][DATA][9] , \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] , 
        \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] , \chs_in_f[1][DATA][4] , 
        \chs_in_f[1][DATA][3] , \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] , 
        \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] , 
        \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] , 
        \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] , 
        \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] , 
        \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] , 
        \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] , 
        \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] , 
        \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] , 
        \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] , 
        \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] , 
        \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] , 
        \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] , 
        \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] , 
        \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] , \chs_in_f[0][DATA][7] , 
        \chs_in_f[0][DATA][6] , \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] , 
        \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] , \chs_in_f[0][DATA][1] , 
        \chs_in_f[0][DATA][0] }), .chs_in_b({\chs_in_b[4][ACK] , 
        \chs_in_b[3][ACK] , \chs_in_b[2][ACK] , \chs_in_b[1][ACK] , 
        \chs_in_b[0][ACK] }), .chs_out_f({\latches_in_f[4][REQ] , 
        \latches_in_f[4][DATA][34] , \latches_in_f[4][DATA][33] , 
        \latches_in_f[4][DATA][32] , \latches_in_f[4][DATA][31] , 
        \latches_in_f[4][DATA][30] , \latches_in_f[4][DATA][29] , 
        \latches_in_f[4][DATA][28] , \latches_in_f[4][DATA][27] , 
        \latches_in_f[4][DATA][26] , \latches_in_f[4][DATA][25] , 
        \latches_in_f[4][DATA][24] , \latches_in_f[4][DATA][23] , 
        \latches_in_f[4][DATA][22] , \latches_in_f[4][DATA][21] , 
        \latches_in_f[4][DATA][20] , \latches_in_f[4][DATA][19] , 
        \latches_in_f[4][DATA][18] , \latches_in_f[4][DATA][17] , 
        \latches_in_f[4][DATA][16] , \latches_in_f[4][DATA][15] , 
        \latches_in_f[4][DATA][14] , \latches_in_f[4][DATA][13] , 
        \latches_in_f[4][DATA][12] , \latches_in_f[4][DATA][11] , 
        \latches_in_f[4][DATA][10] , \latches_in_f[4][DATA][9] , 
        \latches_in_f[4][DATA][8] , \latches_in_f[4][DATA][7] , 
        \latches_in_f[4][DATA][6] , \latches_in_f[4][DATA][5] , 
        \latches_in_f[4][DATA][4] , \latches_in_f[4][DATA][3] , 
        \latches_in_f[4][DATA][2] , \latches_in_f[4][DATA][1] , 
        \latches_in_f[4][DATA][0] , \latches_in_f[3][REQ] , 
        \latches_in_f[3][DATA][34] , \latches_in_f[3][DATA][33] , 
        \latches_in_f[3][DATA][32] , \latches_in_f[3][DATA][31] , 
        \latches_in_f[3][DATA][30] , \latches_in_f[3][DATA][29] , 
        \latches_in_f[3][DATA][28] , \latches_in_f[3][DATA][27] , 
        \latches_in_f[3][DATA][26] , \latches_in_f[3][DATA][25] , 
        \latches_in_f[3][DATA][24] , \latches_in_f[3][DATA][23] , 
        \latches_in_f[3][DATA][22] , \latches_in_f[3][DATA][21] , 
        \latches_in_f[3][DATA][20] , \latches_in_f[3][DATA][19] , 
        \latches_in_f[3][DATA][18] , \latches_in_f[3][DATA][17] , 
        \latches_in_f[3][DATA][16] , \latches_in_f[3][DATA][15] , 
        \latches_in_f[3][DATA][14] , \latches_in_f[3][DATA][13] , 
        \latches_in_f[3][DATA][12] , \latches_in_f[3][DATA][11] , 
        \latches_in_f[3][DATA][10] , \latches_in_f[3][DATA][9] , 
        \latches_in_f[3][DATA][8] , \latches_in_f[3][DATA][7] , 
        \latches_in_f[3][DATA][6] , \latches_in_f[3][DATA][5] , 
        \latches_in_f[3][DATA][4] , \latches_in_f[3][DATA][3] , 
        \latches_in_f[3][DATA][2] , \latches_in_f[3][DATA][1] , 
        \latches_in_f[3][DATA][0] , \latches_in_f[2][REQ] , 
        \latches_in_f[2][DATA][34] , \latches_in_f[2][DATA][33] , 
        \latches_in_f[2][DATA][32] , \latches_in_f[2][DATA][31] , 
        \latches_in_f[2][DATA][30] , \latches_in_f[2][DATA][29] , 
        \latches_in_f[2][DATA][28] , \latches_in_f[2][DATA][27] , 
        \latches_in_f[2][DATA][26] , \latches_in_f[2][DATA][25] , 
        \latches_in_f[2][DATA][24] , \latches_in_f[2][DATA][23] , 
        \latches_in_f[2][DATA][22] , \latches_in_f[2][DATA][21] , 
        \latches_in_f[2][DATA][20] , \latches_in_f[2][DATA][19] , 
        \latches_in_f[2][DATA][18] , \latches_in_f[2][DATA][17] , 
        \latches_in_f[2][DATA][16] , \latches_in_f[2][DATA][15] , 
        \latches_in_f[2][DATA][14] , \latches_in_f[2][DATA][13] , 
        \latches_in_f[2][DATA][12] , \latches_in_f[2][DATA][11] , 
        \latches_in_f[2][DATA][10] , \latches_in_f[2][DATA][9] , 
        \latches_in_f[2][DATA][8] , \latches_in_f[2][DATA][7] , 
        \latches_in_f[2][DATA][6] , \latches_in_f[2][DATA][5] , 
        \latches_in_f[2][DATA][4] , \latches_in_f[2][DATA][3] , 
        \latches_in_f[2][DATA][2] , \latches_in_f[2][DATA][1] , 
        \latches_in_f[2][DATA][0] , \latches_in_f[1][REQ] , 
        \latches_in_f[1][DATA][34] , \latches_in_f[1][DATA][33] , 
        \latches_in_f[1][DATA][32] , \latches_in_f[1][DATA][31] , 
        \latches_in_f[1][DATA][30] , \latches_in_f[1][DATA][29] , 
        \latches_in_f[1][DATA][28] , \latches_in_f[1][DATA][27] , 
        \latches_in_f[1][DATA][26] , \latches_in_f[1][DATA][25] , 
        \latches_in_f[1][DATA][24] , \latches_in_f[1][DATA][23] , 
        \latches_in_f[1][DATA][22] , \latches_in_f[1][DATA][21] , 
        \latches_in_f[1][DATA][20] , \latches_in_f[1][DATA][19] , 
        \latches_in_f[1][DATA][18] , \latches_in_f[1][DATA][17] , 
        \latches_in_f[1][DATA][16] , \latches_in_f[1][DATA][15] , 
        \latches_in_f[1][DATA][14] , \latches_in_f[1][DATA][13] , 
        \latches_in_f[1][DATA][12] , \latches_in_f[1][DATA][11] , 
        \latches_in_f[1][DATA][10] , \latches_in_f[1][DATA][9] , 
        \latches_in_f[1][DATA][8] , \latches_in_f[1][DATA][7] , 
        \latches_in_f[1][DATA][6] , \latches_in_f[1][DATA][5] , 
        \latches_in_f[1][DATA][4] , \latches_in_f[1][DATA][3] , 
        \latches_in_f[1][DATA][2] , \latches_in_f[1][DATA][1] , 
        \latches_in_f[1][DATA][0] , \latches_in_f[0][REQ] , 
        \latches_in_f[0][DATA][34] , \latches_in_f[0][DATA][33] , 
        \latches_in_f[0][DATA][32] , \latches_in_f[0][DATA][31] , 
        \latches_in_f[0][DATA][30] , \latches_in_f[0][DATA][29] , 
        \latches_in_f[0][DATA][28] , \latches_in_f[0][DATA][27] , 
        \latches_in_f[0][DATA][26] , \latches_in_f[0][DATA][25] , 
        \latches_in_f[0][DATA][24] , \latches_in_f[0][DATA][23] , 
        \latches_in_f[0][DATA][22] , \latches_in_f[0][DATA][21] , 
        \latches_in_f[0][DATA][20] , \latches_in_f[0][DATA][19] , 
        \latches_in_f[0][DATA][18] , \latches_in_f[0][DATA][17] , 
        \latches_in_f[0][DATA][16] , \latches_in_f[0][DATA][15] , 
        \latches_in_f[0][DATA][14] , \latches_in_f[0][DATA][13] , 
        \latches_in_f[0][DATA][12] , \latches_in_f[0][DATA][11] , 
        \latches_in_f[0][DATA][10] , \latches_in_f[0][DATA][9] , 
        \latches_in_f[0][DATA][8] , \latches_in_f[0][DATA][7] , 
        \latches_in_f[0][DATA][6] , \latches_in_f[0][DATA][5] , 
        \latches_in_f[0][DATA][4] , \latches_in_f[0][DATA][3] , 
        \latches_in_f[0][DATA][2] , \latches_in_f[0][DATA][1] , 
        \latches_in_f[0][DATA][0] }), .chs_out_b({\latches_in_b[4][ACK] , 
        \latches_in_b[3][ACK] , \latches_in_b[2][ACK] , \latches_in_b[1][ACK] , 
        \latches_in_b[0][ACK] }) );
  channel_latch_0_000000000_5 ch_latch_4 ( .preset(n1), .left_in({
        \latches_in_f[4][REQ] , \latches_in_f[4][DATA][34] , 
        \latches_in_f[4][DATA][33] , \latches_in_f[4][DATA][32] , 
        \latches_in_f[4][DATA][31] , \latches_in_f[4][DATA][30] , 
        \latches_in_f[4][DATA][29] , \latches_in_f[4][DATA][28] , 
        \latches_in_f[4][DATA][27] , \latches_in_f[4][DATA][26] , 
        \latches_in_f[4][DATA][25] , \latches_in_f[4][DATA][24] , 
        \latches_in_f[4][DATA][23] , \latches_in_f[4][DATA][22] , 
        \latches_in_f[4][DATA][21] , \latches_in_f[4][DATA][20] , 
        \latches_in_f[4][DATA][19] , \latches_in_f[4][DATA][18] , 
        \latches_in_f[4][DATA][17] , \latches_in_f[4][DATA][16] , 
        \latches_in_f[4][DATA][15] , \latches_in_f[4][DATA][14] , 
        \latches_in_f[4][DATA][13] , \latches_in_f[4][DATA][12] , 
        \latches_in_f[4][DATA][11] , \latches_in_f[4][DATA][10] , 
        \latches_in_f[4][DATA][9] , \latches_in_f[4][DATA][8] , 
        \latches_in_f[4][DATA][7] , \latches_in_f[4][DATA][6] , 
        \latches_in_f[4][DATA][5] , \latches_in_f[4][DATA][4] , 
        \latches_in_f[4][DATA][3] , \latches_in_f[4][DATA][2] , 
        \latches_in_f[4][DATA][1] , \latches_in_f[4][DATA][0] }), .left_out(
        \latches_in_b[4][ACK] ), .right_out({\latches_out_f[4][REQ] , 
        \latches_out_f[4][DATA][34] , \latches_out_f[4][DATA][33] , 
        \latches_out_f[4][DATA][32] , \latches_out_f[4][DATA][31] , 
        \latches_out_f[4][DATA][30] , \latches_out_f[4][DATA][29] , 
        \latches_out_f[4][DATA][28] , \latches_out_f[4][DATA][27] , 
        \latches_out_f[4][DATA][26] , \latches_out_f[4][DATA][25] , 
        \latches_out_f[4][DATA][24] , \latches_out_f[4][DATA][23] , 
        \latches_out_f[4][DATA][22] , \latches_out_f[4][DATA][21] , 
        \latches_out_f[4][DATA][20] , \latches_out_f[4][DATA][19] , 
        \latches_out_f[4][DATA][18] , \latches_out_f[4][DATA][17] , 
        \latches_out_f[4][DATA][16] , \latches_out_f[4][DATA][15] , 
        \latches_out_f[4][DATA][14] , \latches_out_f[4][DATA][13] , 
        \latches_out_f[4][DATA][12] , \latches_out_f[4][DATA][11] , 
        \latches_out_f[4][DATA][10] , \latches_out_f[4][DATA][9] , 
        \latches_out_f[4][DATA][8] , \latches_out_f[4][DATA][7] , 
        \latches_out_f[4][DATA][6] , \latches_out_f[4][DATA][5] , 
        \latches_out_f[4][DATA][4] , \latches_out_f[4][DATA][3] , 
        \latches_out_f[4][DATA][2] , \latches_out_f[4][DATA][1] , 
        \latches_out_f[4][DATA][0] }), .right_in(\latches_out_b[4][ACK] ) );
  channel_latch_0_000000000_4 ch_latch_3 ( .preset(n1), .left_in({
        \latches_in_f[3][REQ] , \latches_in_f[3][DATA][34] , 
        \latches_in_f[3][DATA][33] , \latches_in_f[3][DATA][32] , 
        \latches_in_f[3][DATA][31] , \latches_in_f[3][DATA][30] , 
        \latches_in_f[3][DATA][29] , \latches_in_f[3][DATA][28] , 
        \latches_in_f[3][DATA][27] , \latches_in_f[3][DATA][26] , 
        \latches_in_f[3][DATA][25] , \latches_in_f[3][DATA][24] , 
        \latches_in_f[3][DATA][23] , \latches_in_f[3][DATA][22] , 
        \latches_in_f[3][DATA][21] , \latches_in_f[3][DATA][20] , 
        \latches_in_f[3][DATA][19] , \latches_in_f[3][DATA][18] , 
        \latches_in_f[3][DATA][17] , \latches_in_f[3][DATA][16] , 
        \latches_in_f[3][DATA][15] , \latches_in_f[3][DATA][14] , 
        \latches_in_f[3][DATA][13] , \latches_in_f[3][DATA][12] , 
        \latches_in_f[3][DATA][11] , \latches_in_f[3][DATA][10] , 
        \latches_in_f[3][DATA][9] , \latches_in_f[3][DATA][8] , 
        \latches_in_f[3][DATA][7] , \latches_in_f[3][DATA][6] , 
        \latches_in_f[3][DATA][5] , \latches_in_f[3][DATA][4] , 
        \latches_in_f[3][DATA][3] , \latches_in_f[3][DATA][2] , 
        \latches_in_f[3][DATA][1] , \latches_in_f[3][DATA][0] }), .left_out(
        \latches_in_b[3][ACK] ), .right_out({\latches_out_f[3][REQ] , 
        \latches_out_f[3][DATA][34] , \latches_out_f[3][DATA][33] , 
        \latches_out_f[3][DATA][32] , \latches_out_f[3][DATA][31] , 
        \latches_out_f[3][DATA][30] , \latches_out_f[3][DATA][29] , 
        \latches_out_f[3][DATA][28] , \latches_out_f[3][DATA][27] , 
        \latches_out_f[3][DATA][26] , \latches_out_f[3][DATA][25] , 
        \latches_out_f[3][DATA][24] , \latches_out_f[3][DATA][23] , 
        \latches_out_f[3][DATA][22] , \latches_out_f[3][DATA][21] , 
        \latches_out_f[3][DATA][20] , \latches_out_f[3][DATA][19] , 
        \latches_out_f[3][DATA][18] , \latches_out_f[3][DATA][17] , 
        \latches_out_f[3][DATA][16] , \latches_out_f[3][DATA][15] , 
        \latches_out_f[3][DATA][14] , \latches_out_f[3][DATA][13] , 
        \latches_out_f[3][DATA][12] , \latches_out_f[3][DATA][11] , 
        \latches_out_f[3][DATA][10] , \latches_out_f[3][DATA][9] , 
        \latches_out_f[3][DATA][8] , \latches_out_f[3][DATA][7] , 
        \latches_out_f[3][DATA][6] , \latches_out_f[3][DATA][5] , 
        \latches_out_f[3][DATA][4] , \latches_out_f[3][DATA][3] , 
        \latches_out_f[3][DATA][2] , \latches_out_f[3][DATA][1] , 
        \latches_out_f[3][DATA][0] }), .right_in(\latches_out_b[3][ACK] ) );
  channel_latch_0_000000000_3 ch_latch_2 ( .preset(n1), .left_in({
        \latches_in_f[2][REQ] , \latches_in_f[2][DATA][34] , 
        \latches_in_f[2][DATA][33] , \latches_in_f[2][DATA][32] , 
        \latches_in_f[2][DATA][31] , \latches_in_f[2][DATA][30] , 
        \latches_in_f[2][DATA][29] , \latches_in_f[2][DATA][28] , 
        \latches_in_f[2][DATA][27] , \latches_in_f[2][DATA][26] , 
        \latches_in_f[2][DATA][25] , \latches_in_f[2][DATA][24] , 
        \latches_in_f[2][DATA][23] , \latches_in_f[2][DATA][22] , 
        \latches_in_f[2][DATA][21] , \latches_in_f[2][DATA][20] , 
        \latches_in_f[2][DATA][19] , \latches_in_f[2][DATA][18] , 
        \latches_in_f[2][DATA][17] , \latches_in_f[2][DATA][16] , 
        \latches_in_f[2][DATA][15] , \latches_in_f[2][DATA][14] , 
        \latches_in_f[2][DATA][13] , \latches_in_f[2][DATA][12] , 
        \latches_in_f[2][DATA][11] , \latches_in_f[2][DATA][10] , 
        \latches_in_f[2][DATA][9] , \latches_in_f[2][DATA][8] , 
        \latches_in_f[2][DATA][7] , \latches_in_f[2][DATA][6] , 
        \latches_in_f[2][DATA][5] , \latches_in_f[2][DATA][4] , 
        \latches_in_f[2][DATA][3] , \latches_in_f[2][DATA][2] , 
        \latches_in_f[2][DATA][1] , \latches_in_f[2][DATA][0] }), .left_out(
        \latches_in_b[2][ACK] ), .right_out({\latches_out_f[2][REQ] , 
        \latches_out_f[2][DATA][34] , \latches_out_f[2][DATA][33] , 
        \latches_out_f[2][DATA][32] , \latches_out_f[2][DATA][31] , 
        \latches_out_f[2][DATA][30] , \latches_out_f[2][DATA][29] , 
        \latches_out_f[2][DATA][28] , \latches_out_f[2][DATA][27] , 
        \latches_out_f[2][DATA][26] , \latches_out_f[2][DATA][25] , 
        \latches_out_f[2][DATA][24] , \latches_out_f[2][DATA][23] , 
        \latches_out_f[2][DATA][22] , \latches_out_f[2][DATA][21] , 
        \latches_out_f[2][DATA][20] , \latches_out_f[2][DATA][19] , 
        \latches_out_f[2][DATA][18] , \latches_out_f[2][DATA][17] , 
        \latches_out_f[2][DATA][16] , \latches_out_f[2][DATA][15] , 
        \latches_out_f[2][DATA][14] , \latches_out_f[2][DATA][13] , 
        \latches_out_f[2][DATA][12] , \latches_out_f[2][DATA][11] , 
        \latches_out_f[2][DATA][10] , \latches_out_f[2][DATA][9] , 
        \latches_out_f[2][DATA][8] , \latches_out_f[2][DATA][7] , 
        \latches_out_f[2][DATA][6] , \latches_out_f[2][DATA][5] , 
        \latches_out_f[2][DATA][4] , \latches_out_f[2][DATA][3] , 
        \latches_out_f[2][DATA][2] , \latches_out_f[2][DATA][1] , 
        \latches_out_f[2][DATA][0] }), .right_in(\latches_out_b[2][ACK] ) );
  channel_latch_0_000000000_2 ch_latch_1 ( .preset(n1), .left_in({
        \latches_in_f[1][REQ] , \latches_in_f[1][DATA][34] , 
        \latches_in_f[1][DATA][33] , \latches_in_f[1][DATA][32] , 
        \latches_in_f[1][DATA][31] , \latches_in_f[1][DATA][30] , 
        \latches_in_f[1][DATA][29] , \latches_in_f[1][DATA][28] , 
        \latches_in_f[1][DATA][27] , \latches_in_f[1][DATA][26] , 
        \latches_in_f[1][DATA][25] , \latches_in_f[1][DATA][24] , 
        \latches_in_f[1][DATA][23] , \latches_in_f[1][DATA][22] , 
        \latches_in_f[1][DATA][21] , \latches_in_f[1][DATA][20] , 
        \latches_in_f[1][DATA][19] , \latches_in_f[1][DATA][18] , 
        \latches_in_f[1][DATA][17] , \latches_in_f[1][DATA][16] , 
        \latches_in_f[1][DATA][15] , \latches_in_f[1][DATA][14] , 
        \latches_in_f[1][DATA][13] , \latches_in_f[1][DATA][12] , 
        \latches_in_f[1][DATA][11] , \latches_in_f[1][DATA][10] , 
        \latches_in_f[1][DATA][9] , \latches_in_f[1][DATA][8] , 
        \latches_in_f[1][DATA][7] , \latches_in_f[1][DATA][6] , 
        \latches_in_f[1][DATA][5] , \latches_in_f[1][DATA][4] , 
        \latches_in_f[1][DATA][3] , \latches_in_f[1][DATA][2] , 
        \latches_in_f[1][DATA][1] , \latches_in_f[1][DATA][0] }), .left_out(
        \latches_in_b[1][ACK] ), .right_out({\latches_out_f[1][REQ] , 
        \latches_out_f[1][DATA][34] , \latches_out_f[1][DATA][33] , 
        \latches_out_f[1][DATA][32] , \latches_out_f[1][DATA][31] , 
        \latches_out_f[1][DATA][30] , \latches_out_f[1][DATA][29] , 
        \latches_out_f[1][DATA][28] , \latches_out_f[1][DATA][27] , 
        \latches_out_f[1][DATA][26] , \latches_out_f[1][DATA][25] , 
        \latches_out_f[1][DATA][24] , \latches_out_f[1][DATA][23] , 
        \latches_out_f[1][DATA][22] , \latches_out_f[1][DATA][21] , 
        \latches_out_f[1][DATA][20] , \latches_out_f[1][DATA][19] , 
        \latches_out_f[1][DATA][18] , \latches_out_f[1][DATA][17] , 
        \latches_out_f[1][DATA][16] , \latches_out_f[1][DATA][15] , 
        \latches_out_f[1][DATA][14] , \latches_out_f[1][DATA][13] , 
        \latches_out_f[1][DATA][12] , \latches_out_f[1][DATA][11] , 
        \latches_out_f[1][DATA][10] , \latches_out_f[1][DATA][9] , 
        \latches_out_f[1][DATA][8] , \latches_out_f[1][DATA][7] , 
        \latches_out_f[1][DATA][6] , \latches_out_f[1][DATA][5] , 
        \latches_out_f[1][DATA][4] , \latches_out_f[1][DATA][3] , 
        \latches_out_f[1][DATA][2] , \latches_out_f[1][DATA][1] , 
        \latches_out_f[1][DATA][0] }), .right_in(\latches_out_b[1][ACK] ) );
  channel_latch_0_000000000_1 ch_latch_0 ( .preset(n1), .left_in({
        \latches_in_f[0][REQ] , \latches_in_f[0][DATA][34] , 
        \latches_in_f[0][DATA][33] , \latches_in_f[0][DATA][32] , 
        \latches_in_f[0][DATA][31] , \latches_in_f[0][DATA][30] , 
        \latches_in_f[0][DATA][29] , \latches_in_f[0][DATA][28] , 
        \latches_in_f[0][DATA][27] , \latches_in_f[0][DATA][26] , 
        \latches_in_f[0][DATA][25] , \latches_in_f[0][DATA][24] , 
        \latches_in_f[0][DATA][23] , \latches_in_f[0][DATA][22] , 
        \latches_in_f[0][DATA][21] , \latches_in_f[0][DATA][20] , 
        \latches_in_f[0][DATA][19] , \latches_in_f[0][DATA][18] , 
        \latches_in_f[0][DATA][17] , \latches_in_f[0][DATA][16] , 
        \latches_in_f[0][DATA][15] , \latches_in_f[0][DATA][14] , 
        \latches_in_f[0][DATA][13] , \latches_in_f[0][DATA][12] , 
        \latches_in_f[0][DATA][11] , \latches_in_f[0][DATA][10] , 
        \latches_in_f[0][DATA][9] , \latches_in_f[0][DATA][8] , 
        \latches_in_f[0][DATA][7] , \latches_in_f[0][DATA][6] , 
        \latches_in_f[0][DATA][5] , \latches_in_f[0][DATA][4] , 
        \latches_in_f[0][DATA][3] , \latches_in_f[0][DATA][2] , 
        \latches_in_f[0][DATA][1] , \latches_in_f[0][DATA][0] }), .left_out(
        \latches_in_b[0][ACK] ), .right_out({\latches_out_f[0][REQ] , 
        \latches_out_f[0][DATA][34] , \latches_out_f[0][DATA][33] , 
        \latches_out_f[0][DATA][32] , \latches_out_f[0][DATA][31] , 
        \latches_out_f[0][DATA][30] , \latches_out_f[0][DATA][29] , 
        \latches_out_f[0][DATA][28] , \latches_out_f[0][DATA][27] , 
        \latches_out_f[0][DATA][26] , \latches_out_f[0][DATA][25] , 
        \latches_out_f[0][DATA][24] , \latches_out_f[0][DATA][23] , 
        \latches_out_f[0][DATA][22] , \latches_out_f[0][DATA][21] , 
        \latches_out_f[0][DATA][20] , \latches_out_f[0][DATA][19] , 
        \latches_out_f[0][DATA][18] , \latches_out_f[0][DATA][17] , 
        \latches_out_f[0][DATA][16] , \latches_out_f[0][DATA][15] , 
        \latches_out_f[0][DATA][14] , \latches_out_f[0][DATA][13] , 
        \latches_out_f[0][DATA][12] , \latches_out_f[0][DATA][11] , 
        \latches_out_f[0][DATA][10] , \latches_out_f[0][DATA][9] , 
        \latches_out_f[0][DATA][8] , \latches_out_f[0][DATA][7] , 
        \latches_out_f[0][DATA][6] , \latches_out_f[0][DATA][5] , 
        \latches_out_f[0][DATA][4] , \latches_out_f[0][DATA][3] , 
        \latches_out_f[0][DATA][2] , \latches_out_f[0][DATA][1] , 
        \latches_out_f[0][DATA][0] }), .right_in(\latches_out_b[0][ACK] ) );
  HS65_LS_BFX9 U1 ( .A(preset), .Z(n1) );
endmodule


module noc_switch_1 ( preset, .north_in_f({\north_in_f[REQ] , 
        \north_in_f[DATA][34] , \north_in_f[DATA][33] , \north_in_f[DATA][32] , 
        \north_in_f[DATA][31] , \north_in_f[DATA][30] , \north_in_f[DATA][29] , 
        \north_in_f[DATA][28] , \north_in_f[DATA][27] , \north_in_f[DATA][26] , 
        \north_in_f[DATA][25] , \north_in_f[DATA][24] , \north_in_f[DATA][23] , 
        \north_in_f[DATA][22] , \north_in_f[DATA][21] , \north_in_f[DATA][20] , 
        \north_in_f[DATA][19] , \north_in_f[DATA][18] , \north_in_f[DATA][17] , 
        \north_in_f[DATA][16] , \north_in_f[DATA][15] , \north_in_f[DATA][14] , 
        \north_in_f[DATA][13] , \north_in_f[DATA][12] , \north_in_f[DATA][11] , 
        \north_in_f[DATA][10] , \north_in_f[DATA][9] , \north_in_f[DATA][8] , 
        \north_in_f[DATA][7] , \north_in_f[DATA][6] , \north_in_f[DATA][5] , 
        \north_in_f[DATA][4] , \north_in_f[DATA][3] , \north_in_f[DATA][2] , 
        \north_in_f[DATA][1] , \north_in_f[DATA][0] }), .north_in_b(
        \north_in_b[ACK] ), .east_in_f({\east_in_f[REQ] , 
        \east_in_f[DATA][34] , \east_in_f[DATA][33] , \east_in_f[DATA][32] , 
        \east_in_f[DATA][31] , \east_in_f[DATA][30] , \east_in_f[DATA][29] , 
        \east_in_f[DATA][28] , \east_in_f[DATA][27] , \east_in_f[DATA][26] , 
        \east_in_f[DATA][25] , \east_in_f[DATA][24] , \east_in_f[DATA][23] , 
        \east_in_f[DATA][22] , \east_in_f[DATA][21] , \east_in_f[DATA][20] , 
        \east_in_f[DATA][19] , \east_in_f[DATA][18] , \east_in_f[DATA][17] , 
        \east_in_f[DATA][16] , \east_in_f[DATA][15] , \east_in_f[DATA][14] , 
        \east_in_f[DATA][13] , \east_in_f[DATA][12] , \east_in_f[DATA][11] , 
        \east_in_f[DATA][10] , \east_in_f[DATA][9] , \east_in_f[DATA][8] , 
        \east_in_f[DATA][7] , \east_in_f[DATA][6] , \east_in_f[DATA][5] , 
        \east_in_f[DATA][4] , \east_in_f[DATA][3] , \east_in_f[DATA][2] , 
        \east_in_f[DATA][1] , \east_in_f[DATA][0] }), .east_in_b(
        \east_in_b[ACK] ), .south_in_f({\south_in_f[REQ] , 
        \south_in_f[DATA][34] , \south_in_f[DATA][33] , \south_in_f[DATA][32] , 
        \south_in_f[DATA][31] , \south_in_f[DATA][30] , \south_in_f[DATA][29] , 
        \south_in_f[DATA][28] , \south_in_f[DATA][27] , \south_in_f[DATA][26] , 
        \south_in_f[DATA][25] , \south_in_f[DATA][24] , \south_in_f[DATA][23] , 
        \south_in_f[DATA][22] , \south_in_f[DATA][21] , \south_in_f[DATA][20] , 
        \south_in_f[DATA][19] , \south_in_f[DATA][18] , \south_in_f[DATA][17] , 
        \south_in_f[DATA][16] , \south_in_f[DATA][15] , \south_in_f[DATA][14] , 
        \south_in_f[DATA][13] , \south_in_f[DATA][12] , \south_in_f[DATA][11] , 
        \south_in_f[DATA][10] , \south_in_f[DATA][9] , \south_in_f[DATA][8] , 
        \south_in_f[DATA][7] , \south_in_f[DATA][6] , \south_in_f[DATA][5] , 
        \south_in_f[DATA][4] , \south_in_f[DATA][3] , \south_in_f[DATA][2] , 
        \south_in_f[DATA][1] , \south_in_f[DATA][0] }), .south_in_b(
        \south_in_b[ACK] ), .west_in_f({\west_in_f[REQ] , 
        \west_in_f[DATA][34] , \west_in_f[DATA][33] , \west_in_f[DATA][32] , 
        \west_in_f[DATA][31] , \west_in_f[DATA][30] , \west_in_f[DATA][29] , 
        \west_in_f[DATA][28] , \west_in_f[DATA][27] , \west_in_f[DATA][26] , 
        \west_in_f[DATA][25] , \west_in_f[DATA][24] , \west_in_f[DATA][23] , 
        \west_in_f[DATA][22] , \west_in_f[DATA][21] , \west_in_f[DATA][20] , 
        \west_in_f[DATA][19] , \west_in_f[DATA][18] , \west_in_f[DATA][17] , 
        \west_in_f[DATA][16] , \west_in_f[DATA][15] , \west_in_f[DATA][14] , 
        \west_in_f[DATA][13] , \west_in_f[DATA][12] , \west_in_f[DATA][11] , 
        \west_in_f[DATA][10] , \west_in_f[DATA][9] , \west_in_f[DATA][8] , 
        \west_in_f[DATA][7] , \west_in_f[DATA][6] , \west_in_f[DATA][5] , 
        \west_in_f[DATA][4] , \west_in_f[DATA][3] , \west_in_f[DATA][2] , 
        \west_in_f[DATA][1] , \west_in_f[DATA][0] }), .west_in_b(
        \west_in_b[ACK] ), .resource_in_f({\resource_in_f[REQ] , 
        \resource_in_f[DATA][34] , \resource_in_f[DATA][33] , 
        \resource_in_f[DATA][32] , \resource_in_f[DATA][31] , 
        \resource_in_f[DATA][30] , \resource_in_f[DATA][29] , 
        \resource_in_f[DATA][28] , \resource_in_f[DATA][27] , 
        \resource_in_f[DATA][26] , \resource_in_f[DATA][25] , 
        \resource_in_f[DATA][24] , \resource_in_f[DATA][23] , 
        \resource_in_f[DATA][22] , \resource_in_f[DATA][21] , 
        \resource_in_f[DATA][20] , \resource_in_f[DATA][19] , 
        \resource_in_f[DATA][18] , \resource_in_f[DATA][17] , 
        \resource_in_f[DATA][16] , \resource_in_f[DATA][15] , 
        \resource_in_f[DATA][14] , \resource_in_f[DATA][13] , 
        \resource_in_f[DATA][12] , \resource_in_f[DATA][11] , 
        \resource_in_f[DATA][10] , \resource_in_f[DATA][9] , 
        \resource_in_f[DATA][8] , \resource_in_f[DATA][7] , 
        \resource_in_f[DATA][6] , \resource_in_f[DATA][5] , 
        \resource_in_f[DATA][4] , \resource_in_f[DATA][3] , 
        \resource_in_f[DATA][2] , \resource_in_f[DATA][1] , 
        \resource_in_f[DATA][0] }), .resource_in_b(\resource_in_b[ACK] ), 
    .north_out_f({\north_out_f[REQ] , \north_out_f[DATA][34] , 
        \north_out_f[DATA][33] , \north_out_f[DATA][32] , 
        \north_out_f[DATA][31] , \north_out_f[DATA][30] , 
        \north_out_f[DATA][29] , \north_out_f[DATA][28] , 
        \north_out_f[DATA][27] , \north_out_f[DATA][26] , 
        \north_out_f[DATA][25] , \north_out_f[DATA][24] , 
        \north_out_f[DATA][23] , \north_out_f[DATA][22] , 
        \north_out_f[DATA][21] , \north_out_f[DATA][20] , 
        \north_out_f[DATA][19] , \north_out_f[DATA][18] , 
        \north_out_f[DATA][17] , \north_out_f[DATA][16] , 
        \north_out_f[DATA][15] , \north_out_f[DATA][14] , 
        \north_out_f[DATA][13] , \north_out_f[DATA][12] , 
        \north_out_f[DATA][11] , \north_out_f[DATA][10] , 
        \north_out_f[DATA][9] , \north_out_f[DATA][8] , \north_out_f[DATA][7] , 
        \north_out_f[DATA][6] , \north_out_f[DATA][5] , \north_out_f[DATA][4] , 
        \north_out_f[DATA][3] , \north_out_f[DATA][2] , \north_out_f[DATA][1] , 
        \north_out_f[DATA][0] }), .north_out_b(\north_out_b[ACK] ), 
    .east_out_f({\east_out_f[REQ] , \east_out_f[DATA][34] , 
        \east_out_f[DATA][33] , \east_out_f[DATA][32] , \east_out_f[DATA][31] , 
        \east_out_f[DATA][30] , \east_out_f[DATA][29] , \east_out_f[DATA][28] , 
        \east_out_f[DATA][27] , \east_out_f[DATA][26] , \east_out_f[DATA][25] , 
        \east_out_f[DATA][24] , \east_out_f[DATA][23] , \east_out_f[DATA][22] , 
        \east_out_f[DATA][21] , \east_out_f[DATA][20] , \east_out_f[DATA][19] , 
        \east_out_f[DATA][18] , \east_out_f[DATA][17] , \east_out_f[DATA][16] , 
        \east_out_f[DATA][15] , \east_out_f[DATA][14] , \east_out_f[DATA][13] , 
        \east_out_f[DATA][12] , \east_out_f[DATA][11] , \east_out_f[DATA][10] , 
        \east_out_f[DATA][9] , \east_out_f[DATA][8] , \east_out_f[DATA][7] , 
        \east_out_f[DATA][6] , \east_out_f[DATA][5] , \east_out_f[DATA][4] , 
        \east_out_f[DATA][3] , \east_out_f[DATA][2] , \east_out_f[DATA][1] , 
        \east_out_f[DATA][0] }), .east_out_b(\east_out_b[ACK] ), 
    .south_out_f({\south_out_f[REQ] , \south_out_f[DATA][34] , 
        \south_out_f[DATA][33] , \south_out_f[DATA][32] , 
        \south_out_f[DATA][31] , \south_out_f[DATA][30] , 
        \south_out_f[DATA][29] , \south_out_f[DATA][28] , 
        \south_out_f[DATA][27] , \south_out_f[DATA][26] , 
        \south_out_f[DATA][25] , \south_out_f[DATA][24] , 
        \south_out_f[DATA][23] , \south_out_f[DATA][22] , 
        \south_out_f[DATA][21] , \south_out_f[DATA][20] , 
        \south_out_f[DATA][19] , \south_out_f[DATA][18] , 
        \south_out_f[DATA][17] , \south_out_f[DATA][16] , 
        \south_out_f[DATA][15] , \south_out_f[DATA][14] , 
        \south_out_f[DATA][13] , \south_out_f[DATA][12] , 
        \south_out_f[DATA][11] , \south_out_f[DATA][10] , 
        \south_out_f[DATA][9] , \south_out_f[DATA][8] , \south_out_f[DATA][7] , 
        \south_out_f[DATA][6] , \south_out_f[DATA][5] , \south_out_f[DATA][4] , 
        \south_out_f[DATA][3] , \south_out_f[DATA][2] , \south_out_f[DATA][1] , 
        \south_out_f[DATA][0] }), .south_out_b(\south_out_b[ACK] ), 
    .west_out_f({\west_out_f[REQ] , \west_out_f[DATA][34] , 
        \west_out_f[DATA][33] , \west_out_f[DATA][32] , \west_out_f[DATA][31] , 
        \west_out_f[DATA][30] , \west_out_f[DATA][29] , \west_out_f[DATA][28] , 
        \west_out_f[DATA][27] , \west_out_f[DATA][26] , \west_out_f[DATA][25] , 
        \west_out_f[DATA][24] , \west_out_f[DATA][23] , \west_out_f[DATA][22] , 
        \west_out_f[DATA][21] , \west_out_f[DATA][20] , \west_out_f[DATA][19] , 
        \west_out_f[DATA][18] , \west_out_f[DATA][17] , \west_out_f[DATA][16] , 
        \west_out_f[DATA][15] , \west_out_f[DATA][14] , \west_out_f[DATA][13] , 
        \west_out_f[DATA][12] , \west_out_f[DATA][11] , \west_out_f[DATA][10] , 
        \west_out_f[DATA][9] , \west_out_f[DATA][8] , \west_out_f[DATA][7] , 
        \west_out_f[DATA][6] , \west_out_f[DATA][5] , \west_out_f[DATA][4] , 
        \west_out_f[DATA][3] , \west_out_f[DATA][2] , \west_out_f[DATA][1] , 
        \west_out_f[DATA][0] }), .west_out_b(\west_out_b[ACK] ), 
    .resource_out_f({\resource_out_f[REQ] , \resource_out_f[DATA][34] , 
        \resource_out_f[DATA][33] , \resource_out_f[DATA][32] , 
        \resource_out_f[DATA][31] , \resource_out_f[DATA][30] , 
        \resource_out_f[DATA][29] , \resource_out_f[DATA][28] , 
        \resource_out_f[DATA][27] , \resource_out_f[DATA][26] , 
        \resource_out_f[DATA][25] , \resource_out_f[DATA][24] , 
        \resource_out_f[DATA][23] , \resource_out_f[DATA][22] , 
        \resource_out_f[DATA][21] , \resource_out_f[DATA][20] , 
        \resource_out_f[DATA][19] , \resource_out_f[DATA][18] , 
        \resource_out_f[DATA][17] , \resource_out_f[DATA][16] , 
        \resource_out_f[DATA][15] , \resource_out_f[DATA][14] , 
        \resource_out_f[DATA][13] , \resource_out_f[DATA][12] , 
        \resource_out_f[DATA][11] , \resource_out_f[DATA][10] , 
        \resource_out_f[DATA][9] , \resource_out_f[DATA][8] , 
        \resource_out_f[DATA][7] , \resource_out_f[DATA][6] , 
        \resource_out_f[DATA][5] , \resource_out_f[DATA][4] , 
        \resource_out_f[DATA][3] , \resource_out_f[DATA][2] , 
        \resource_out_f[DATA][1] , \resource_out_f[DATA][0] }), 
    .resource_out_b(\resource_out_b[ACK] ) );
  input preset, \north_in_f[REQ] , \north_in_f[DATA][34] ,
         \north_in_f[DATA][33] , \north_in_f[DATA][32] ,
         \north_in_f[DATA][31] , \north_in_f[DATA][30] ,
         \north_in_f[DATA][29] , \north_in_f[DATA][28] ,
         \north_in_f[DATA][27] , \north_in_f[DATA][26] ,
         \north_in_f[DATA][25] , \north_in_f[DATA][24] ,
         \north_in_f[DATA][23] , \north_in_f[DATA][22] ,
         \north_in_f[DATA][21] , \north_in_f[DATA][20] ,
         \north_in_f[DATA][19] , \north_in_f[DATA][18] ,
         \north_in_f[DATA][17] , \north_in_f[DATA][16] ,
         \north_in_f[DATA][15] , \north_in_f[DATA][14] ,
         \north_in_f[DATA][13] , \north_in_f[DATA][12] ,
         \north_in_f[DATA][11] , \north_in_f[DATA][10] , \north_in_f[DATA][9] ,
         \north_in_f[DATA][8] , \north_in_f[DATA][7] , \north_in_f[DATA][6] ,
         \north_in_f[DATA][5] , \north_in_f[DATA][4] , \north_in_f[DATA][3] ,
         \north_in_f[DATA][2] , \north_in_f[DATA][1] , \north_in_f[DATA][0] ,
         \east_in_f[REQ] , \east_in_f[DATA][34] , \east_in_f[DATA][33] ,
         \east_in_f[DATA][32] , \east_in_f[DATA][31] , \east_in_f[DATA][30] ,
         \east_in_f[DATA][29] , \east_in_f[DATA][28] , \east_in_f[DATA][27] ,
         \east_in_f[DATA][26] , \east_in_f[DATA][25] , \east_in_f[DATA][24] ,
         \east_in_f[DATA][23] , \east_in_f[DATA][22] , \east_in_f[DATA][21] ,
         \east_in_f[DATA][20] , \east_in_f[DATA][19] , \east_in_f[DATA][18] ,
         \east_in_f[DATA][17] , \east_in_f[DATA][16] , \east_in_f[DATA][15] ,
         \east_in_f[DATA][14] , \east_in_f[DATA][13] , \east_in_f[DATA][12] ,
         \east_in_f[DATA][11] , \east_in_f[DATA][10] , \east_in_f[DATA][9] ,
         \east_in_f[DATA][8] , \east_in_f[DATA][7] , \east_in_f[DATA][6] ,
         \east_in_f[DATA][5] , \east_in_f[DATA][4] , \east_in_f[DATA][3] ,
         \east_in_f[DATA][2] , \east_in_f[DATA][1] , \east_in_f[DATA][0] ,
         \south_in_f[REQ] , \south_in_f[DATA][34] , \south_in_f[DATA][33] ,
         \south_in_f[DATA][32] , \south_in_f[DATA][31] ,
         \south_in_f[DATA][30] , \south_in_f[DATA][29] ,
         \south_in_f[DATA][28] , \south_in_f[DATA][27] ,
         \south_in_f[DATA][26] , \south_in_f[DATA][25] ,
         \south_in_f[DATA][24] , \south_in_f[DATA][23] ,
         \south_in_f[DATA][22] , \south_in_f[DATA][21] ,
         \south_in_f[DATA][20] , \south_in_f[DATA][19] ,
         \south_in_f[DATA][18] , \south_in_f[DATA][17] ,
         \south_in_f[DATA][16] , \south_in_f[DATA][15] ,
         \south_in_f[DATA][14] , \south_in_f[DATA][13] ,
         \south_in_f[DATA][12] , \south_in_f[DATA][11] ,
         \south_in_f[DATA][10] , \south_in_f[DATA][9] , \south_in_f[DATA][8] ,
         \south_in_f[DATA][7] , \south_in_f[DATA][6] , \south_in_f[DATA][5] ,
         \south_in_f[DATA][4] , \south_in_f[DATA][3] , \south_in_f[DATA][2] ,
         \south_in_f[DATA][1] , \south_in_f[DATA][0] , \west_in_f[REQ] ,
         \west_in_f[DATA][34] , \west_in_f[DATA][33] , \west_in_f[DATA][32] ,
         \west_in_f[DATA][31] , \west_in_f[DATA][30] , \west_in_f[DATA][29] ,
         \west_in_f[DATA][28] , \west_in_f[DATA][27] , \west_in_f[DATA][26] ,
         \west_in_f[DATA][25] , \west_in_f[DATA][24] , \west_in_f[DATA][23] ,
         \west_in_f[DATA][22] , \west_in_f[DATA][21] , \west_in_f[DATA][20] ,
         \west_in_f[DATA][19] , \west_in_f[DATA][18] , \west_in_f[DATA][17] ,
         \west_in_f[DATA][16] , \west_in_f[DATA][15] , \west_in_f[DATA][14] ,
         \west_in_f[DATA][13] , \west_in_f[DATA][12] , \west_in_f[DATA][11] ,
         \west_in_f[DATA][10] , \west_in_f[DATA][9] , \west_in_f[DATA][8] ,
         \west_in_f[DATA][7] , \west_in_f[DATA][6] , \west_in_f[DATA][5] ,
         \west_in_f[DATA][4] , \west_in_f[DATA][3] , \west_in_f[DATA][2] ,
         \west_in_f[DATA][1] , \west_in_f[DATA][0] , \resource_in_f[REQ] ,
         \resource_in_f[DATA][34] , \resource_in_f[DATA][33] ,
         \resource_in_f[DATA][32] , \resource_in_f[DATA][31] ,
         \resource_in_f[DATA][30] , \resource_in_f[DATA][29] ,
         \resource_in_f[DATA][28] , \resource_in_f[DATA][27] ,
         \resource_in_f[DATA][26] , \resource_in_f[DATA][25] ,
         \resource_in_f[DATA][24] , \resource_in_f[DATA][23] ,
         \resource_in_f[DATA][22] , \resource_in_f[DATA][21] ,
         \resource_in_f[DATA][20] , \resource_in_f[DATA][19] ,
         \resource_in_f[DATA][18] , \resource_in_f[DATA][17] ,
         \resource_in_f[DATA][16] , \resource_in_f[DATA][15] ,
         \resource_in_f[DATA][14] , \resource_in_f[DATA][13] ,
         \resource_in_f[DATA][12] , \resource_in_f[DATA][11] ,
         \resource_in_f[DATA][10] , \resource_in_f[DATA][9] ,
         \resource_in_f[DATA][8] , \resource_in_f[DATA][7] ,
         \resource_in_f[DATA][6] , \resource_in_f[DATA][5] ,
         \resource_in_f[DATA][4] , \resource_in_f[DATA][3] ,
         \resource_in_f[DATA][2] , \resource_in_f[DATA][1] ,
         \resource_in_f[DATA][0] , \north_out_b[ACK] , \east_out_b[ACK] ,
         \south_out_b[ACK] , \west_out_b[ACK] , \resource_out_b[ACK] ;
  output \north_in_b[ACK] , \east_in_b[ACK] , \south_in_b[ACK] ,
         \west_in_b[ACK] , \resource_in_b[ACK] , \north_out_f[REQ] ,
         \north_out_f[DATA][34] , \north_out_f[DATA][33] ,
         \north_out_f[DATA][32] , \north_out_f[DATA][31] ,
         \north_out_f[DATA][30] , \north_out_f[DATA][29] ,
         \north_out_f[DATA][28] , \north_out_f[DATA][27] ,
         \north_out_f[DATA][26] , \north_out_f[DATA][25] ,
         \north_out_f[DATA][24] , \north_out_f[DATA][23] ,
         \north_out_f[DATA][22] , \north_out_f[DATA][21] ,
         \north_out_f[DATA][20] , \north_out_f[DATA][19] ,
         \north_out_f[DATA][18] , \north_out_f[DATA][17] ,
         \north_out_f[DATA][16] , \north_out_f[DATA][15] ,
         \north_out_f[DATA][14] , \north_out_f[DATA][13] ,
         \north_out_f[DATA][12] , \north_out_f[DATA][11] ,
         \north_out_f[DATA][10] , \north_out_f[DATA][9] ,
         \north_out_f[DATA][8] , \north_out_f[DATA][7] ,
         \north_out_f[DATA][6] , \north_out_f[DATA][5] ,
         \north_out_f[DATA][4] , \north_out_f[DATA][3] ,
         \north_out_f[DATA][2] , \north_out_f[DATA][1] ,
         \north_out_f[DATA][0] , \east_out_f[REQ] , \east_out_f[DATA][34] ,
         \east_out_f[DATA][33] , \east_out_f[DATA][32] ,
         \east_out_f[DATA][31] , \east_out_f[DATA][30] ,
         \east_out_f[DATA][29] , \east_out_f[DATA][28] ,
         \east_out_f[DATA][27] , \east_out_f[DATA][26] ,
         \east_out_f[DATA][25] , \east_out_f[DATA][24] ,
         \east_out_f[DATA][23] , \east_out_f[DATA][22] ,
         \east_out_f[DATA][21] , \east_out_f[DATA][20] ,
         \east_out_f[DATA][19] , \east_out_f[DATA][18] ,
         \east_out_f[DATA][17] , \east_out_f[DATA][16] ,
         \east_out_f[DATA][15] , \east_out_f[DATA][14] ,
         \east_out_f[DATA][13] , \east_out_f[DATA][12] ,
         \east_out_f[DATA][11] , \east_out_f[DATA][10] , \east_out_f[DATA][9] ,
         \east_out_f[DATA][8] , \east_out_f[DATA][7] , \east_out_f[DATA][6] ,
         \east_out_f[DATA][5] , \east_out_f[DATA][4] , \east_out_f[DATA][3] ,
         \east_out_f[DATA][2] , \east_out_f[DATA][1] , \east_out_f[DATA][0] ,
         \south_out_f[REQ] , \south_out_f[DATA][34] , \south_out_f[DATA][33] ,
         \south_out_f[DATA][32] , \south_out_f[DATA][31] ,
         \south_out_f[DATA][30] , \south_out_f[DATA][29] ,
         \south_out_f[DATA][28] , \south_out_f[DATA][27] ,
         \south_out_f[DATA][26] , \south_out_f[DATA][25] ,
         \south_out_f[DATA][24] , \south_out_f[DATA][23] ,
         \south_out_f[DATA][22] , \south_out_f[DATA][21] ,
         \south_out_f[DATA][20] , \south_out_f[DATA][19] ,
         \south_out_f[DATA][18] , \south_out_f[DATA][17] ,
         \south_out_f[DATA][16] , \south_out_f[DATA][15] ,
         \south_out_f[DATA][14] , \south_out_f[DATA][13] ,
         \south_out_f[DATA][12] , \south_out_f[DATA][11] ,
         \south_out_f[DATA][10] , \south_out_f[DATA][9] ,
         \south_out_f[DATA][8] , \south_out_f[DATA][7] ,
         \south_out_f[DATA][6] , \south_out_f[DATA][5] ,
         \south_out_f[DATA][4] , \south_out_f[DATA][3] ,
         \south_out_f[DATA][2] , \south_out_f[DATA][1] ,
         \south_out_f[DATA][0] , \west_out_f[REQ] , \west_out_f[DATA][34] ,
         \west_out_f[DATA][33] , \west_out_f[DATA][32] ,
         \west_out_f[DATA][31] , \west_out_f[DATA][30] ,
         \west_out_f[DATA][29] , \west_out_f[DATA][28] ,
         \west_out_f[DATA][27] , \west_out_f[DATA][26] ,
         \west_out_f[DATA][25] , \west_out_f[DATA][24] ,
         \west_out_f[DATA][23] , \west_out_f[DATA][22] ,
         \west_out_f[DATA][21] , \west_out_f[DATA][20] ,
         \west_out_f[DATA][19] , \west_out_f[DATA][18] ,
         \west_out_f[DATA][17] , \west_out_f[DATA][16] ,
         \west_out_f[DATA][15] , \west_out_f[DATA][14] ,
         \west_out_f[DATA][13] , \west_out_f[DATA][12] ,
         \west_out_f[DATA][11] , \west_out_f[DATA][10] , \west_out_f[DATA][9] ,
         \west_out_f[DATA][8] , \west_out_f[DATA][7] , \west_out_f[DATA][6] ,
         \west_out_f[DATA][5] , \west_out_f[DATA][4] , \west_out_f[DATA][3] ,
         \west_out_f[DATA][2] , \west_out_f[DATA][1] , \west_out_f[DATA][0] ,
         \resource_out_f[REQ] , \resource_out_f[DATA][34] ,
         \resource_out_f[DATA][33] , \resource_out_f[DATA][32] ,
         \resource_out_f[DATA][31] , \resource_out_f[DATA][30] ,
         \resource_out_f[DATA][29] , \resource_out_f[DATA][28] ,
         \resource_out_f[DATA][27] , \resource_out_f[DATA][26] ,
         \resource_out_f[DATA][25] , \resource_out_f[DATA][24] ,
         \resource_out_f[DATA][23] , \resource_out_f[DATA][22] ,
         \resource_out_f[DATA][21] , \resource_out_f[DATA][20] ,
         \resource_out_f[DATA][19] , \resource_out_f[DATA][18] ,
         \resource_out_f[DATA][17] , \resource_out_f[DATA][16] ,
         \resource_out_f[DATA][15] , \resource_out_f[DATA][14] ,
         \resource_out_f[DATA][13] , \resource_out_f[DATA][12] ,
         \resource_out_f[DATA][11] , \resource_out_f[DATA][10] ,
         \resource_out_f[DATA][9] , \resource_out_f[DATA][8] ,
         \resource_out_f[DATA][7] , \resource_out_f[DATA][6] ,
         \resource_out_f[DATA][5] , \resource_out_f[DATA][4] ,
         \resource_out_f[DATA][3] , \resource_out_f[DATA][2] ,
         \resource_out_f[DATA][1] , \resource_out_f[DATA][0] ;
  wire   \north_hpu_f[REQ] , \north_hpu_f[DATA][34] , \north_hpu_f[DATA][33] ,
         \north_hpu_f[DATA][32] , \north_hpu_f[DATA][31] ,
         \north_hpu_f[DATA][30] , \north_hpu_f[DATA][29] ,
         \north_hpu_f[DATA][28] , \north_hpu_f[DATA][27] ,
         \north_hpu_f[DATA][26] , \north_hpu_f[DATA][25] ,
         \north_hpu_f[DATA][24] , \north_hpu_f[DATA][23] ,
         \north_hpu_f[DATA][22] , \north_hpu_f[DATA][21] ,
         \north_hpu_f[DATA][20] , \north_hpu_f[DATA][19] ,
         \north_hpu_f[DATA][18] , \north_hpu_f[DATA][17] ,
         \north_hpu_f[DATA][16] , \north_hpu_f[DATA][15] ,
         \north_hpu_f[DATA][14] , \north_hpu_f[DATA][13] ,
         \north_hpu_f[DATA][12] , \north_hpu_f[DATA][11] ,
         \north_hpu_f[DATA][10] , \north_hpu_f[DATA][9] ,
         \north_hpu_f[DATA][8] , \north_hpu_f[DATA][7] ,
         \north_hpu_f[DATA][6] , \north_hpu_f[DATA][5] ,
         \north_hpu_f[DATA][4] , \north_hpu_f[DATA][3] ,
         \north_hpu_f[DATA][2] , \north_hpu_f[DATA][1] ,
         \north_hpu_f[DATA][0] , \north_hpu_b[ACK] , \south_hpu_f[REQ] ,
         \south_hpu_f[DATA][34] , \south_hpu_f[DATA][33] ,
         \south_hpu_f[DATA][32] , \south_hpu_f[DATA][31] ,
         \south_hpu_f[DATA][30] , \south_hpu_f[DATA][29] ,
         \south_hpu_f[DATA][28] , \south_hpu_f[DATA][27] ,
         \south_hpu_f[DATA][26] , \south_hpu_f[DATA][25] ,
         \south_hpu_f[DATA][24] , \south_hpu_f[DATA][23] ,
         \south_hpu_f[DATA][22] , \south_hpu_f[DATA][21] ,
         \south_hpu_f[DATA][20] , \south_hpu_f[DATA][19] ,
         \south_hpu_f[DATA][18] , \south_hpu_f[DATA][17] ,
         \south_hpu_f[DATA][16] , \south_hpu_f[DATA][15] ,
         \south_hpu_f[DATA][14] , \south_hpu_f[DATA][13] ,
         \south_hpu_f[DATA][12] , \south_hpu_f[DATA][11] ,
         \south_hpu_f[DATA][10] , \south_hpu_f[DATA][9] ,
         \south_hpu_f[DATA][8] , \south_hpu_f[DATA][7] ,
         \south_hpu_f[DATA][6] , \south_hpu_f[DATA][5] ,
         \south_hpu_f[DATA][4] , \south_hpu_f[DATA][3] ,
         \south_hpu_f[DATA][2] , \south_hpu_f[DATA][1] ,
         \south_hpu_f[DATA][0] , \south_hpu_b[ACK] , \east_hpu_f[REQ] ,
         \east_hpu_f[DATA][34] , \east_hpu_f[DATA][33] ,
         \east_hpu_f[DATA][32] , \east_hpu_f[DATA][31] ,
         \east_hpu_f[DATA][30] , \east_hpu_f[DATA][29] ,
         \east_hpu_f[DATA][28] , \east_hpu_f[DATA][27] ,
         \east_hpu_f[DATA][26] , \east_hpu_f[DATA][25] ,
         \east_hpu_f[DATA][24] , \east_hpu_f[DATA][23] ,
         \east_hpu_f[DATA][22] , \east_hpu_f[DATA][21] ,
         \east_hpu_f[DATA][20] , \east_hpu_f[DATA][19] ,
         \east_hpu_f[DATA][18] , \east_hpu_f[DATA][17] ,
         \east_hpu_f[DATA][16] , \east_hpu_f[DATA][15] ,
         \east_hpu_f[DATA][14] , \east_hpu_f[DATA][13] ,
         \east_hpu_f[DATA][12] , \east_hpu_f[DATA][11] ,
         \east_hpu_f[DATA][10] , \east_hpu_f[DATA][9] , \east_hpu_f[DATA][8] ,
         \east_hpu_f[DATA][7] , \east_hpu_f[DATA][6] , \east_hpu_f[DATA][5] ,
         \east_hpu_f[DATA][4] , \east_hpu_f[DATA][3] , \east_hpu_f[DATA][2] ,
         \east_hpu_f[DATA][1] , \east_hpu_f[DATA][0] , \east_hpu_b[ACK] ,
         \west_hpu_f[REQ] , \west_hpu_f[DATA][34] , \west_hpu_f[DATA][33] ,
         \west_hpu_f[DATA][32] , \west_hpu_f[DATA][31] ,
         \west_hpu_f[DATA][30] , \west_hpu_f[DATA][29] ,
         \west_hpu_f[DATA][28] , \west_hpu_f[DATA][27] ,
         \west_hpu_f[DATA][26] , \west_hpu_f[DATA][25] ,
         \west_hpu_f[DATA][24] , \west_hpu_f[DATA][23] ,
         \west_hpu_f[DATA][22] , \west_hpu_f[DATA][21] ,
         \west_hpu_f[DATA][20] , \west_hpu_f[DATA][19] ,
         \west_hpu_f[DATA][18] , \west_hpu_f[DATA][17] ,
         \west_hpu_f[DATA][16] , \west_hpu_f[DATA][15] ,
         \west_hpu_f[DATA][14] , \west_hpu_f[DATA][13] ,
         \west_hpu_f[DATA][12] , \west_hpu_f[DATA][11] ,
         \west_hpu_f[DATA][10] , \west_hpu_f[DATA][9] , \west_hpu_f[DATA][8] ,
         \west_hpu_f[DATA][7] , \west_hpu_f[DATA][6] , \west_hpu_f[DATA][5] ,
         \west_hpu_f[DATA][4] , \west_hpu_f[DATA][3] , \west_hpu_f[DATA][2] ,
         \west_hpu_f[DATA][1] , \west_hpu_f[DATA][0] , \west_hpu_b[ACK] ,
         \resource_hpu_f[REQ] , \resource_hpu_f[DATA][34] ,
         \resource_hpu_f[DATA][33] , \resource_hpu_f[DATA][32] ,
         \resource_hpu_f[DATA][31] , \resource_hpu_f[DATA][30] ,
         \resource_hpu_f[DATA][29] , \resource_hpu_f[DATA][28] ,
         \resource_hpu_f[DATA][27] , \resource_hpu_f[DATA][26] ,
         \resource_hpu_f[DATA][25] , \resource_hpu_f[DATA][24] ,
         \resource_hpu_f[DATA][23] , \resource_hpu_f[DATA][22] ,
         \resource_hpu_f[DATA][21] , \resource_hpu_f[DATA][20] ,
         \resource_hpu_f[DATA][19] , \resource_hpu_f[DATA][18] ,
         \resource_hpu_f[DATA][17] , \resource_hpu_f[DATA][16] ,
         \resource_hpu_f[DATA][15] , \resource_hpu_f[DATA][14] ,
         \resource_hpu_f[DATA][13] , \resource_hpu_f[DATA][12] ,
         \resource_hpu_f[DATA][11] , \resource_hpu_f[DATA][10] ,
         \resource_hpu_f[DATA][9] , \resource_hpu_f[DATA][8] ,
         \resource_hpu_f[DATA][7] , \resource_hpu_f[DATA][6] ,
         \resource_hpu_f[DATA][5] , \resource_hpu_f[DATA][4] ,
         \resource_hpu_f[DATA][3] , \resource_hpu_f[DATA][2] ,
         \resource_hpu_f[DATA][1] , \resource_hpu_f[DATA][0] ,
         \resource_hpu_b[ACK] , \chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] ,
         \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] ,
         \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] ,
         \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] ,
         \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] ,
         \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] ,
         \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] ,
         \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] ,
         \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] ,
         \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] ,
         \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] ,
         \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] ,
         \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] ,
         \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] ,
         \chs_in_f[4][DATA][7] , \chs_in_f[4][DATA][6] ,
         \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] ,
         \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] ,
         \chs_in_f[4][DATA][1] , \chs_in_f[4][DATA][0] , \chs_in_f[3][REQ] ,
         \chs_in_f[3][DATA][34] , \chs_in_f[3][DATA][33] ,
         \chs_in_f[3][DATA][32] , \chs_in_f[3][DATA][31] ,
         \chs_in_f[3][DATA][30] , \chs_in_f[3][DATA][29] ,
         \chs_in_f[3][DATA][28] , \chs_in_f[3][DATA][27] ,
         \chs_in_f[3][DATA][26] , \chs_in_f[3][DATA][25] ,
         \chs_in_f[3][DATA][24] , \chs_in_f[3][DATA][23] ,
         \chs_in_f[3][DATA][22] , \chs_in_f[3][DATA][21] ,
         \chs_in_f[3][DATA][20] , \chs_in_f[3][DATA][19] ,
         \chs_in_f[3][DATA][18] , \chs_in_f[3][DATA][17] ,
         \chs_in_f[3][DATA][16] , \chs_in_f[3][DATA][15] ,
         \chs_in_f[3][DATA][14] , \chs_in_f[3][DATA][13] ,
         \chs_in_f[3][DATA][12] , \chs_in_f[3][DATA][11] ,
         \chs_in_f[3][DATA][10] , \chs_in_f[3][DATA][9] ,
         \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] ,
         \chs_in_f[3][DATA][6] , \chs_in_f[3][DATA][5] ,
         \chs_in_f[3][DATA][4] , \chs_in_f[3][DATA][3] ,
         \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] ,
         \chs_in_f[3][DATA][0] , \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] ,
         \chs_in_f[2][DATA][33] , \chs_in_f[2][DATA][32] ,
         \chs_in_f[2][DATA][31] , \chs_in_f[2][DATA][30] ,
         \chs_in_f[2][DATA][29] , \chs_in_f[2][DATA][28] ,
         \chs_in_f[2][DATA][27] , \chs_in_f[2][DATA][26] ,
         \chs_in_f[2][DATA][25] , \chs_in_f[2][DATA][24] ,
         \chs_in_f[2][DATA][23] , \chs_in_f[2][DATA][22] ,
         \chs_in_f[2][DATA][21] , \chs_in_f[2][DATA][20] ,
         \chs_in_f[2][DATA][19] , \chs_in_f[2][DATA][18] ,
         \chs_in_f[2][DATA][17] , \chs_in_f[2][DATA][16] ,
         \chs_in_f[2][DATA][15] , \chs_in_f[2][DATA][14] ,
         \chs_in_f[2][DATA][13] , \chs_in_f[2][DATA][12] ,
         \chs_in_f[2][DATA][11] , \chs_in_f[2][DATA][10] ,
         \chs_in_f[2][DATA][9] , \chs_in_f[2][DATA][8] ,
         \chs_in_f[2][DATA][7] , \chs_in_f[2][DATA][6] ,
         \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] ,
         \chs_in_f[2][DATA][3] , \chs_in_f[2][DATA][2] ,
         \chs_in_f[2][DATA][1] , \chs_in_f[2][DATA][0] , \chs_in_f[1][REQ] ,
         \chs_in_f[1][DATA][34] , \chs_in_f[1][DATA][33] ,
         \chs_in_f[1][DATA][32] , \chs_in_f[1][DATA][31] ,
         \chs_in_f[1][DATA][30] , \chs_in_f[1][DATA][29] ,
         \chs_in_f[1][DATA][28] , \chs_in_f[1][DATA][27] ,
         \chs_in_f[1][DATA][26] , \chs_in_f[1][DATA][25] ,
         \chs_in_f[1][DATA][24] , \chs_in_f[1][DATA][23] ,
         \chs_in_f[1][DATA][22] , \chs_in_f[1][DATA][21] ,
         \chs_in_f[1][DATA][20] , \chs_in_f[1][DATA][19] ,
         \chs_in_f[1][DATA][18] , \chs_in_f[1][DATA][17] ,
         \chs_in_f[1][DATA][16] , \chs_in_f[1][DATA][15] ,
         \chs_in_f[1][DATA][14] , \chs_in_f[1][DATA][13] ,
         \chs_in_f[1][DATA][12] , \chs_in_f[1][DATA][11] ,
         \chs_in_f[1][DATA][10] , \chs_in_f[1][DATA][9] ,
         \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] ,
         \chs_in_f[1][DATA][6] , \chs_in_f[1][DATA][5] ,
         \chs_in_f[1][DATA][4] , \chs_in_f[1][DATA][3] ,
         \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] ,
         \chs_in_f[1][DATA][0] , \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] ,
         \chs_in_f[0][DATA][33] , \chs_in_f[0][DATA][32] ,
         \chs_in_f[0][DATA][31] , \chs_in_f[0][DATA][30] ,
         \chs_in_f[0][DATA][29] , \chs_in_f[0][DATA][28] ,
         \chs_in_f[0][DATA][27] , \chs_in_f[0][DATA][26] ,
         \chs_in_f[0][DATA][25] , \chs_in_f[0][DATA][24] ,
         \chs_in_f[0][DATA][23] , \chs_in_f[0][DATA][22] ,
         \chs_in_f[0][DATA][21] , \chs_in_f[0][DATA][20] ,
         \chs_in_f[0][DATA][19] , \chs_in_f[0][DATA][18] ,
         \chs_in_f[0][DATA][17] , \chs_in_f[0][DATA][16] ,
         \chs_in_f[0][DATA][15] , \chs_in_f[0][DATA][14] ,
         \chs_in_f[0][DATA][13] , \chs_in_f[0][DATA][12] ,
         \chs_in_f[0][DATA][11] , \chs_in_f[0][DATA][10] ,
         \chs_in_f[0][DATA][9] , \chs_in_f[0][DATA][8] ,
         \chs_in_f[0][DATA][7] , \chs_in_f[0][DATA][6] ,
         \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] ,
         \chs_in_f[0][DATA][3] , \chs_in_f[0][DATA][2] ,
         \chs_in_f[0][DATA][1] , \chs_in_f[0][DATA][0] , \chs_in_b[4][ACK] ,
         \chs_in_b[3][ACK] , \chs_in_b[2][ACK] , \chs_in_b[1][ACK] ,
         \chs_in_b[0][ACK] , \switch_sel[4][4] , \switch_sel[4][3] ,
         \switch_sel[4][2] , \switch_sel[4][1] , \switch_sel[4][0] ,
         \switch_sel[3][4] , \switch_sel[3][3] , \switch_sel[3][2] ,
         \switch_sel[3][1] , \switch_sel[3][0] , \switch_sel[2][4] ,
         \switch_sel[2][3] , \switch_sel[2][2] , \switch_sel[2][1] ,
         \switch_sel[2][0] , \switch_sel[1][4] , \switch_sel[1][3] ,
         \switch_sel[1][2] , \switch_sel[1][1] , \switch_sel[1][0] ,
         \switch_sel[0][4] , \switch_sel[0][3] , \switch_sel[0][2] ,
         \switch_sel[0][1] , \switch_sel[0][0] , n2, n3;

  channel_latch_1_xxxxxxxxx_25 north_in_latch ( .preset(n3), .left_in({
        \north_in_f[REQ] , \north_in_f[DATA][34] , \north_in_f[DATA][33] , 
        \north_in_f[DATA][32] , \north_in_f[DATA][31] , \north_in_f[DATA][30] , 
        \north_in_f[DATA][29] , \north_in_f[DATA][28] , \north_in_f[DATA][27] , 
        \north_in_f[DATA][26] , \north_in_f[DATA][25] , \north_in_f[DATA][24] , 
        \north_in_f[DATA][23] , \north_in_f[DATA][22] , \north_in_f[DATA][21] , 
        \north_in_f[DATA][20] , \north_in_f[DATA][19] , \north_in_f[DATA][18] , 
        \north_in_f[DATA][17] , \north_in_f[DATA][16] , \north_in_f[DATA][15] , 
        \north_in_f[DATA][14] , \north_in_f[DATA][13] , \north_in_f[DATA][12] , 
        \north_in_f[DATA][11] , \north_in_f[DATA][10] , \north_in_f[DATA][9] , 
        \north_in_f[DATA][8] , \north_in_f[DATA][7] , \north_in_f[DATA][6] , 
        \north_in_f[DATA][5] , \north_in_f[DATA][4] , \north_in_f[DATA][3] , 
        \north_in_f[DATA][2] , \north_in_f[DATA][1] , \north_in_f[DATA][0] }), 
        .left_out(\north_in_b[ACK] ), .right_out({\north_hpu_f[REQ] , 
        \north_hpu_f[DATA][34] , \north_hpu_f[DATA][33] , 
        \north_hpu_f[DATA][32] , \north_hpu_f[DATA][31] , 
        \north_hpu_f[DATA][30] , \north_hpu_f[DATA][29] , 
        \north_hpu_f[DATA][28] , \north_hpu_f[DATA][27] , 
        \north_hpu_f[DATA][26] , \north_hpu_f[DATA][25] , 
        \north_hpu_f[DATA][24] , \north_hpu_f[DATA][23] , 
        \north_hpu_f[DATA][22] , \north_hpu_f[DATA][21] , 
        \north_hpu_f[DATA][20] , \north_hpu_f[DATA][19] , 
        \north_hpu_f[DATA][18] , \north_hpu_f[DATA][17] , 
        \north_hpu_f[DATA][16] , \north_hpu_f[DATA][15] , 
        \north_hpu_f[DATA][14] , \north_hpu_f[DATA][13] , 
        \north_hpu_f[DATA][12] , \north_hpu_f[DATA][11] , 
        \north_hpu_f[DATA][10] , \north_hpu_f[DATA][9] , 
        \north_hpu_f[DATA][8] , \north_hpu_f[DATA][7] , \north_hpu_f[DATA][6] , 
        \north_hpu_f[DATA][5] , \north_hpu_f[DATA][4] , \north_hpu_f[DATA][3] , 
        \north_hpu_f[DATA][2] , \north_hpu_f[DATA][1] , \north_hpu_f[DATA][0] }), .right_in(\north_hpu_b[ACK] ) );
  channel_latch_1_xxxxxxxxx_24 south_in_latch ( .preset(n3), .left_in({
        \south_in_f[REQ] , \south_in_f[DATA][34] , \south_in_f[DATA][33] , 
        \south_in_f[DATA][32] , \south_in_f[DATA][31] , \south_in_f[DATA][30] , 
        \south_in_f[DATA][29] , \south_in_f[DATA][28] , \south_in_f[DATA][27] , 
        \south_in_f[DATA][26] , \south_in_f[DATA][25] , \south_in_f[DATA][24] , 
        \south_in_f[DATA][23] , \south_in_f[DATA][22] , \south_in_f[DATA][21] , 
        \south_in_f[DATA][20] , \south_in_f[DATA][19] , \south_in_f[DATA][18] , 
        \south_in_f[DATA][17] , \south_in_f[DATA][16] , \south_in_f[DATA][15] , 
        \south_in_f[DATA][14] , \south_in_f[DATA][13] , \south_in_f[DATA][12] , 
        \south_in_f[DATA][11] , \south_in_f[DATA][10] , \south_in_f[DATA][9] , 
        \south_in_f[DATA][8] , \south_in_f[DATA][7] , \south_in_f[DATA][6] , 
        \south_in_f[DATA][5] , \south_in_f[DATA][4] , \south_in_f[DATA][3] , 
        \south_in_f[DATA][2] , \south_in_f[DATA][1] , \south_in_f[DATA][0] }), 
        .left_out(\south_in_b[ACK] ), .right_out({\south_hpu_f[REQ] , 
        \south_hpu_f[DATA][34] , \south_hpu_f[DATA][33] , 
        \south_hpu_f[DATA][32] , \south_hpu_f[DATA][31] , 
        \south_hpu_f[DATA][30] , \south_hpu_f[DATA][29] , 
        \south_hpu_f[DATA][28] , \south_hpu_f[DATA][27] , 
        \south_hpu_f[DATA][26] , \south_hpu_f[DATA][25] , 
        \south_hpu_f[DATA][24] , \south_hpu_f[DATA][23] , 
        \south_hpu_f[DATA][22] , \south_hpu_f[DATA][21] , 
        \south_hpu_f[DATA][20] , \south_hpu_f[DATA][19] , 
        \south_hpu_f[DATA][18] , \south_hpu_f[DATA][17] , 
        \south_hpu_f[DATA][16] , \south_hpu_f[DATA][15] , 
        \south_hpu_f[DATA][14] , \south_hpu_f[DATA][13] , 
        \south_hpu_f[DATA][12] , \south_hpu_f[DATA][11] , 
        \south_hpu_f[DATA][10] , \south_hpu_f[DATA][9] , 
        \south_hpu_f[DATA][8] , \south_hpu_f[DATA][7] , \south_hpu_f[DATA][6] , 
        \south_hpu_f[DATA][5] , \south_hpu_f[DATA][4] , \south_hpu_f[DATA][3] , 
        \south_hpu_f[DATA][2] , \south_hpu_f[DATA][1] , \south_hpu_f[DATA][0] }), .right_in(\south_hpu_b[ACK] ) );
  channel_latch_1_xxxxxxxxx_23 east_in_latch ( .preset(n3), .left_in({
        \east_in_f[REQ] , \east_in_f[DATA][34] , \east_in_f[DATA][33] , 
        \east_in_f[DATA][32] , \east_in_f[DATA][31] , \east_in_f[DATA][30] , 
        \east_in_f[DATA][29] , \east_in_f[DATA][28] , \east_in_f[DATA][27] , 
        \east_in_f[DATA][26] , \east_in_f[DATA][25] , \east_in_f[DATA][24] , 
        \east_in_f[DATA][23] , \east_in_f[DATA][22] , \east_in_f[DATA][21] , 
        \east_in_f[DATA][20] , \east_in_f[DATA][19] , \east_in_f[DATA][18] , 
        \east_in_f[DATA][17] , \east_in_f[DATA][16] , \east_in_f[DATA][15] , 
        \east_in_f[DATA][14] , \east_in_f[DATA][13] , \east_in_f[DATA][12] , 
        \east_in_f[DATA][11] , \east_in_f[DATA][10] , \east_in_f[DATA][9] , 
        \east_in_f[DATA][8] , \east_in_f[DATA][7] , \east_in_f[DATA][6] , 
        \east_in_f[DATA][5] , \east_in_f[DATA][4] , \east_in_f[DATA][3] , 
        \east_in_f[DATA][2] , \east_in_f[DATA][1] , \east_in_f[DATA][0] }), 
        .left_out(\east_in_b[ACK] ), .right_out({\east_hpu_f[REQ] , 
        \east_hpu_f[DATA][34] , \east_hpu_f[DATA][33] , \east_hpu_f[DATA][32] , 
        \east_hpu_f[DATA][31] , \east_hpu_f[DATA][30] , \east_hpu_f[DATA][29] , 
        \east_hpu_f[DATA][28] , \east_hpu_f[DATA][27] , \east_hpu_f[DATA][26] , 
        \east_hpu_f[DATA][25] , \east_hpu_f[DATA][24] , \east_hpu_f[DATA][23] , 
        \east_hpu_f[DATA][22] , \east_hpu_f[DATA][21] , \east_hpu_f[DATA][20] , 
        \east_hpu_f[DATA][19] , \east_hpu_f[DATA][18] , \east_hpu_f[DATA][17] , 
        \east_hpu_f[DATA][16] , \east_hpu_f[DATA][15] , \east_hpu_f[DATA][14] , 
        \east_hpu_f[DATA][13] , \east_hpu_f[DATA][12] , \east_hpu_f[DATA][11] , 
        \east_hpu_f[DATA][10] , \east_hpu_f[DATA][9] , \east_hpu_f[DATA][8] , 
        \east_hpu_f[DATA][7] , \east_hpu_f[DATA][6] , \east_hpu_f[DATA][5] , 
        \east_hpu_f[DATA][4] , \east_hpu_f[DATA][3] , \east_hpu_f[DATA][2] , 
        \east_hpu_f[DATA][1] , \east_hpu_f[DATA][0] }), .right_in(
        \east_hpu_b[ACK] ) );
  channel_latch_1_xxxxxxxxx_22 west_in_latch ( .preset(n3), .left_in({
        \west_in_f[REQ] , \west_in_f[DATA][34] , \west_in_f[DATA][33] , 
        \west_in_f[DATA][32] , \west_in_f[DATA][31] , \west_in_f[DATA][30] , 
        \west_in_f[DATA][29] , \west_in_f[DATA][28] , \west_in_f[DATA][27] , 
        \west_in_f[DATA][26] , \west_in_f[DATA][25] , \west_in_f[DATA][24] , 
        \west_in_f[DATA][23] , \west_in_f[DATA][22] , \west_in_f[DATA][21] , 
        \west_in_f[DATA][20] , \west_in_f[DATA][19] , \west_in_f[DATA][18] , 
        \west_in_f[DATA][17] , \west_in_f[DATA][16] , \west_in_f[DATA][15] , 
        \west_in_f[DATA][14] , \west_in_f[DATA][13] , \west_in_f[DATA][12] , 
        \west_in_f[DATA][11] , \west_in_f[DATA][10] , \west_in_f[DATA][9] , 
        \west_in_f[DATA][8] , \west_in_f[DATA][7] , \west_in_f[DATA][6] , 
        \west_in_f[DATA][5] , \west_in_f[DATA][4] , \west_in_f[DATA][3] , 
        \west_in_f[DATA][2] , \west_in_f[DATA][1] , \west_in_f[DATA][0] }), 
        .left_out(\west_in_b[ACK] ), .right_out({\west_hpu_f[REQ] , 
        \west_hpu_f[DATA][34] , \west_hpu_f[DATA][33] , \west_hpu_f[DATA][32] , 
        \west_hpu_f[DATA][31] , \west_hpu_f[DATA][30] , \west_hpu_f[DATA][29] , 
        \west_hpu_f[DATA][28] , \west_hpu_f[DATA][27] , \west_hpu_f[DATA][26] , 
        \west_hpu_f[DATA][25] , \west_hpu_f[DATA][24] , \west_hpu_f[DATA][23] , 
        \west_hpu_f[DATA][22] , \west_hpu_f[DATA][21] , \west_hpu_f[DATA][20] , 
        \west_hpu_f[DATA][19] , \west_hpu_f[DATA][18] , \west_hpu_f[DATA][17] , 
        \west_hpu_f[DATA][16] , \west_hpu_f[DATA][15] , \west_hpu_f[DATA][14] , 
        \west_hpu_f[DATA][13] , \west_hpu_f[DATA][12] , \west_hpu_f[DATA][11] , 
        \west_hpu_f[DATA][10] , \west_hpu_f[DATA][9] , \west_hpu_f[DATA][8] , 
        \west_hpu_f[DATA][7] , \west_hpu_f[DATA][6] , \west_hpu_f[DATA][5] , 
        \west_hpu_f[DATA][4] , \west_hpu_f[DATA][3] , \west_hpu_f[DATA][2] , 
        \west_hpu_f[DATA][1] , \west_hpu_f[DATA][0] }), .right_in(
        \west_hpu_b[ACK] ) );
  channel_latch_1_xxxxxxxxx_21 resource_in_latch ( .preset(n3), .left_in({
        \resource_in_f[REQ] , \resource_in_f[DATA][34] , 
        \resource_in_f[DATA][33] , \resource_in_f[DATA][32] , 
        \resource_in_f[DATA][31] , \resource_in_f[DATA][30] , 
        \resource_in_f[DATA][29] , \resource_in_f[DATA][28] , 
        \resource_in_f[DATA][27] , \resource_in_f[DATA][26] , 
        \resource_in_f[DATA][25] , \resource_in_f[DATA][24] , 
        \resource_in_f[DATA][23] , \resource_in_f[DATA][22] , 
        \resource_in_f[DATA][21] , \resource_in_f[DATA][20] , 
        \resource_in_f[DATA][19] , \resource_in_f[DATA][18] , 
        \resource_in_f[DATA][17] , \resource_in_f[DATA][16] , 
        \resource_in_f[DATA][15] , \resource_in_f[DATA][14] , 
        \resource_in_f[DATA][13] , \resource_in_f[DATA][12] , 
        \resource_in_f[DATA][11] , \resource_in_f[DATA][10] , 
        \resource_in_f[DATA][9] , \resource_in_f[DATA][8] , 
        \resource_in_f[DATA][7] , \resource_in_f[DATA][6] , 
        \resource_in_f[DATA][5] , \resource_in_f[DATA][4] , 
        \resource_in_f[DATA][3] , \resource_in_f[DATA][2] , 
        \resource_in_f[DATA][1] , \resource_in_f[DATA][0] }), .left_out(
        \resource_in_b[ACK] ), .right_out({\resource_hpu_f[REQ] , 
        \resource_hpu_f[DATA][34] , \resource_hpu_f[DATA][33] , 
        \resource_hpu_f[DATA][32] , \resource_hpu_f[DATA][31] , 
        \resource_hpu_f[DATA][30] , \resource_hpu_f[DATA][29] , 
        \resource_hpu_f[DATA][28] , \resource_hpu_f[DATA][27] , 
        \resource_hpu_f[DATA][26] , \resource_hpu_f[DATA][25] , 
        \resource_hpu_f[DATA][24] , \resource_hpu_f[DATA][23] , 
        \resource_hpu_f[DATA][22] , \resource_hpu_f[DATA][21] , 
        \resource_hpu_f[DATA][20] , \resource_hpu_f[DATA][19] , 
        \resource_hpu_f[DATA][18] , \resource_hpu_f[DATA][17] , 
        \resource_hpu_f[DATA][16] , \resource_hpu_f[DATA][15] , 
        \resource_hpu_f[DATA][14] , \resource_hpu_f[DATA][13] , 
        \resource_hpu_f[DATA][12] , \resource_hpu_f[DATA][11] , 
        \resource_hpu_f[DATA][10] , \resource_hpu_f[DATA][9] , 
        \resource_hpu_f[DATA][8] , \resource_hpu_f[DATA][7] , 
        \resource_hpu_f[DATA][6] , \resource_hpu_f[DATA][5] , 
        \resource_hpu_f[DATA][4] , \resource_hpu_f[DATA][3] , 
        \resource_hpu_f[DATA][2] , \resource_hpu_f[DATA][1] , 
        \resource_hpu_f[DATA][0] }), .right_in(\resource_hpu_b[ACK] ) );
  hpu_0_0_1 north_hpu ( .preset(n2), .chan_in_f({\north_hpu_f[REQ] , 
        \north_hpu_f[DATA][34] , \north_hpu_f[DATA][33] , 
        \north_hpu_f[DATA][32] , \north_hpu_f[DATA][31] , 
        \north_hpu_f[DATA][30] , \north_hpu_f[DATA][29] , 
        \north_hpu_f[DATA][28] , \north_hpu_f[DATA][27] , 
        \north_hpu_f[DATA][26] , \north_hpu_f[DATA][25] , 
        \north_hpu_f[DATA][24] , \north_hpu_f[DATA][23] , 
        \north_hpu_f[DATA][22] , \north_hpu_f[DATA][21] , 
        \north_hpu_f[DATA][20] , \north_hpu_f[DATA][19] , 
        \north_hpu_f[DATA][18] , \north_hpu_f[DATA][17] , 
        \north_hpu_f[DATA][16] , \north_hpu_f[DATA][15] , 
        \north_hpu_f[DATA][14] , \north_hpu_f[DATA][13] , 
        \north_hpu_f[DATA][12] , \north_hpu_f[DATA][11] , 
        \north_hpu_f[DATA][10] , \north_hpu_f[DATA][9] , 
        \north_hpu_f[DATA][8] , \north_hpu_f[DATA][7] , \north_hpu_f[DATA][6] , 
        \north_hpu_f[DATA][5] , \north_hpu_f[DATA][4] , \north_hpu_f[DATA][3] , 
        \north_hpu_f[DATA][2] , \north_hpu_f[DATA][1] , \north_hpu_f[DATA][0] }), .chan_in_b(\north_hpu_b[ACK] ), .chan_out_f({\chs_in_f[0][REQ] , 
        \chs_in_f[0][DATA][34] , \chs_in_f[0][DATA][33] , 
        \chs_in_f[0][DATA][32] , \chs_in_f[0][DATA][31] , 
        \chs_in_f[0][DATA][30] , \chs_in_f[0][DATA][29] , 
        \chs_in_f[0][DATA][28] , \chs_in_f[0][DATA][27] , 
        \chs_in_f[0][DATA][26] , \chs_in_f[0][DATA][25] , 
        \chs_in_f[0][DATA][24] , \chs_in_f[0][DATA][23] , 
        \chs_in_f[0][DATA][22] , \chs_in_f[0][DATA][21] , 
        \chs_in_f[0][DATA][20] , \chs_in_f[0][DATA][19] , 
        \chs_in_f[0][DATA][18] , \chs_in_f[0][DATA][17] , 
        \chs_in_f[0][DATA][16] , \chs_in_f[0][DATA][15] , 
        \chs_in_f[0][DATA][14] , \chs_in_f[0][DATA][13] , 
        \chs_in_f[0][DATA][12] , \chs_in_f[0][DATA][11] , 
        \chs_in_f[0][DATA][10] , \chs_in_f[0][DATA][9] , 
        \chs_in_f[0][DATA][8] , \chs_in_f[0][DATA][7] , \chs_in_f[0][DATA][6] , 
        \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] , \chs_in_f[0][DATA][3] , 
        \chs_in_f[0][DATA][2] , \chs_in_f[0][DATA][1] , \chs_in_f[0][DATA][0] }), .chan_out_b(\chs_in_b[0][ACK] ), .sel({\switch_sel[0][4] , 
        \switch_sel[0][3] , \switch_sel[0][2] , \switch_sel[0][1] , 
        \switch_sel[0][0] }) );
  hpu_0_2_1 south_hpu ( .preset(n2), .chan_in_f({\south_hpu_f[REQ] , 
        \south_hpu_f[DATA][34] , \south_hpu_f[DATA][33] , 
        \south_hpu_f[DATA][32] , \south_hpu_f[DATA][31] , 
        \south_hpu_f[DATA][30] , \south_hpu_f[DATA][29] , 
        \south_hpu_f[DATA][28] , \south_hpu_f[DATA][27] , 
        \south_hpu_f[DATA][26] , \south_hpu_f[DATA][25] , 
        \south_hpu_f[DATA][24] , \south_hpu_f[DATA][23] , 
        \south_hpu_f[DATA][22] , \south_hpu_f[DATA][21] , 
        \south_hpu_f[DATA][20] , \south_hpu_f[DATA][19] , 
        \south_hpu_f[DATA][18] , \south_hpu_f[DATA][17] , 
        \south_hpu_f[DATA][16] , \south_hpu_f[DATA][15] , 
        \south_hpu_f[DATA][14] , \south_hpu_f[DATA][13] , 
        \south_hpu_f[DATA][12] , \south_hpu_f[DATA][11] , 
        \south_hpu_f[DATA][10] , \south_hpu_f[DATA][9] , 
        \south_hpu_f[DATA][8] , \south_hpu_f[DATA][7] , \south_hpu_f[DATA][6] , 
        \south_hpu_f[DATA][5] , \south_hpu_f[DATA][4] , \south_hpu_f[DATA][3] , 
        \south_hpu_f[DATA][2] , \south_hpu_f[DATA][1] , \south_hpu_f[DATA][0] }), .chan_in_b(\south_hpu_b[ACK] ), .chan_out_f({\chs_in_f[2][REQ] , 
        \chs_in_f[2][DATA][34] , \chs_in_f[2][DATA][33] , 
        \chs_in_f[2][DATA][32] , \chs_in_f[2][DATA][31] , 
        \chs_in_f[2][DATA][30] , \chs_in_f[2][DATA][29] , 
        \chs_in_f[2][DATA][28] , \chs_in_f[2][DATA][27] , 
        \chs_in_f[2][DATA][26] , \chs_in_f[2][DATA][25] , 
        \chs_in_f[2][DATA][24] , \chs_in_f[2][DATA][23] , 
        \chs_in_f[2][DATA][22] , \chs_in_f[2][DATA][21] , 
        \chs_in_f[2][DATA][20] , \chs_in_f[2][DATA][19] , 
        \chs_in_f[2][DATA][18] , \chs_in_f[2][DATA][17] , 
        \chs_in_f[2][DATA][16] , \chs_in_f[2][DATA][15] , 
        \chs_in_f[2][DATA][14] , \chs_in_f[2][DATA][13] , 
        \chs_in_f[2][DATA][12] , \chs_in_f[2][DATA][11] , 
        \chs_in_f[2][DATA][10] , \chs_in_f[2][DATA][9] , 
        \chs_in_f[2][DATA][8] , \chs_in_f[2][DATA][7] , \chs_in_f[2][DATA][6] , 
        \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] , \chs_in_f[2][DATA][3] , 
        \chs_in_f[2][DATA][2] , \chs_in_f[2][DATA][1] , \chs_in_f[2][DATA][0] }), .chan_out_b(\chs_in_b[2][ACK] ), .sel({\switch_sel[2][4] , 
        \switch_sel[2][3] , \switch_sel[2][2] , \switch_sel[2][1] , 
        \switch_sel[2][0] }) );
  hpu_0_1_1 east_hpu ( .preset(n2), .chan_in_f({\east_hpu_f[REQ] , 
        \east_hpu_f[DATA][34] , \east_hpu_f[DATA][33] , \east_hpu_f[DATA][32] , 
        \east_hpu_f[DATA][31] , \east_hpu_f[DATA][30] , \east_hpu_f[DATA][29] , 
        \east_hpu_f[DATA][28] , \east_hpu_f[DATA][27] , \east_hpu_f[DATA][26] , 
        \east_hpu_f[DATA][25] , \east_hpu_f[DATA][24] , \east_hpu_f[DATA][23] , 
        \east_hpu_f[DATA][22] , \east_hpu_f[DATA][21] , \east_hpu_f[DATA][20] , 
        \east_hpu_f[DATA][19] , \east_hpu_f[DATA][18] , \east_hpu_f[DATA][17] , 
        \east_hpu_f[DATA][16] , \east_hpu_f[DATA][15] , \east_hpu_f[DATA][14] , 
        \east_hpu_f[DATA][13] , \east_hpu_f[DATA][12] , \east_hpu_f[DATA][11] , 
        \east_hpu_f[DATA][10] , \east_hpu_f[DATA][9] , \east_hpu_f[DATA][8] , 
        \east_hpu_f[DATA][7] , \east_hpu_f[DATA][6] , \east_hpu_f[DATA][5] , 
        \east_hpu_f[DATA][4] , \east_hpu_f[DATA][3] , \east_hpu_f[DATA][2] , 
        \east_hpu_f[DATA][1] , \east_hpu_f[DATA][0] }), .chan_in_b(
        \east_hpu_b[ACK] ), .chan_out_f({\chs_in_f[1][REQ] , 
        \chs_in_f[1][DATA][34] , \chs_in_f[1][DATA][33] , 
        \chs_in_f[1][DATA][32] , \chs_in_f[1][DATA][31] , 
        \chs_in_f[1][DATA][30] , \chs_in_f[1][DATA][29] , 
        \chs_in_f[1][DATA][28] , \chs_in_f[1][DATA][27] , 
        \chs_in_f[1][DATA][26] , \chs_in_f[1][DATA][25] , 
        \chs_in_f[1][DATA][24] , \chs_in_f[1][DATA][23] , 
        \chs_in_f[1][DATA][22] , \chs_in_f[1][DATA][21] , 
        \chs_in_f[1][DATA][20] , \chs_in_f[1][DATA][19] , 
        \chs_in_f[1][DATA][18] , \chs_in_f[1][DATA][17] , 
        \chs_in_f[1][DATA][16] , \chs_in_f[1][DATA][15] , 
        \chs_in_f[1][DATA][14] , \chs_in_f[1][DATA][13] , 
        \chs_in_f[1][DATA][12] , \chs_in_f[1][DATA][11] , 
        \chs_in_f[1][DATA][10] , \chs_in_f[1][DATA][9] , 
        \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] , \chs_in_f[1][DATA][6] , 
        \chs_in_f[1][DATA][5] , \chs_in_f[1][DATA][4] , \chs_in_f[1][DATA][3] , 
        \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] , \chs_in_f[1][DATA][0] }), .chan_out_b(\chs_in_b[1][ACK] ), .sel({\switch_sel[1][4] , 
        \switch_sel[1][3] , \switch_sel[1][2] , \switch_sel[1][1] , 
        \switch_sel[1][0] }) );
  hpu_0_3_1 west_hpu ( .preset(n2), .chan_in_f({\west_hpu_f[REQ] , 
        \west_hpu_f[DATA][34] , \west_hpu_f[DATA][33] , \west_hpu_f[DATA][32] , 
        \west_hpu_f[DATA][31] , \west_hpu_f[DATA][30] , \west_hpu_f[DATA][29] , 
        \west_hpu_f[DATA][28] , \west_hpu_f[DATA][27] , \west_hpu_f[DATA][26] , 
        \west_hpu_f[DATA][25] , \west_hpu_f[DATA][24] , \west_hpu_f[DATA][23] , 
        \west_hpu_f[DATA][22] , \west_hpu_f[DATA][21] , \west_hpu_f[DATA][20] , 
        \west_hpu_f[DATA][19] , \west_hpu_f[DATA][18] , \west_hpu_f[DATA][17] , 
        \west_hpu_f[DATA][16] , \west_hpu_f[DATA][15] , \west_hpu_f[DATA][14] , 
        \west_hpu_f[DATA][13] , \west_hpu_f[DATA][12] , \west_hpu_f[DATA][11] , 
        \west_hpu_f[DATA][10] , \west_hpu_f[DATA][9] , \west_hpu_f[DATA][8] , 
        \west_hpu_f[DATA][7] , \west_hpu_f[DATA][6] , \west_hpu_f[DATA][5] , 
        \west_hpu_f[DATA][4] , \west_hpu_f[DATA][3] , \west_hpu_f[DATA][2] , 
        \west_hpu_f[DATA][1] , \west_hpu_f[DATA][0] }), .chan_in_b(
        \west_hpu_b[ACK] ), .chan_out_f({\chs_in_f[3][REQ] , 
        \chs_in_f[3][DATA][34] , \chs_in_f[3][DATA][33] , 
        \chs_in_f[3][DATA][32] , \chs_in_f[3][DATA][31] , 
        \chs_in_f[3][DATA][30] , \chs_in_f[3][DATA][29] , 
        \chs_in_f[3][DATA][28] , \chs_in_f[3][DATA][27] , 
        \chs_in_f[3][DATA][26] , \chs_in_f[3][DATA][25] , 
        \chs_in_f[3][DATA][24] , \chs_in_f[3][DATA][23] , 
        \chs_in_f[3][DATA][22] , \chs_in_f[3][DATA][21] , 
        \chs_in_f[3][DATA][20] , \chs_in_f[3][DATA][19] , 
        \chs_in_f[3][DATA][18] , \chs_in_f[3][DATA][17] , 
        \chs_in_f[3][DATA][16] , \chs_in_f[3][DATA][15] , 
        \chs_in_f[3][DATA][14] , \chs_in_f[3][DATA][13] , 
        \chs_in_f[3][DATA][12] , \chs_in_f[3][DATA][11] , 
        \chs_in_f[3][DATA][10] , \chs_in_f[3][DATA][9] , 
        \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] , \chs_in_f[3][DATA][6] , 
        \chs_in_f[3][DATA][5] , \chs_in_f[3][DATA][4] , \chs_in_f[3][DATA][3] , 
        \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] , \chs_in_f[3][DATA][0] }), .chan_out_b(\chs_in_b[3][ACK] ), .sel({\switch_sel[3][4] , 
        \switch_sel[3][3] , \switch_sel[3][2] , \switch_sel[3][1] , 
        \switch_sel[3][0] }) );
  hpu_1_x_1 resource_hpu ( .preset(n2), .chan_in_f({\resource_hpu_f[REQ] , 
        \resource_hpu_f[DATA][34] , \resource_hpu_f[DATA][33] , 
        \resource_hpu_f[DATA][32] , \resource_hpu_f[DATA][31] , 
        \resource_hpu_f[DATA][30] , \resource_hpu_f[DATA][29] , 
        \resource_hpu_f[DATA][28] , \resource_hpu_f[DATA][27] , 
        \resource_hpu_f[DATA][26] , \resource_hpu_f[DATA][25] , 
        \resource_hpu_f[DATA][24] , \resource_hpu_f[DATA][23] , 
        \resource_hpu_f[DATA][22] , \resource_hpu_f[DATA][21] , 
        \resource_hpu_f[DATA][20] , \resource_hpu_f[DATA][19] , 
        \resource_hpu_f[DATA][18] , \resource_hpu_f[DATA][17] , 
        \resource_hpu_f[DATA][16] , \resource_hpu_f[DATA][15] , 
        \resource_hpu_f[DATA][14] , \resource_hpu_f[DATA][13] , 
        \resource_hpu_f[DATA][12] , \resource_hpu_f[DATA][11] , 
        \resource_hpu_f[DATA][10] , \resource_hpu_f[DATA][9] , 
        \resource_hpu_f[DATA][8] , \resource_hpu_f[DATA][7] , 
        \resource_hpu_f[DATA][6] , \resource_hpu_f[DATA][5] , 
        \resource_hpu_f[DATA][4] , \resource_hpu_f[DATA][3] , 
        \resource_hpu_f[DATA][2] , \resource_hpu_f[DATA][1] , 
        \resource_hpu_f[DATA][0] }), .chan_in_b(\resource_hpu_b[ACK] ), 
        .chan_out_f({\chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] , 
        \chs_in_f[4][DATA][33] , \chs_in_f[4][DATA][32] , 
        \chs_in_f[4][DATA][31] , \chs_in_f[4][DATA][30] , 
        \chs_in_f[4][DATA][29] , \chs_in_f[4][DATA][28] , 
        \chs_in_f[4][DATA][27] , \chs_in_f[4][DATA][26] , 
        \chs_in_f[4][DATA][25] , \chs_in_f[4][DATA][24] , 
        \chs_in_f[4][DATA][23] , \chs_in_f[4][DATA][22] , 
        \chs_in_f[4][DATA][21] , \chs_in_f[4][DATA][20] , 
        \chs_in_f[4][DATA][19] , \chs_in_f[4][DATA][18] , 
        \chs_in_f[4][DATA][17] , \chs_in_f[4][DATA][16] , 
        \chs_in_f[4][DATA][15] , \chs_in_f[4][DATA][14] , 
        \chs_in_f[4][DATA][13] , \chs_in_f[4][DATA][12] , 
        \chs_in_f[4][DATA][11] , \chs_in_f[4][DATA][10] , 
        \chs_in_f[4][DATA][9] , \chs_in_f[4][DATA][8] , \chs_in_f[4][DATA][7] , 
        \chs_in_f[4][DATA][6] , \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] , 
        \chs_in_f[4][DATA][3] , \chs_in_f[4][DATA][2] , \chs_in_f[4][DATA][1] , 
        \chs_in_f[4][DATA][0] }), .chan_out_b(\chs_in_b[4][ACK] ), .sel({
        \switch_sel[4][4] , \switch_sel[4][3] , \switch_sel[4][2] , 
        \switch_sel[4][1] , \switch_sel[4][0] }) );
  crossbar_stage_1 xbar_with_latches ( .preset(n3), .switch_sel({1'b0, 
        \switch_sel[4][3] , \switch_sel[4][2] , \switch_sel[4][1] , 
        \switch_sel[4][0] , \switch_sel[3][4] , 1'b0, \switch_sel[3][2] , 
        \switch_sel[3][1] , \switch_sel[3][0] , \switch_sel[2][4] , 
        \switch_sel[2][3] , 1'b0, \switch_sel[2][1] , \switch_sel[2][0] , 
        \switch_sel[1][4] , \switch_sel[1][3] , \switch_sel[1][2] , 1'b0, 
        \switch_sel[1][0] , \switch_sel[0][4] , \switch_sel[0][3] , 
        \switch_sel[0][2] , \switch_sel[0][1] , 1'b0}), .chs_in_f({
        \chs_in_f[4][REQ] , \chs_in_f[4][DATA][34] , \chs_in_f[4][DATA][33] , 
        \chs_in_f[4][DATA][32] , \chs_in_f[4][DATA][31] , 
        \chs_in_f[4][DATA][30] , \chs_in_f[4][DATA][29] , 
        \chs_in_f[4][DATA][28] , \chs_in_f[4][DATA][27] , 
        \chs_in_f[4][DATA][26] , \chs_in_f[4][DATA][25] , 
        \chs_in_f[4][DATA][24] , \chs_in_f[4][DATA][23] , 
        \chs_in_f[4][DATA][22] , \chs_in_f[4][DATA][21] , 
        \chs_in_f[4][DATA][20] , \chs_in_f[4][DATA][19] , 
        \chs_in_f[4][DATA][18] , \chs_in_f[4][DATA][17] , 
        \chs_in_f[4][DATA][16] , \chs_in_f[4][DATA][15] , 
        \chs_in_f[4][DATA][14] , \chs_in_f[4][DATA][13] , 
        \chs_in_f[4][DATA][12] , \chs_in_f[4][DATA][11] , 
        \chs_in_f[4][DATA][10] , \chs_in_f[4][DATA][9] , 
        \chs_in_f[4][DATA][8] , \chs_in_f[4][DATA][7] , \chs_in_f[4][DATA][6] , 
        \chs_in_f[4][DATA][5] , \chs_in_f[4][DATA][4] , \chs_in_f[4][DATA][3] , 
        \chs_in_f[4][DATA][2] , \chs_in_f[4][DATA][1] , \chs_in_f[4][DATA][0] , 
        \chs_in_f[3][REQ] , \chs_in_f[3][DATA][34] , \chs_in_f[3][DATA][33] , 
        \chs_in_f[3][DATA][32] , \chs_in_f[3][DATA][31] , 
        \chs_in_f[3][DATA][30] , \chs_in_f[3][DATA][29] , 
        \chs_in_f[3][DATA][28] , \chs_in_f[3][DATA][27] , 
        \chs_in_f[3][DATA][26] , \chs_in_f[3][DATA][25] , 
        \chs_in_f[3][DATA][24] , \chs_in_f[3][DATA][23] , 
        \chs_in_f[3][DATA][22] , \chs_in_f[3][DATA][21] , 
        \chs_in_f[3][DATA][20] , \chs_in_f[3][DATA][19] , 
        \chs_in_f[3][DATA][18] , \chs_in_f[3][DATA][17] , 
        \chs_in_f[3][DATA][16] , \chs_in_f[3][DATA][15] , 
        \chs_in_f[3][DATA][14] , \chs_in_f[3][DATA][13] , 
        \chs_in_f[3][DATA][12] , \chs_in_f[3][DATA][11] , 
        \chs_in_f[3][DATA][10] , \chs_in_f[3][DATA][9] , 
        \chs_in_f[3][DATA][8] , \chs_in_f[3][DATA][7] , \chs_in_f[3][DATA][6] , 
        \chs_in_f[3][DATA][5] , \chs_in_f[3][DATA][4] , \chs_in_f[3][DATA][3] , 
        \chs_in_f[3][DATA][2] , \chs_in_f[3][DATA][1] , \chs_in_f[3][DATA][0] , 
        \chs_in_f[2][REQ] , \chs_in_f[2][DATA][34] , \chs_in_f[2][DATA][33] , 
        \chs_in_f[2][DATA][32] , \chs_in_f[2][DATA][31] , 
        \chs_in_f[2][DATA][30] , \chs_in_f[2][DATA][29] , 
        \chs_in_f[2][DATA][28] , \chs_in_f[2][DATA][27] , 
        \chs_in_f[2][DATA][26] , \chs_in_f[2][DATA][25] , 
        \chs_in_f[2][DATA][24] , \chs_in_f[2][DATA][23] , 
        \chs_in_f[2][DATA][22] , \chs_in_f[2][DATA][21] , 
        \chs_in_f[2][DATA][20] , \chs_in_f[2][DATA][19] , 
        \chs_in_f[2][DATA][18] , \chs_in_f[2][DATA][17] , 
        \chs_in_f[2][DATA][16] , \chs_in_f[2][DATA][15] , 
        \chs_in_f[2][DATA][14] , \chs_in_f[2][DATA][13] , 
        \chs_in_f[2][DATA][12] , \chs_in_f[2][DATA][11] , 
        \chs_in_f[2][DATA][10] , \chs_in_f[2][DATA][9] , 
        \chs_in_f[2][DATA][8] , \chs_in_f[2][DATA][7] , \chs_in_f[2][DATA][6] , 
        \chs_in_f[2][DATA][5] , \chs_in_f[2][DATA][4] , \chs_in_f[2][DATA][3] , 
        \chs_in_f[2][DATA][2] , \chs_in_f[2][DATA][1] , \chs_in_f[2][DATA][0] , 
        \chs_in_f[1][REQ] , \chs_in_f[1][DATA][34] , \chs_in_f[1][DATA][33] , 
        \chs_in_f[1][DATA][32] , \chs_in_f[1][DATA][31] , 
        \chs_in_f[1][DATA][30] , \chs_in_f[1][DATA][29] , 
        \chs_in_f[1][DATA][28] , \chs_in_f[1][DATA][27] , 
        \chs_in_f[1][DATA][26] , \chs_in_f[1][DATA][25] , 
        \chs_in_f[1][DATA][24] , \chs_in_f[1][DATA][23] , 
        \chs_in_f[1][DATA][22] , \chs_in_f[1][DATA][21] , 
        \chs_in_f[1][DATA][20] , \chs_in_f[1][DATA][19] , 
        \chs_in_f[1][DATA][18] , \chs_in_f[1][DATA][17] , 
        \chs_in_f[1][DATA][16] , \chs_in_f[1][DATA][15] , 
        \chs_in_f[1][DATA][14] , \chs_in_f[1][DATA][13] , 
        \chs_in_f[1][DATA][12] , \chs_in_f[1][DATA][11] , 
        \chs_in_f[1][DATA][10] , \chs_in_f[1][DATA][9] , 
        \chs_in_f[1][DATA][8] , \chs_in_f[1][DATA][7] , \chs_in_f[1][DATA][6] , 
        \chs_in_f[1][DATA][5] , \chs_in_f[1][DATA][4] , \chs_in_f[1][DATA][3] , 
        \chs_in_f[1][DATA][2] , \chs_in_f[1][DATA][1] , \chs_in_f[1][DATA][0] , 
        \chs_in_f[0][REQ] , \chs_in_f[0][DATA][34] , \chs_in_f[0][DATA][33] , 
        \chs_in_f[0][DATA][32] , \chs_in_f[0][DATA][31] , 
        \chs_in_f[0][DATA][30] , \chs_in_f[0][DATA][29] , 
        \chs_in_f[0][DATA][28] , \chs_in_f[0][DATA][27] , 
        \chs_in_f[0][DATA][26] , \chs_in_f[0][DATA][25] , 
        \chs_in_f[0][DATA][24] , \chs_in_f[0][DATA][23] , 
        \chs_in_f[0][DATA][22] , \chs_in_f[0][DATA][21] , 
        \chs_in_f[0][DATA][20] , \chs_in_f[0][DATA][19] , 
        \chs_in_f[0][DATA][18] , \chs_in_f[0][DATA][17] , 
        \chs_in_f[0][DATA][16] , \chs_in_f[0][DATA][15] , 
        \chs_in_f[0][DATA][14] , \chs_in_f[0][DATA][13] , 
        \chs_in_f[0][DATA][12] , \chs_in_f[0][DATA][11] , 
        \chs_in_f[0][DATA][10] , \chs_in_f[0][DATA][9] , 
        \chs_in_f[0][DATA][8] , \chs_in_f[0][DATA][7] , \chs_in_f[0][DATA][6] , 
        \chs_in_f[0][DATA][5] , \chs_in_f[0][DATA][4] , \chs_in_f[0][DATA][3] , 
        \chs_in_f[0][DATA][2] , \chs_in_f[0][DATA][1] , \chs_in_f[0][DATA][0] }), .chs_in_b({\chs_in_b[4][ACK] , \chs_in_b[3][ACK] , \chs_in_b[2][ACK] , 
        \chs_in_b[1][ACK] , \chs_in_b[0][ACK] }), .latches_out_f({
        \resource_out_f[REQ] , \resource_out_f[DATA][34] , 
        \resource_out_f[DATA][33] , \resource_out_f[DATA][32] , 
        \resource_out_f[DATA][31] , \resource_out_f[DATA][30] , 
        \resource_out_f[DATA][29] , \resource_out_f[DATA][28] , 
        \resource_out_f[DATA][27] , \resource_out_f[DATA][26] , 
        \resource_out_f[DATA][25] , \resource_out_f[DATA][24] , 
        \resource_out_f[DATA][23] , \resource_out_f[DATA][22] , 
        \resource_out_f[DATA][21] , \resource_out_f[DATA][20] , 
        \resource_out_f[DATA][19] , \resource_out_f[DATA][18] , 
        \resource_out_f[DATA][17] , \resource_out_f[DATA][16] , 
        \resource_out_f[DATA][15] , \resource_out_f[DATA][14] , 
        \resource_out_f[DATA][13] , \resource_out_f[DATA][12] , 
        \resource_out_f[DATA][11] , \resource_out_f[DATA][10] , 
        \resource_out_f[DATA][9] , \resource_out_f[DATA][8] , 
        \resource_out_f[DATA][7] , \resource_out_f[DATA][6] , 
        \resource_out_f[DATA][5] , \resource_out_f[DATA][4] , 
        \resource_out_f[DATA][3] , \resource_out_f[DATA][2] , 
        \resource_out_f[DATA][1] , \resource_out_f[DATA][0] , 
        \west_out_f[REQ] , \west_out_f[DATA][34] , \west_out_f[DATA][33] , 
        \west_out_f[DATA][32] , \west_out_f[DATA][31] , \west_out_f[DATA][30] , 
        \west_out_f[DATA][29] , \west_out_f[DATA][28] , \west_out_f[DATA][27] , 
        \west_out_f[DATA][26] , \west_out_f[DATA][25] , \west_out_f[DATA][24] , 
        \west_out_f[DATA][23] , \west_out_f[DATA][22] , \west_out_f[DATA][21] , 
        \west_out_f[DATA][20] , \west_out_f[DATA][19] , \west_out_f[DATA][18] , 
        \west_out_f[DATA][17] , \west_out_f[DATA][16] , \west_out_f[DATA][15] , 
        \west_out_f[DATA][14] , \west_out_f[DATA][13] , \west_out_f[DATA][12] , 
        \west_out_f[DATA][11] , \west_out_f[DATA][10] , \west_out_f[DATA][9] , 
        \west_out_f[DATA][8] , \west_out_f[DATA][7] , \west_out_f[DATA][6] , 
        \west_out_f[DATA][5] , \west_out_f[DATA][4] , \west_out_f[DATA][3] , 
        \west_out_f[DATA][2] , \west_out_f[DATA][1] , \west_out_f[DATA][0] , 
        \south_out_f[REQ] , \south_out_f[DATA][34] , \south_out_f[DATA][33] , 
        \south_out_f[DATA][32] , \south_out_f[DATA][31] , 
        \south_out_f[DATA][30] , \south_out_f[DATA][29] , 
        \south_out_f[DATA][28] , \south_out_f[DATA][27] , 
        \south_out_f[DATA][26] , \south_out_f[DATA][25] , 
        \south_out_f[DATA][24] , \south_out_f[DATA][23] , 
        \south_out_f[DATA][22] , \south_out_f[DATA][21] , 
        \south_out_f[DATA][20] , \south_out_f[DATA][19] , 
        \south_out_f[DATA][18] , \south_out_f[DATA][17] , 
        \south_out_f[DATA][16] , \south_out_f[DATA][15] , 
        \south_out_f[DATA][14] , \south_out_f[DATA][13] , 
        \south_out_f[DATA][12] , \south_out_f[DATA][11] , 
        \south_out_f[DATA][10] , \south_out_f[DATA][9] , 
        \south_out_f[DATA][8] , \south_out_f[DATA][7] , \south_out_f[DATA][6] , 
        \south_out_f[DATA][5] , \south_out_f[DATA][4] , \south_out_f[DATA][3] , 
        \south_out_f[DATA][2] , \south_out_f[DATA][1] , \south_out_f[DATA][0] , 
        \east_out_f[REQ] , \east_out_f[DATA][34] , \east_out_f[DATA][33] , 
        \east_out_f[DATA][32] , \east_out_f[DATA][31] , \east_out_f[DATA][30] , 
        \east_out_f[DATA][29] , \east_out_f[DATA][28] , \east_out_f[DATA][27] , 
        \east_out_f[DATA][26] , \east_out_f[DATA][25] , \east_out_f[DATA][24] , 
        \east_out_f[DATA][23] , \east_out_f[DATA][22] , \east_out_f[DATA][21] , 
        \east_out_f[DATA][20] , \east_out_f[DATA][19] , \east_out_f[DATA][18] , 
        \east_out_f[DATA][17] , \east_out_f[DATA][16] , \east_out_f[DATA][15] , 
        \east_out_f[DATA][14] , \east_out_f[DATA][13] , \east_out_f[DATA][12] , 
        \east_out_f[DATA][11] , \east_out_f[DATA][10] , \east_out_f[DATA][9] , 
        \east_out_f[DATA][8] , \east_out_f[DATA][7] , \east_out_f[DATA][6] , 
        \east_out_f[DATA][5] , \east_out_f[DATA][4] , \east_out_f[DATA][3] , 
        \east_out_f[DATA][2] , \east_out_f[DATA][1] , \east_out_f[DATA][0] , 
        \north_out_f[REQ] , \north_out_f[DATA][34] , \north_out_f[DATA][33] , 
        \north_out_f[DATA][32] , \north_out_f[DATA][31] , 
        \north_out_f[DATA][30] , \north_out_f[DATA][29] , 
        \north_out_f[DATA][28] , \north_out_f[DATA][27] , 
        \north_out_f[DATA][26] , \north_out_f[DATA][25] , 
        \north_out_f[DATA][24] , \north_out_f[DATA][23] , 
        \north_out_f[DATA][22] , \north_out_f[DATA][21] , 
        \north_out_f[DATA][20] , \north_out_f[DATA][19] , 
        \north_out_f[DATA][18] , \north_out_f[DATA][17] , 
        \north_out_f[DATA][16] , \north_out_f[DATA][15] , 
        \north_out_f[DATA][14] , \north_out_f[DATA][13] , 
        \north_out_f[DATA][12] , \north_out_f[DATA][11] , 
        \north_out_f[DATA][10] , \north_out_f[DATA][9] , 
        \north_out_f[DATA][8] , \north_out_f[DATA][7] , \north_out_f[DATA][6] , 
        \north_out_f[DATA][5] , \north_out_f[DATA][4] , \north_out_f[DATA][3] , 
        \north_out_f[DATA][2] , \north_out_f[DATA][1] , \north_out_f[DATA][0] }), .latches_out_b({\resource_out_b[ACK] , \west_out_b[ACK] , 
        \south_out_b[ACK] , \east_out_b[ACK] , \north_out_b[ACK] }) );
  HS65_LS_BFX9 U1 ( .A(preset), .Z(n3) );
  HS65_LS_BFX9 U2 ( .A(preset), .Z(n2) );
endmodule


module noc_node_1 ( p_clk, n_clk, reset, .proc_in({\proc_in[MCMD][1] , 
        \proc_in[MCMD][0] , \proc_in[MADDR][31] , \proc_in[MADDR][30] , 
        \proc_in[MADDR][29] , \proc_in[MADDR][28] , \proc_in[MADDR][27] , 
        \proc_in[MADDR][26] , \proc_in[MADDR][25] , \proc_in[MADDR][24] , 
        \proc_in[MADDR][23] , \proc_in[MADDR][22] , \proc_in[MADDR][21] , 
        \proc_in[MADDR][20] , \proc_in[MADDR][19] , \proc_in[MADDR][18] , 
        \proc_in[MADDR][17] , \proc_in[MADDR][16] , \proc_in[MADDR][15] , 
        \proc_in[MADDR][14] , \proc_in[MADDR][13] , \proc_in[MADDR][12] , 
        \proc_in[MADDR][11] , \proc_in[MADDR][10] , \proc_in[MADDR][9] , 
        \proc_in[MADDR][8] , \proc_in[MADDR][7] , \proc_in[MADDR][6] , 
        \proc_in[MADDR][5] , \proc_in[MADDR][4] , \proc_in[MADDR][3] , 
        \proc_in[MADDR][2] , \proc_in[MADDR][1] , \proc_in[MADDR][0] , 
        \proc_in[MDATA][31] , \proc_in[MDATA][30] , \proc_in[MDATA][29] , 
        \proc_in[MDATA][28] , \proc_in[MDATA][27] , \proc_in[MDATA][26] , 
        \proc_in[MDATA][25] , \proc_in[MDATA][24] , \proc_in[MDATA][23] , 
        \proc_in[MDATA][22] , \proc_in[MDATA][21] , \proc_in[MDATA][20] , 
        \proc_in[MDATA][19] , \proc_in[MDATA][18] , \proc_in[MDATA][17] , 
        \proc_in[MDATA][16] , \proc_in[MDATA][15] , \proc_in[MDATA][14] , 
        \proc_in[MDATA][13] , \proc_in[MDATA][12] , \proc_in[MDATA][11] , 
        \proc_in[MDATA][10] , \proc_in[MDATA][9] , \proc_in[MDATA][8] , 
        \proc_in[MDATA][7] , \proc_in[MDATA][6] , \proc_in[MDATA][5] , 
        \proc_in[MDATA][4] , \proc_in[MDATA][3] , \proc_in[MDATA][2] , 
        \proc_in[MDATA][1] , \proc_in[MDATA][0] }), .proc_out({
        \proc_out[SCMDACCEPT] , \proc_out[SRESP] , \proc_out[SDATA][31] , 
        \proc_out[SDATA][30] , \proc_out[SDATA][29] , \proc_out[SDATA][28] , 
        \proc_out[SDATA][27] , \proc_out[SDATA][26] , \proc_out[SDATA][25] , 
        \proc_out[SDATA][24] , \proc_out[SDATA][23] , \proc_out[SDATA][22] , 
        \proc_out[SDATA][21] , \proc_out[SDATA][20] , \proc_out[SDATA][19] , 
        \proc_out[SDATA][18] , \proc_out[SDATA][17] , \proc_out[SDATA][16] , 
        \proc_out[SDATA][15] , \proc_out[SDATA][14] , \proc_out[SDATA][13] , 
        \proc_out[SDATA][12] , \proc_out[SDATA][11] , \proc_out[SDATA][10] , 
        \proc_out[SDATA][9] , \proc_out[SDATA][8] , \proc_out[SDATA][7] , 
        \proc_out[SDATA][6] , \proc_out[SDATA][5] , \proc_out[SDATA][4] , 
        \proc_out[SDATA][3] , \proc_out[SDATA][2] , \proc_out[SDATA][1] , 
        \proc_out[SDATA][0] }), .spm_in({\spm_in[SCMDACCEPT] , \spm_in[SRESP] , 
        \spm_in[SDATA][63] , \spm_in[SDATA][62] , \spm_in[SDATA][61] , 
        \spm_in[SDATA][60] , \spm_in[SDATA][59] , \spm_in[SDATA][58] , 
        \spm_in[SDATA][57] , \spm_in[SDATA][56] , \spm_in[SDATA][55] , 
        \spm_in[SDATA][54] , \spm_in[SDATA][53] , \spm_in[SDATA][52] , 
        \spm_in[SDATA][51] , \spm_in[SDATA][50] , \spm_in[SDATA][49] , 
        \spm_in[SDATA][48] , \spm_in[SDATA][47] , \spm_in[SDATA][46] , 
        \spm_in[SDATA][45] , \spm_in[SDATA][44] , \spm_in[SDATA][43] , 
        \spm_in[SDATA][42] , \spm_in[SDATA][41] , \spm_in[SDATA][40] , 
        \spm_in[SDATA][39] , \spm_in[SDATA][38] , \spm_in[SDATA][37] , 
        \spm_in[SDATA][36] , \spm_in[SDATA][35] , \spm_in[SDATA][34] , 
        \spm_in[SDATA][33] , \spm_in[SDATA][32] , \spm_in[SDATA][31] , 
        \spm_in[SDATA][30] , \spm_in[SDATA][29] , \spm_in[SDATA][28] , 
        \spm_in[SDATA][27] , \spm_in[SDATA][26] , \spm_in[SDATA][25] , 
        \spm_in[SDATA][24] , \spm_in[SDATA][23] , \spm_in[SDATA][22] , 
        \spm_in[SDATA][21] , \spm_in[SDATA][20] , \spm_in[SDATA][19] , 
        \spm_in[SDATA][18] , \spm_in[SDATA][17] , \spm_in[SDATA][16] , 
        \spm_in[SDATA][15] , \spm_in[SDATA][14] , \spm_in[SDATA][13] , 
        \spm_in[SDATA][12] , \spm_in[SDATA][11] , \spm_in[SDATA][10] , 
        \spm_in[SDATA][9] , \spm_in[SDATA][8] , \spm_in[SDATA][7] , 
        \spm_in[SDATA][6] , \spm_in[SDATA][5] , \spm_in[SDATA][4] , 
        \spm_in[SDATA][3] , \spm_in[SDATA][2] , \spm_in[SDATA][1] , 
        \spm_in[SDATA][0] }), .spm_out({\spm_out[MCMD][1] , \spm_out[MCMD][0] , 
        \spm_out[MADDR][31] , \spm_out[MADDR][30] , \spm_out[MADDR][29] , 
        \spm_out[MADDR][28] , \spm_out[MADDR][27] , \spm_out[MADDR][26] , 
        \spm_out[MADDR][25] , \spm_out[MADDR][24] , \spm_out[MADDR][23] , 
        \spm_out[MADDR][22] , \spm_out[MADDR][21] , \spm_out[MADDR][20] , 
        \spm_out[MADDR][19] , \spm_out[MADDR][18] , \spm_out[MADDR][17] , 
        \spm_out[MADDR][16] , \spm_out[MADDR][15] , \spm_out[MADDR][14] , 
        \spm_out[MADDR][13] , \spm_out[MADDR][12] , \spm_out[MADDR][11] , 
        \spm_out[MADDR][10] , \spm_out[MADDR][9] , \spm_out[MADDR][8] , 
        \spm_out[MADDR][7] , \spm_out[MADDR][6] , \spm_out[MADDR][5] , 
        \spm_out[MADDR][4] , \spm_out[MADDR][3] , \spm_out[MADDR][2] , 
        \spm_out[MADDR][1] , \spm_out[MADDR][0] , \spm_out[MDATA][63] , 
        \spm_out[MDATA][62] , \spm_out[MDATA][61] , \spm_out[MDATA][60] , 
        \spm_out[MDATA][59] , \spm_out[MDATA][58] , \spm_out[MDATA][57] , 
        \spm_out[MDATA][56] , \spm_out[MDATA][55] , \spm_out[MDATA][54] , 
        \spm_out[MDATA][53] , \spm_out[MDATA][52] , \spm_out[MDATA][51] , 
        \spm_out[MDATA][50] , \spm_out[MDATA][49] , \spm_out[MDATA][48] , 
        \spm_out[MDATA][47] , \spm_out[MDATA][46] , \spm_out[MDATA][45] , 
        \spm_out[MDATA][44] , \spm_out[MDATA][43] , \spm_out[MDATA][42] , 
        \spm_out[MDATA][41] , \spm_out[MDATA][40] , \spm_out[MDATA][39] , 
        \spm_out[MDATA][38] , \spm_out[MDATA][37] , \spm_out[MDATA][36] , 
        \spm_out[MDATA][35] , \spm_out[MDATA][34] , \spm_out[MDATA][33] , 
        \spm_out[MDATA][32] , \spm_out[MDATA][31] , \spm_out[MDATA][30] , 
        \spm_out[MDATA][29] , \spm_out[MDATA][28] , \spm_out[MDATA][27] , 
        \spm_out[MDATA][26] , \spm_out[MDATA][25] , \spm_out[MDATA][24] , 
        \spm_out[MDATA][23] , \spm_out[MDATA][22] , \spm_out[MDATA][21] , 
        \spm_out[MDATA][20] , \spm_out[MDATA][19] , \spm_out[MDATA][18] , 
        \spm_out[MDATA][17] , \spm_out[MDATA][16] , \spm_out[MDATA][15] , 
        \spm_out[MDATA][14] , \spm_out[MDATA][13] , \spm_out[MDATA][12] , 
        \spm_out[MDATA][11] , \spm_out[MDATA][10] , \spm_out[MDATA][9] , 
        \spm_out[MDATA][8] , \spm_out[MDATA][7] , \spm_out[MDATA][6] , 
        \spm_out[MDATA][5] , \spm_out[MDATA][4] , \spm_out[MDATA][3] , 
        \spm_out[MDATA][2] , \spm_out[MDATA][1] , \spm_out[MDATA][0] }), 
    .north_in_f({\north_in_f[REQ] , \north_in_f[DATA][34] , 
        \north_in_f[DATA][33] , \north_in_f[DATA][32] , \north_in_f[DATA][31] , 
        \north_in_f[DATA][30] , \north_in_f[DATA][29] , \north_in_f[DATA][28] , 
        \north_in_f[DATA][27] , \north_in_f[DATA][26] , \north_in_f[DATA][25] , 
        \north_in_f[DATA][24] , \north_in_f[DATA][23] , \north_in_f[DATA][22] , 
        \north_in_f[DATA][21] , \north_in_f[DATA][20] , \north_in_f[DATA][19] , 
        \north_in_f[DATA][18] , \north_in_f[DATA][17] , \north_in_f[DATA][16] , 
        \north_in_f[DATA][15] , \north_in_f[DATA][14] , \north_in_f[DATA][13] , 
        \north_in_f[DATA][12] , \north_in_f[DATA][11] , \north_in_f[DATA][10] , 
        \north_in_f[DATA][9] , \north_in_f[DATA][8] , \north_in_f[DATA][7] , 
        \north_in_f[DATA][6] , \north_in_f[DATA][5] , \north_in_f[DATA][4] , 
        \north_in_f[DATA][3] , \north_in_f[DATA][2] , \north_in_f[DATA][1] , 
        \north_in_f[DATA][0] }), .north_in_b(\north_in_b[ACK] ), .east_in_f({
        \east_in_f[REQ] , \east_in_f[DATA][34] , \east_in_f[DATA][33] , 
        \east_in_f[DATA][32] , \east_in_f[DATA][31] , \east_in_f[DATA][30] , 
        \east_in_f[DATA][29] , \east_in_f[DATA][28] , \east_in_f[DATA][27] , 
        \east_in_f[DATA][26] , \east_in_f[DATA][25] , \east_in_f[DATA][24] , 
        \east_in_f[DATA][23] , \east_in_f[DATA][22] , \east_in_f[DATA][21] , 
        \east_in_f[DATA][20] , \east_in_f[DATA][19] , \east_in_f[DATA][18] , 
        \east_in_f[DATA][17] , \east_in_f[DATA][16] , \east_in_f[DATA][15] , 
        \east_in_f[DATA][14] , \east_in_f[DATA][13] , \east_in_f[DATA][12] , 
        \east_in_f[DATA][11] , \east_in_f[DATA][10] , \east_in_f[DATA][9] , 
        \east_in_f[DATA][8] , \east_in_f[DATA][7] , \east_in_f[DATA][6] , 
        \east_in_f[DATA][5] , \east_in_f[DATA][4] , \east_in_f[DATA][3] , 
        \east_in_f[DATA][2] , \east_in_f[DATA][1] , \east_in_f[DATA][0] }), 
    .east_in_b(\east_in_b[ACK] ), .south_in_f({\south_in_f[REQ] , 
        \south_in_f[DATA][34] , \south_in_f[DATA][33] , \south_in_f[DATA][32] , 
        \south_in_f[DATA][31] , \south_in_f[DATA][30] , \south_in_f[DATA][29] , 
        \south_in_f[DATA][28] , \south_in_f[DATA][27] , \south_in_f[DATA][26] , 
        \south_in_f[DATA][25] , \south_in_f[DATA][24] , \south_in_f[DATA][23] , 
        \south_in_f[DATA][22] , \south_in_f[DATA][21] , \south_in_f[DATA][20] , 
        \south_in_f[DATA][19] , \south_in_f[DATA][18] , \south_in_f[DATA][17] , 
        \south_in_f[DATA][16] , \south_in_f[DATA][15] , \south_in_f[DATA][14] , 
        \south_in_f[DATA][13] , \south_in_f[DATA][12] , \south_in_f[DATA][11] , 
        \south_in_f[DATA][10] , \south_in_f[DATA][9] , \south_in_f[DATA][8] , 
        \south_in_f[DATA][7] , \south_in_f[DATA][6] , \south_in_f[DATA][5] , 
        \south_in_f[DATA][4] , \south_in_f[DATA][3] , \south_in_f[DATA][2] , 
        \south_in_f[DATA][1] , \south_in_f[DATA][0] }), .south_in_b(
        \south_in_b[ACK] ), .west_in_f({\west_in_f[REQ] , 
        \west_in_f[DATA][34] , \west_in_f[DATA][33] , \west_in_f[DATA][32] , 
        \west_in_f[DATA][31] , \west_in_f[DATA][30] , \west_in_f[DATA][29] , 
        \west_in_f[DATA][28] , \west_in_f[DATA][27] , \west_in_f[DATA][26] , 
        \west_in_f[DATA][25] , \west_in_f[DATA][24] , \west_in_f[DATA][23] , 
        \west_in_f[DATA][22] , \west_in_f[DATA][21] , \west_in_f[DATA][20] , 
        \west_in_f[DATA][19] , \west_in_f[DATA][18] , \west_in_f[DATA][17] , 
        \west_in_f[DATA][16] , \west_in_f[DATA][15] , \west_in_f[DATA][14] , 
        \west_in_f[DATA][13] , \west_in_f[DATA][12] , \west_in_f[DATA][11] , 
        \west_in_f[DATA][10] , \west_in_f[DATA][9] , \west_in_f[DATA][8] , 
        \west_in_f[DATA][7] , \west_in_f[DATA][6] , \west_in_f[DATA][5] , 
        \west_in_f[DATA][4] , \west_in_f[DATA][3] , \west_in_f[DATA][2] , 
        \west_in_f[DATA][1] , \west_in_f[DATA][0] }), .west_in_b(
        \west_in_b[ACK] ), .north_out_f({\north_out_f[REQ] , 
        \north_out_f[DATA][34] , \north_out_f[DATA][33] , 
        \north_out_f[DATA][32] , \north_out_f[DATA][31] , 
        \north_out_f[DATA][30] , \north_out_f[DATA][29] , 
        \north_out_f[DATA][28] , \north_out_f[DATA][27] , 
        \north_out_f[DATA][26] , \north_out_f[DATA][25] , 
        \north_out_f[DATA][24] , \north_out_f[DATA][23] , 
        \north_out_f[DATA][22] , \north_out_f[DATA][21] , 
        \north_out_f[DATA][20] , \north_out_f[DATA][19] , 
        \north_out_f[DATA][18] , \north_out_f[DATA][17] , 
        \north_out_f[DATA][16] , \north_out_f[DATA][15] , 
        \north_out_f[DATA][14] , \north_out_f[DATA][13] , 
        \north_out_f[DATA][12] , \north_out_f[DATA][11] , 
        \north_out_f[DATA][10] , \north_out_f[DATA][9] , 
        \north_out_f[DATA][8] , \north_out_f[DATA][7] , \north_out_f[DATA][6] , 
        \north_out_f[DATA][5] , \north_out_f[DATA][4] , \north_out_f[DATA][3] , 
        \north_out_f[DATA][2] , \north_out_f[DATA][1] , \north_out_f[DATA][0] 
        }), .north_out_b(\north_out_b[ACK] ), .east_out_f({\east_out_f[REQ] , 
        \east_out_f[DATA][34] , \east_out_f[DATA][33] , \east_out_f[DATA][32] , 
        \east_out_f[DATA][31] , \east_out_f[DATA][30] , \east_out_f[DATA][29] , 
        \east_out_f[DATA][28] , \east_out_f[DATA][27] , \east_out_f[DATA][26] , 
        \east_out_f[DATA][25] , \east_out_f[DATA][24] , \east_out_f[DATA][23] , 
        \east_out_f[DATA][22] , \east_out_f[DATA][21] , \east_out_f[DATA][20] , 
        \east_out_f[DATA][19] , \east_out_f[DATA][18] , \east_out_f[DATA][17] , 
        \east_out_f[DATA][16] , \east_out_f[DATA][15] , \east_out_f[DATA][14] , 
        \east_out_f[DATA][13] , \east_out_f[DATA][12] , \east_out_f[DATA][11] , 
        \east_out_f[DATA][10] , \east_out_f[DATA][9] , \east_out_f[DATA][8] , 
        \east_out_f[DATA][7] , \east_out_f[DATA][6] , \east_out_f[DATA][5] , 
        \east_out_f[DATA][4] , \east_out_f[DATA][3] , \east_out_f[DATA][2] , 
        \east_out_f[DATA][1] , \east_out_f[DATA][0] }), .east_out_b(
        \east_out_b[ACK] ), .south_out_f({\south_out_f[REQ] , 
        \south_out_f[DATA][34] , \south_out_f[DATA][33] , 
        \south_out_f[DATA][32] , \south_out_f[DATA][31] , 
        \south_out_f[DATA][30] , \south_out_f[DATA][29] , 
        \south_out_f[DATA][28] , \south_out_f[DATA][27] , 
        \south_out_f[DATA][26] , \south_out_f[DATA][25] , 
        \south_out_f[DATA][24] , \south_out_f[DATA][23] , 
        \south_out_f[DATA][22] , \south_out_f[DATA][21] , 
        \south_out_f[DATA][20] , \south_out_f[DATA][19] , 
        \south_out_f[DATA][18] , \south_out_f[DATA][17] , 
        \south_out_f[DATA][16] , \south_out_f[DATA][15] , 
        \south_out_f[DATA][14] , \south_out_f[DATA][13] , 
        \south_out_f[DATA][12] , \south_out_f[DATA][11] , 
        \south_out_f[DATA][10] , \south_out_f[DATA][9] , 
        \south_out_f[DATA][8] , \south_out_f[DATA][7] , \south_out_f[DATA][6] , 
        \south_out_f[DATA][5] , \south_out_f[DATA][4] , \south_out_f[DATA][3] , 
        \south_out_f[DATA][2] , \south_out_f[DATA][1] , \south_out_f[DATA][0] 
        }), .south_out_b(\south_out_b[ACK] ), .west_out_f({\west_out_f[REQ] , 
        \west_out_f[DATA][34] , \west_out_f[DATA][33] , \west_out_f[DATA][32] , 
        \west_out_f[DATA][31] , \west_out_f[DATA][30] , \west_out_f[DATA][29] , 
        \west_out_f[DATA][28] , \west_out_f[DATA][27] , \west_out_f[DATA][26] , 
        \west_out_f[DATA][25] , \west_out_f[DATA][24] , \west_out_f[DATA][23] , 
        \west_out_f[DATA][22] , \west_out_f[DATA][21] , \west_out_f[DATA][20] , 
        \west_out_f[DATA][19] , \west_out_f[DATA][18] , \west_out_f[DATA][17] , 
        \west_out_f[DATA][16] , \west_out_f[DATA][15] , \west_out_f[DATA][14] , 
        \west_out_f[DATA][13] , \west_out_f[DATA][12] , \west_out_f[DATA][11] , 
        \west_out_f[DATA][10] , \west_out_f[DATA][9] , \west_out_f[DATA][8] , 
        \west_out_f[DATA][7] , \west_out_f[DATA][6] , \west_out_f[DATA][5] , 
        \west_out_f[DATA][4] , \west_out_f[DATA][3] , \west_out_f[DATA][2] , 
        \west_out_f[DATA][1] , \west_out_f[DATA][0] }), .west_out_b(
        \west_out_b[ACK] ) );
  input p_clk, n_clk, reset, \proc_in[MCMD][1] , \proc_in[MCMD][0] ,
         \proc_in[MADDR][31] , \proc_in[MADDR][30] , \proc_in[MADDR][29] ,
         \proc_in[MADDR][28] , \proc_in[MADDR][27] , \proc_in[MADDR][26] ,
         \proc_in[MADDR][25] , \proc_in[MADDR][24] , \proc_in[MADDR][23] ,
         \proc_in[MADDR][22] , \proc_in[MADDR][21] , \proc_in[MADDR][20] ,
         \proc_in[MADDR][19] , \proc_in[MADDR][18] , \proc_in[MADDR][17] ,
         \proc_in[MADDR][16] , \proc_in[MADDR][15] , \proc_in[MADDR][14] ,
         \proc_in[MADDR][13] , \proc_in[MADDR][12] , \proc_in[MADDR][11] ,
         \proc_in[MADDR][10] , \proc_in[MADDR][9] , \proc_in[MADDR][8] ,
         \proc_in[MADDR][7] , \proc_in[MADDR][6] , \proc_in[MADDR][5] ,
         \proc_in[MADDR][4] , \proc_in[MADDR][3] , \proc_in[MADDR][2] ,
         \proc_in[MADDR][1] , \proc_in[MADDR][0] , \proc_in[MDATA][31] ,
         \proc_in[MDATA][30] , \proc_in[MDATA][29] , \proc_in[MDATA][28] ,
         \proc_in[MDATA][27] , \proc_in[MDATA][26] , \proc_in[MDATA][25] ,
         \proc_in[MDATA][24] , \proc_in[MDATA][23] , \proc_in[MDATA][22] ,
         \proc_in[MDATA][21] , \proc_in[MDATA][20] , \proc_in[MDATA][19] ,
         \proc_in[MDATA][18] , \proc_in[MDATA][17] , \proc_in[MDATA][16] ,
         \proc_in[MDATA][15] , \proc_in[MDATA][14] , \proc_in[MDATA][13] ,
         \proc_in[MDATA][12] , \proc_in[MDATA][11] , \proc_in[MDATA][10] ,
         \proc_in[MDATA][9] , \proc_in[MDATA][8] , \proc_in[MDATA][7] ,
         \proc_in[MDATA][6] , \proc_in[MDATA][5] , \proc_in[MDATA][4] ,
         \proc_in[MDATA][3] , \proc_in[MDATA][2] , \proc_in[MDATA][1] ,
         \proc_in[MDATA][0] , \spm_in[SCMDACCEPT] , \spm_in[SRESP] ,
         \spm_in[SDATA][63] , \spm_in[SDATA][62] , \spm_in[SDATA][61] ,
         \spm_in[SDATA][60] , \spm_in[SDATA][59] , \spm_in[SDATA][58] ,
         \spm_in[SDATA][57] , \spm_in[SDATA][56] , \spm_in[SDATA][55] ,
         \spm_in[SDATA][54] , \spm_in[SDATA][53] , \spm_in[SDATA][52] ,
         \spm_in[SDATA][51] , \spm_in[SDATA][50] , \spm_in[SDATA][49] ,
         \spm_in[SDATA][48] , \spm_in[SDATA][47] , \spm_in[SDATA][46] ,
         \spm_in[SDATA][45] , \spm_in[SDATA][44] , \spm_in[SDATA][43] ,
         \spm_in[SDATA][42] , \spm_in[SDATA][41] , \spm_in[SDATA][40] ,
         \spm_in[SDATA][39] , \spm_in[SDATA][38] , \spm_in[SDATA][37] ,
         \spm_in[SDATA][36] , \spm_in[SDATA][35] , \spm_in[SDATA][34] ,
         \spm_in[SDATA][33] , \spm_in[SDATA][32] , \spm_in[SDATA][31] ,
         \spm_in[SDATA][30] , \spm_in[SDATA][29] , \spm_in[SDATA][28] ,
         \spm_in[SDATA][27] , \spm_in[SDATA][26] , \spm_in[SDATA][25] ,
         \spm_in[SDATA][24] , \spm_in[SDATA][23] , \spm_in[SDATA][22] ,
         \spm_in[SDATA][21] , \spm_in[SDATA][20] , \spm_in[SDATA][19] ,
         \spm_in[SDATA][18] , \spm_in[SDATA][17] , \spm_in[SDATA][16] ,
         \spm_in[SDATA][15] , \spm_in[SDATA][14] , \spm_in[SDATA][13] ,
         \spm_in[SDATA][12] , \spm_in[SDATA][11] , \spm_in[SDATA][10] ,
         \spm_in[SDATA][9] , \spm_in[SDATA][8] , \spm_in[SDATA][7] ,
         \spm_in[SDATA][6] , \spm_in[SDATA][5] , \spm_in[SDATA][4] ,
         \spm_in[SDATA][3] , \spm_in[SDATA][2] , \spm_in[SDATA][1] ,
         \spm_in[SDATA][0] , \north_in_f[REQ] , \north_in_f[DATA][34] ,
         \north_in_f[DATA][33] , \north_in_f[DATA][32] ,
         \north_in_f[DATA][31] , \north_in_f[DATA][30] ,
         \north_in_f[DATA][29] , \north_in_f[DATA][28] ,
         \north_in_f[DATA][27] , \north_in_f[DATA][26] ,
         \north_in_f[DATA][25] , \north_in_f[DATA][24] ,
         \north_in_f[DATA][23] , \north_in_f[DATA][22] ,
         \north_in_f[DATA][21] , \north_in_f[DATA][20] ,
         \north_in_f[DATA][19] , \north_in_f[DATA][18] ,
         \north_in_f[DATA][17] , \north_in_f[DATA][16] ,
         \north_in_f[DATA][15] , \north_in_f[DATA][14] ,
         \north_in_f[DATA][13] , \north_in_f[DATA][12] ,
         \north_in_f[DATA][11] , \north_in_f[DATA][10] , \north_in_f[DATA][9] ,
         \north_in_f[DATA][8] , \north_in_f[DATA][7] , \north_in_f[DATA][6] ,
         \north_in_f[DATA][5] , \north_in_f[DATA][4] , \north_in_f[DATA][3] ,
         \north_in_f[DATA][2] , \north_in_f[DATA][1] , \north_in_f[DATA][0] ,
         \east_in_f[REQ] , \east_in_f[DATA][34] , \east_in_f[DATA][33] ,
         \east_in_f[DATA][32] , \east_in_f[DATA][31] , \east_in_f[DATA][30] ,
         \east_in_f[DATA][29] , \east_in_f[DATA][28] , \east_in_f[DATA][27] ,
         \east_in_f[DATA][26] , \east_in_f[DATA][25] , \east_in_f[DATA][24] ,
         \east_in_f[DATA][23] , \east_in_f[DATA][22] , \east_in_f[DATA][21] ,
         \east_in_f[DATA][20] , \east_in_f[DATA][19] , \east_in_f[DATA][18] ,
         \east_in_f[DATA][17] , \east_in_f[DATA][16] , \east_in_f[DATA][15] ,
         \east_in_f[DATA][14] , \east_in_f[DATA][13] , \east_in_f[DATA][12] ,
         \east_in_f[DATA][11] , \east_in_f[DATA][10] , \east_in_f[DATA][9] ,
         \east_in_f[DATA][8] , \east_in_f[DATA][7] , \east_in_f[DATA][6] ,
         \east_in_f[DATA][5] , \east_in_f[DATA][4] , \east_in_f[DATA][3] ,
         \east_in_f[DATA][2] , \east_in_f[DATA][1] , \east_in_f[DATA][0] ,
         \south_in_f[REQ] , \south_in_f[DATA][34] , \south_in_f[DATA][33] ,
         \south_in_f[DATA][32] , \south_in_f[DATA][31] ,
         \south_in_f[DATA][30] , \south_in_f[DATA][29] ,
         \south_in_f[DATA][28] , \south_in_f[DATA][27] ,
         \south_in_f[DATA][26] , \south_in_f[DATA][25] ,
         \south_in_f[DATA][24] , \south_in_f[DATA][23] ,
         \south_in_f[DATA][22] , \south_in_f[DATA][21] ,
         \south_in_f[DATA][20] , \south_in_f[DATA][19] ,
         \south_in_f[DATA][18] , \south_in_f[DATA][17] ,
         \south_in_f[DATA][16] , \south_in_f[DATA][15] ,
         \south_in_f[DATA][14] , \south_in_f[DATA][13] ,
         \south_in_f[DATA][12] , \south_in_f[DATA][11] ,
         \south_in_f[DATA][10] , \south_in_f[DATA][9] , \south_in_f[DATA][8] ,
         \south_in_f[DATA][7] , \south_in_f[DATA][6] , \south_in_f[DATA][5] ,
         \south_in_f[DATA][4] , \south_in_f[DATA][3] , \south_in_f[DATA][2] ,
         \south_in_f[DATA][1] , \south_in_f[DATA][0] , \west_in_f[REQ] ,
         \west_in_f[DATA][34] , \west_in_f[DATA][33] , \west_in_f[DATA][32] ,
         \west_in_f[DATA][31] , \west_in_f[DATA][30] , \west_in_f[DATA][29] ,
         \west_in_f[DATA][28] , \west_in_f[DATA][27] , \west_in_f[DATA][26] ,
         \west_in_f[DATA][25] , \west_in_f[DATA][24] , \west_in_f[DATA][23] ,
         \west_in_f[DATA][22] , \west_in_f[DATA][21] , \west_in_f[DATA][20] ,
         \west_in_f[DATA][19] , \west_in_f[DATA][18] , \west_in_f[DATA][17] ,
         \west_in_f[DATA][16] , \west_in_f[DATA][15] , \west_in_f[DATA][14] ,
         \west_in_f[DATA][13] , \west_in_f[DATA][12] , \west_in_f[DATA][11] ,
         \west_in_f[DATA][10] , \west_in_f[DATA][9] , \west_in_f[DATA][8] ,
         \west_in_f[DATA][7] , \west_in_f[DATA][6] , \west_in_f[DATA][5] ,
         \west_in_f[DATA][4] , \west_in_f[DATA][3] , \west_in_f[DATA][2] ,
         \west_in_f[DATA][1] , \west_in_f[DATA][0] , \north_out_b[ACK] ,
         \east_out_b[ACK] , \south_out_b[ACK] , \west_out_b[ACK] ;
  output \proc_out[SCMDACCEPT] , \proc_out[SRESP] , \proc_out[SDATA][31] ,
         \proc_out[SDATA][30] , \proc_out[SDATA][29] , \proc_out[SDATA][28] ,
         \proc_out[SDATA][27] , \proc_out[SDATA][26] , \proc_out[SDATA][25] ,
         \proc_out[SDATA][24] , \proc_out[SDATA][23] , \proc_out[SDATA][22] ,
         \proc_out[SDATA][21] , \proc_out[SDATA][20] , \proc_out[SDATA][19] ,
         \proc_out[SDATA][18] , \proc_out[SDATA][17] , \proc_out[SDATA][16] ,
         \proc_out[SDATA][15] , \proc_out[SDATA][14] , \proc_out[SDATA][13] ,
         \proc_out[SDATA][12] , \proc_out[SDATA][11] , \proc_out[SDATA][10] ,
         \proc_out[SDATA][9] , \proc_out[SDATA][8] , \proc_out[SDATA][7] ,
         \proc_out[SDATA][6] , \proc_out[SDATA][5] , \proc_out[SDATA][4] ,
         \proc_out[SDATA][3] , \proc_out[SDATA][2] , \proc_out[SDATA][1] ,
         \proc_out[SDATA][0] , \spm_out[MCMD][1] , \spm_out[MCMD][0] ,
         \spm_out[MADDR][31] , \spm_out[MADDR][30] , \spm_out[MADDR][29] ,
         \spm_out[MADDR][28] , \spm_out[MADDR][27] , \spm_out[MADDR][26] ,
         \spm_out[MADDR][25] , \spm_out[MADDR][24] , \spm_out[MADDR][23] ,
         \spm_out[MADDR][22] , \spm_out[MADDR][21] , \spm_out[MADDR][20] ,
         \spm_out[MADDR][19] , \spm_out[MADDR][18] , \spm_out[MADDR][17] ,
         \spm_out[MADDR][16] , \spm_out[MADDR][15] , \spm_out[MADDR][14] ,
         \spm_out[MADDR][13] , \spm_out[MADDR][12] , \spm_out[MADDR][11] ,
         \spm_out[MADDR][10] , \spm_out[MADDR][9] , \spm_out[MADDR][8] ,
         \spm_out[MADDR][7] , \spm_out[MADDR][6] , \spm_out[MADDR][5] ,
         \spm_out[MADDR][4] , \spm_out[MADDR][3] , \spm_out[MADDR][2] ,
         \spm_out[MADDR][1] , \spm_out[MADDR][0] , \spm_out[MDATA][63] ,
         \spm_out[MDATA][62] , \spm_out[MDATA][61] , \spm_out[MDATA][60] ,
         \spm_out[MDATA][59] , \spm_out[MDATA][58] , \spm_out[MDATA][57] ,
         \spm_out[MDATA][56] , \spm_out[MDATA][55] , \spm_out[MDATA][54] ,
         \spm_out[MDATA][53] , \spm_out[MDATA][52] , \spm_out[MDATA][51] ,
         \spm_out[MDATA][50] , \spm_out[MDATA][49] , \spm_out[MDATA][48] ,
         \spm_out[MDATA][47] , \spm_out[MDATA][46] , \spm_out[MDATA][45] ,
         \spm_out[MDATA][44] , \spm_out[MDATA][43] , \spm_out[MDATA][42] ,
         \spm_out[MDATA][41] , \spm_out[MDATA][40] , \spm_out[MDATA][39] ,
         \spm_out[MDATA][38] , \spm_out[MDATA][37] , \spm_out[MDATA][36] ,
         \spm_out[MDATA][35] , \spm_out[MDATA][34] , \spm_out[MDATA][33] ,
         \spm_out[MDATA][32] , \spm_out[MDATA][31] , \spm_out[MDATA][30] ,
         \spm_out[MDATA][29] , \spm_out[MDATA][28] , \spm_out[MDATA][27] ,
         \spm_out[MDATA][26] , \spm_out[MDATA][25] , \spm_out[MDATA][24] ,
         \spm_out[MDATA][23] , \spm_out[MDATA][22] , \spm_out[MDATA][21] ,
         \spm_out[MDATA][20] , \spm_out[MDATA][19] , \spm_out[MDATA][18] ,
         \spm_out[MDATA][17] , \spm_out[MDATA][16] , \spm_out[MDATA][15] ,
         \spm_out[MDATA][14] , \spm_out[MDATA][13] , \spm_out[MDATA][12] ,
         \spm_out[MDATA][11] , \spm_out[MDATA][10] , \spm_out[MDATA][9] ,
         \spm_out[MDATA][8] , \spm_out[MDATA][7] , \spm_out[MDATA][6] ,
         \spm_out[MDATA][5] , \spm_out[MDATA][4] , \spm_out[MDATA][3] ,
         \spm_out[MDATA][2] , \spm_out[MDATA][1] , \spm_out[MDATA][0] ,
         \north_in_b[ACK] , \east_in_b[ACK] , \south_in_b[ACK] ,
         \west_in_b[ACK] , \north_out_f[REQ] , \north_out_f[DATA][34] ,
         \north_out_f[DATA][33] , \north_out_f[DATA][32] ,
         \north_out_f[DATA][31] , \north_out_f[DATA][30] ,
         \north_out_f[DATA][29] , \north_out_f[DATA][28] ,
         \north_out_f[DATA][27] , \north_out_f[DATA][26] ,
         \north_out_f[DATA][25] , \north_out_f[DATA][24] ,
         \north_out_f[DATA][23] , \north_out_f[DATA][22] ,
         \north_out_f[DATA][21] , \north_out_f[DATA][20] ,
         \north_out_f[DATA][19] , \north_out_f[DATA][18] ,
         \north_out_f[DATA][17] , \north_out_f[DATA][16] ,
         \north_out_f[DATA][15] , \north_out_f[DATA][14] ,
         \north_out_f[DATA][13] , \north_out_f[DATA][12] ,
         \north_out_f[DATA][11] , \north_out_f[DATA][10] ,
         \north_out_f[DATA][9] , \north_out_f[DATA][8] ,
         \north_out_f[DATA][7] , \north_out_f[DATA][6] ,
         \north_out_f[DATA][5] , \north_out_f[DATA][4] ,
         \north_out_f[DATA][3] , \north_out_f[DATA][2] ,
         \north_out_f[DATA][1] , \north_out_f[DATA][0] , \east_out_f[REQ] ,
         \east_out_f[DATA][34] , \east_out_f[DATA][33] ,
         \east_out_f[DATA][32] , \east_out_f[DATA][31] ,
         \east_out_f[DATA][30] , \east_out_f[DATA][29] ,
         \east_out_f[DATA][28] , \east_out_f[DATA][27] ,
         \east_out_f[DATA][26] , \east_out_f[DATA][25] ,
         \east_out_f[DATA][24] , \east_out_f[DATA][23] ,
         \east_out_f[DATA][22] , \east_out_f[DATA][21] ,
         \east_out_f[DATA][20] , \east_out_f[DATA][19] ,
         \east_out_f[DATA][18] , \east_out_f[DATA][17] ,
         \east_out_f[DATA][16] , \east_out_f[DATA][15] ,
         \east_out_f[DATA][14] , \east_out_f[DATA][13] ,
         \east_out_f[DATA][12] , \east_out_f[DATA][11] ,
         \east_out_f[DATA][10] , \east_out_f[DATA][9] , \east_out_f[DATA][8] ,
         \east_out_f[DATA][7] , \east_out_f[DATA][6] , \east_out_f[DATA][5] ,
         \east_out_f[DATA][4] , \east_out_f[DATA][3] , \east_out_f[DATA][2] ,
         \east_out_f[DATA][1] , \east_out_f[DATA][0] , \south_out_f[REQ] ,
         \south_out_f[DATA][34] , \south_out_f[DATA][33] ,
         \south_out_f[DATA][32] , \south_out_f[DATA][31] ,
         \south_out_f[DATA][30] , \south_out_f[DATA][29] ,
         \south_out_f[DATA][28] , \south_out_f[DATA][27] ,
         \south_out_f[DATA][26] , \south_out_f[DATA][25] ,
         \south_out_f[DATA][24] , \south_out_f[DATA][23] ,
         \south_out_f[DATA][22] , \south_out_f[DATA][21] ,
         \south_out_f[DATA][20] , \south_out_f[DATA][19] ,
         \south_out_f[DATA][18] , \south_out_f[DATA][17] ,
         \south_out_f[DATA][16] , \south_out_f[DATA][15] ,
         \south_out_f[DATA][14] , \south_out_f[DATA][13] ,
         \south_out_f[DATA][12] , \south_out_f[DATA][11] ,
         \south_out_f[DATA][10] , \south_out_f[DATA][9] ,
         \south_out_f[DATA][8] , \south_out_f[DATA][7] ,
         \south_out_f[DATA][6] , \south_out_f[DATA][5] ,
         \south_out_f[DATA][4] , \south_out_f[DATA][3] ,
         \south_out_f[DATA][2] , \south_out_f[DATA][1] ,
         \south_out_f[DATA][0] , \west_out_f[REQ] , \west_out_f[DATA][34] ,
         \west_out_f[DATA][33] , \west_out_f[DATA][32] ,
         \west_out_f[DATA][31] , \west_out_f[DATA][30] ,
         \west_out_f[DATA][29] , \west_out_f[DATA][28] ,
         \west_out_f[DATA][27] , \west_out_f[DATA][26] ,
         \west_out_f[DATA][25] , \west_out_f[DATA][24] ,
         \west_out_f[DATA][23] , \west_out_f[DATA][22] ,
         \west_out_f[DATA][21] , \west_out_f[DATA][20] ,
         \west_out_f[DATA][19] , \west_out_f[DATA][18] ,
         \west_out_f[DATA][17] , \west_out_f[DATA][16] ,
         \west_out_f[DATA][15] , \west_out_f[DATA][14] ,
         \west_out_f[DATA][13] , \west_out_f[DATA][12] ,
         \west_out_f[DATA][11] , \west_out_f[DATA][10] , \west_out_f[DATA][9] ,
         \west_out_f[DATA][8] , \west_out_f[DATA][7] , \west_out_f[DATA][6] ,
         \west_out_f[DATA][5] , \west_out_f[DATA][4] , \west_out_f[DATA][3] ,
         \west_out_f[DATA][2] , \west_out_f[DATA][1] , \west_out_f[DATA][0] ;
  wire   del_half_clk0, \ip_to_net_f[REQ] , n1, n3, n4, n5, n6, n7, n8, n9,
         n10, n11;
  wire   [34:0] net_to_ip;
  wire   [34:0] ip_to_net;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17;
  assign \spm_out[MADDR][31]  = 1'b0;
  assign \spm_out[MADDR][30]  = 1'b0;
  assign \spm_out[MADDR][29]  = 1'b0;
  assign \spm_out[MADDR][28]  = 1'b0;
  assign \spm_out[MADDR][27]  = 1'b0;
  assign \spm_out[MADDR][26]  = 1'b0;
  assign \spm_out[MADDR][25]  = 1'b0;
  assign \spm_out[MADDR][24]  = 1'b0;
  assign \spm_out[MADDR][23]  = 1'b0;
  assign \spm_out[MADDR][22]  = 1'b0;
  assign \spm_out[MADDR][21]  = 1'b0;
  assign \spm_out[MADDR][20]  = 1'b0;
  assign \spm_out[MADDR][19]  = 1'b0;
  assign \spm_out[MADDR][18]  = 1'b0;
  assign \spm_out[MADDR][17]  = 1'b0;
  assign \spm_out[MADDR][16]  = 1'b0;
  assign \spm_out[MADDR][15]  = 1'b0;

  nAdapter_1 na ( .na_clk(n_clk), .na_reset(reset), .proc_in({
        \proc_in[MCMD][1] , \proc_in[MCMD][0] , \proc_in[MADDR][31] , 
        \proc_in[MADDR][30] , \proc_in[MADDR][29] , \proc_in[MADDR][28] , 
        \proc_in[MADDR][27] , \proc_in[MADDR][26] , \proc_in[MADDR][25] , 
        \proc_in[MADDR][24] , \proc_in[MADDR][23] , \proc_in[MADDR][22] , 
        \proc_in[MADDR][21] , \proc_in[MADDR][20] , \proc_in[MADDR][19] , 
        \proc_in[MADDR][18] , \proc_in[MADDR][17] , \proc_in[MADDR][16] , 
        \proc_in[MADDR][15] , \proc_in[MADDR][14] , \proc_in[MADDR][13] , 
        \proc_in[MADDR][12] , \proc_in[MADDR][11] , \proc_in[MADDR][10] , 
        \proc_in[MADDR][9] , \proc_in[MADDR][8] , \proc_in[MADDR][7] , 
        \proc_in[MADDR][6] , \proc_in[MADDR][5] , \proc_in[MADDR][4] , 
        \proc_in[MADDR][3] , \proc_in[MADDR][2] , \proc_in[MADDR][1] , 
        \proc_in[MADDR][0] , \proc_in[MDATA][31] , \proc_in[MDATA][30] , 
        \proc_in[MDATA][29] , \proc_in[MDATA][28] , \proc_in[MDATA][27] , 
        \proc_in[MDATA][26] , \proc_in[MDATA][25] , \proc_in[MDATA][24] , 
        \proc_in[MDATA][23] , \proc_in[MDATA][22] , \proc_in[MDATA][21] , 
        \proc_in[MDATA][20] , \proc_in[MDATA][19] , \proc_in[MDATA][18] , 
        \proc_in[MDATA][17] , \proc_in[MDATA][16] , \proc_in[MDATA][15] , 
        \proc_in[MDATA][14] , \proc_in[MDATA][13] , \proc_in[MDATA][12] , 
        \proc_in[MDATA][11] , \proc_in[MDATA][10] , \proc_in[MDATA][9] , 
        \proc_in[MDATA][8] , \proc_in[MDATA][7] , \proc_in[MDATA][6] , 
        \proc_in[MDATA][5] , \proc_in[MDATA][4] , \proc_in[MDATA][3] , 
        \proc_in[MDATA][2] , \proc_in[MDATA][1] , \proc_in[MDATA][0] }), 
        .proc_out({\proc_out[SCMDACCEPT] , \proc_out[SRESP] , 
        \proc_out[SDATA][31] , \proc_out[SDATA][30] , \proc_out[SDATA][29] , 
        \proc_out[SDATA][28] , \proc_out[SDATA][27] , \proc_out[SDATA][26] , 
        \proc_out[SDATA][25] , \proc_out[SDATA][24] , \proc_out[SDATA][23] , 
        \proc_out[SDATA][22] , \proc_out[SDATA][21] , \proc_out[SDATA][20] , 
        \proc_out[SDATA][19] , \proc_out[SDATA][18] , \proc_out[SDATA][17] , 
        \proc_out[SDATA][16] , \proc_out[SDATA][15] , \proc_out[SDATA][14] , 
        \proc_out[SDATA][13] , \proc_out[SDATA][12] , \proc_out[SDATA][11] , 
        \proc_out[SDATA][10] , \proc_out[SDATA][9] , \proc_out[SDATA][8] , 
        \proc_out[SDATA][7] , \proc_out[SDATA][6] , \proc_out[SDATA][5] , 
        \proc_out[SDATA][4] , \proc_out[SDATA][3] , \proc_out[SDATA][2] , 
        \proc_out[SDATA][1] , \proc_out[SDATA][0] }), .spm_in({
        \spm_in[SCMDACCEPT] , \spm_in[SRESP] , \spm_in[SDATA][63] , 
        \spm_in[SDATA][62] , \spm_in[SDATA][61] , \spm_in[SDATA][60] , 
        \spm_in[SDATA][59] , \spm_in[SDATA][58] , \spm_in[SDATA][57] , 
        \spm_in[SDATA][56] , \spm_in[SDATA][55] , \spm_in[SDATA][54] , 
        \spm_in[SDATA][53] , \spm_in[SDATA][52] , \spm_in[SDATA][51] , 
        \spm_in[SDATA][50] , \spm_in[SDATA][49] , \spm_in[SDATA][48] , 
        \spm_in[SDATA][47] , \spm_in[SDATA][46] , \spm_in[SDATA][45] , 
        \spm_in[SDATA][44] , \spm_in[SDATA][43] , \spm_in[SDATA][42] , 
        \spm_in[SDATA][41] , \spm_in[SDATA][40] , \spm_in[SDATA][39] , 
        \spm_in[SDATA][38] , \spm_in[SDATA][37] , \spm_in[SDATA][36] , 
        \spm_in[SDATA][35] , \spm_in[SDATA][34] , \spm_in[SDATA][33] , 
        \spm_in[SDATA][32] , \spm_in[SDATA][31] , \spm_in[SDATA][30] , 
        \spm_in[SDATA][29] , \spm_in[SDATA][28] , \spm_in[SDATA][27] , 
        \spm_in[SDATA][26] , \spm_in[SDATA][25] , \spm_in[SDATA][24] , 
        \spm_in[SDATA][23] , \spm_in[SDATA][22] , \spm_in[SDATA][21] , 
        \spm_in[SDATA][20] , \spm_in[SDATA][19] , \spm_in[SDATA][18] , 
        \spm_in[SDATA][17] , \spm_in[SDATA][16] , \spm_in[SDATA][15] , 
        \spm_in[SDATA][14] , \spm_in[SDATA][13] , \spm_in[SDATA][12] , 
        \spm_in[SDATA][11] , \spm_in[SDATA][10] , \spm_in[SDATA][9] , 
        \spm_in[SDATA][8] , \spm_in[SDATA][7] , \spm_in[SDATA][6] , 
        \spm_in[SDATA][5] , \spm_in[SDATA][4] , \spm_in[SDATA][3] , 
        \spm_in[SDATA][2] , \spm_in[SDATA][1] , \spm_in[SDATA][0] }), 
        .spm_out({\spm_out[MCMD][1] , \spm_out[MCMD][0] , 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, \spm_out[MADDR][14] , \spm_out[MADDR][13] , 
        \spm_out[MADDR][12] , \spm_out[MADDR][11] , \spm_out[MADDR][10] , 
        \spm_out[MADDR][9] , \spm_out[MADDR][8] , \spm_out[MADDR][7] , 
        \spm_out[MADDR][6] , \spm_out[MADDR][5] , \spm_out[MADDR][4] , 
        \spm_out[MADDR][3] , \spm_out[MADDR][2] , \spm_out[MADDR][1] , 
        \spm_out[MADDR][0] , \spm_out[MDATA][63] , \spm_out[MDATA][62] , 
        \spm_out[MDATA][61] , \spm_out[MDATA][60] , \spm_out[MDATA][59] , 
        \spm_out[MDATA][58] , \spm_out[MDATA][57] , \spm_out[MDATA][56] , 
        \spm_out[MDATA][55] , \spm_out[MDATA][54] , \spm_out[MDATA][53] , 
        \spm_out[MDATA][52] , \spm_out[MDATA][51] , \spm_out[MDATA][50] , 
        \spm_out[MDATA][49] , \spm_out[MDATA][48] , \spm_out[MDATA][47] , 
        \spm_out[MDATA][46] , \spm_out[MDATA][45] , \spm_out[MDATA][44] , 
        \spm_out[MDATA][43] , \spm_out[MDATA][42] , \spm_out[MDATA][41] , 
        \spm_out[MDATA][40] , \spm_out[MDATA][39] , \spm_out[MDATA][38] , 
        \spm_out[MDATA][37] , \spm_out[MDATA][36] , \spm_out[MDATA][35] , 
        \spm_out[MDATA][34] , \spm_out[MDATA][33] , \spm_out[MDATA][32] , 
        \spm_out[MDATA][31] , \spm_out[MDATA][30] , \spm_out[MDATA][29] , 
        \spm_out[MDATA][28] , \spm_out[MDATA][27] , \spm_out[MDATA][26] , 
        \spm_out[MDATA][25] , \spm_out[MDATA][24] , \spm_out[MDATA][23] , 
        \spm_out[MDATA][22] , \spm_out[MDATA][21] , \spm_out[MDATA][20] , 
        \spm_out[MDATA][19] , \spm_out[MDATA][18] , \spm_out[MDATA][17] , 
        \spm_out[MDATA][16] , \spm_out[MDATA][15] , \spm_out[MDATA][14] , 
        \spm_out[MDATA][13] , \spm_out[MDATA][12] , \spm_out[MDATA][11] , 
        \spm_out[MDATA][10] , \spm_out[MDATA][9] , \spm_out[MDATA][8] , 
        \spm_out[MDATA][7] , \spm_out[MDATA][6] , \spm_out[MDATA][5] , 
        \spm_out[MDATA][4] , \spm_out[MDATA][3] , \spm_out[MDATA][2] , 
        \spm_out[MDATA][1] , \spm_out[MDATA][0] }), .pkt_in(net_to_ip), 
        .pkt_out(ip_to_net) );
  noc_switch_1 r ( .preset(reset), .north_in_f({\north_in_f[REQ] , 
        \north_in_f[DATA][34] , \north_in_f[DATA][33] , \north_in_f[DATA][32] , 
        \north_in_f[DATA][31] , \north_in_f[DATA][30] , \north_in_f[DATA][29] , 
        \north_in_f[DATA][28] , \north_in_f[DATA][27] , \north_in_f[DATA][26] , 
        \north_in_f[DATA][25] , \north_in_f[DATA][24] , \north_in_f[DATA][23] , 
        \north_in_f[DATA][22] , \north_in_f[DATA][21] , \north_in_f[DATA][20] , 
        \north_in_f[DATA][19] , \north_in_f[DATA][18] , \north_in_f[DATA][17] , 
        \north_in_f[DATA][16] , \north_in_f[DATA][15] , \north_in_f[DATA][14] , 
        \north_in_f[DATA][13] , \north_in_f[DATA][12] , \north_in_f[DATA][11] , 
        \north_in_f[DATA][10] , \north_in_f[DATA][9] , \north_in_f[DATA][8] , 
        \north_in_f[DATA][7] , \north_in_f[DATA][6] , \north_in_f[DATA][5] , 
        \north_in_f[DATA][4] , \north_in_f[DATA][3] , \north_in_f[DATA][2] , 
        \north_in_f[DATA][1] , \north_in_f[DATA][0] }), .north_in_b(
        \north_in_b[ACK] ), .east_in_f({\east_in_f[REQ] , 
        \east_in_f[DATA][34] , \east_in_f[DATA][33] , \east_in_f[DATA][32] , 
        \east_in_f[DATA][31] , \east_in_f[DATA][30] , \east_in_f[DATA][29] , 
        \east_in_f[DATA][28] , \east_in_f[DATA][27] , \east_in_f[DATA][26] , 
        \east_in_f[DATA][25] , \east_in_f[DATA][24] , \east_in_f[DATA][23] , 
        \east_in_f[DATA][22] , \east_in_f[DATA][21] , \east_in_f[DATA][20] , 
        \east_in_f[DATA][19] , \east_in_f[DATA][18] , \east_in_f[DATA][17] , 
        \east_in_f[DATA][16] , \east_in_f[DATA][15] , \east_in_f[DATA][14] , 
        \east_in_f[DATA][13] , \east_in_f[DATA][12] , \east_in_f[DATA][11] , 
        \east_in_f[DATA][10] , \east_in_f[DATA][9] , \east_in_f[DATA][8] , 
        \east_in_f[DATA][7] , \east_in_f[DATA][6] , \east_in_f[DATA][5] , 
        \east_in_f[DATA][4] , \east_in_f[DATA][3] , \east_in_f[DATA][2] , 
        \east_in_f[DATA][1] , \east_in_f[DATA][0] }), .east_in_b(
        \east_in_b[ACK] ), .south_in_f({\south_in_f[REQ] , 
        \south_in_f[DATA][34] , \south_in_f[DATA][33] , \south_in_f[DATA][32] , 
        \south_in_f[DATA][31] , \south_in_f[DATA][30] , \south_in_f[DATA][29] , 
        \south_in_f[DATA][28] , \south_in_f[DATA][27] , \south_in_f[DATA][26] , 
        \south_in_f[DATA][25] , \south_in_f[DATA][24] , \south_in_f[DATA][23] , 
        \south_in_f[DATA][22] , \south_in_f[DATA][21] , \south_in_f[DATA][20] , 
        \south_in_f[DATA][19] , \south_in_f[DATA][18] , \south_in_f[DATA][17] , 
        \south_in_f[DATA][16] , \south_in_f[DATA][15] , \south_in_f[DATA][14] , 
        \south_in_f[DATA][13] , \south_in_f[DATA][12] , \south_in_f[DATA][11] , 
        \south_in_f[DATA][10] , \south_in_f[DATA][9] , \south_in_f[DATA][8] , 
        \south_in_f[DATA][7] , \south_in_f[DATA][6] , \south_in_f[DATA][5] , 
        \south_in_f[DATA][4] , \south_in_f[DATA][3] , \south_in_f[DATA][2] , 
        \south_in_f[DATA][1] , \south_in_f[DATA][0] }), .south_in_b(
        \south_in_b[ACK] ), .west_in_f({\west_in_f[REQ] , 
        \west_in_f[DATA][34] , \west_in_f[DATA][33] , \west_in_f[DATA][32] , 
        \west_in_f[DATA][31] , \west_in_f[DATA][30] , \west_in_f[DATA][29] , 
        \west_in_f[DATA][28] , \west_in_f[DATA][27] , \west_in_f[DATA][26] , 
        \west_in_f[DATA][25] , \west_in_f[DATA][24] , \west_in_f[DATA][23] , 
        \west_in_f[DATA][22] , \west_in_f[DATA][21] , \west_in_f[DATA][20] , 
        \west_in_f[DATA][19] , \west_in_f[DATA][18] , \west_in_f[DATA][17] , 
        \west_in_f[DATA][16] , \west_in_f[DATA][15] , \west_in_f[DATA][14] , 
        \west_in_f[DATA][13] , \west_in_f[DATA][12] , \west_in_f[DATA][11] , 
        \west_in_f[DATA][10] , \west_in_f[DATA][9] , \west_in_f[DATA][8] , 
        \west_in_f[DATA][7] , \west_in_f[DATA][6] , \west_in_f[DATA][5] , 
        \west_in_f[DATA][4] , \west_in_f[DATA][3] , \west_in_f[DATA][2] , 
        \west_in_f[DATA][1] , \west_in_f[DATA][0] }), .west_in_b(
        \west_in_b[ACK] ), .resource_in_f({\ip_to_net_f[REQ] , ip_to_net}), 
        .north_out_f({\north_out_f[REQ] , \north_out_f[DATA][34] , 
        \north_out_f[DATA][33] , \north_out_f[DATA][32] , 
        \north_out_f[DATA][31] , \north_out_f[DATA][30] , 
        \north_out_f[DATA][29] , \north_out_f[DATA][28] , 
        \north_out_f[DATA][27] , \north_out_f[DATA][26] , 
        \north_out_f[DATA][25] , \north_out_f[DATA][24] , 
        \north_out_f[DATA][23] , \north_out_f[DATA][22] , 
        \north_out_f[DATA][21] , \north_out_f[DATA][20] , 
        \north_out_f[DATA][19] , \north_out_f[DATA][18] , 
        \north_out_f[DATA][17] , \north_out_f[DATA][16] , 
        \north_out_f[DATA][15] , \north_out_f[DATA][14] , 
        \north_out_f[DATA][13] , \north_out_f[DATA][12] , 
        \north_out_f[DATA][11] , \north_out_f[DATA][10] , 
        \north_out_f[DATA][9] , \north_out_f[DATA][8] , \north_out_f[DATA][7] , 
        \north_out_f[DATA][6] , \north_out_f[DATA][5] , \north_out_f[DATA][4] , 
        \north_out_f[DATA][3] , \north_out_f[DATA][2] , \north_out_f[DATA][1] , 
        \north_out_f[DATA][0] }), .north_out_b(\north_out_b[ACK] ), 
        .east_out_f({\east_out_f[REQ] , \east_out_f[DATA][34] , 
        \east_out_f[DATA][33] , \east_out_f[DATA][32] , \east_out_f[DATA][31] , 
        \east_out_f[DATA][30] , \east_out_f[DATA][29] , \east_out_f[DATA][28] , 
        \east_out_f[DATA][27] , \east_out_f[DATA][26] , \east_out_f[DATA][25] , 
        \east_out_f[DATA][24] , \east_out_f[DATA][23] , \east_out_f[DATA][22] , 
        \east_out_f[DATA][21] , \east_out_f[DATA][20] , \east_out_f[DATA][19] , 
        \east_out_f[DATA][18] , \east_out_f[DATA][17] , \east_out_f[DATA][16] , 
        \east_out_f[DATA][15] , \east_out_f[DATA][14] , \east_out_f[DATA][13] , 
        \east_out_f[DATA][12] , \east_out_f[DATA][11] , \east_out_f[DATA][10] , 
        \east_out_f[DATA][9] , \east_out_f[DATA][8] , \east_out_f[DATA][7] , 
        \east_out_f[DATA][6] , \east_out_f[DATA][5] , \east_out_f[DATA][4] , 
        \east_out_f[DATA][3] , \east_out_f[DATA][2] , \east_out_f[DATA][1] , 
        \east_out_f[DATA][0] }), .east_out_b(\east_out_b[ACK] ), .south_out_f(
        {\south_out_f[REQ] , \south_out_f[DATA][34] , \south_out_f[DATA][33] , 
        \south_out_f[DATA][32] , \south_out_f[DATA][31] , 
        \south_out_f[DATA][30] , \south_out_f[DATA][29] , 
        \south_out_f[DATA][28] , \south_out_f[DATA][27] , 
        \south_out_f[DATA][26] , \south_out_f[DATA][25] , 
        \south_out_f[DATA][24] , \south_out_f[DATA][23] , 
        \south_out_f[DATA][22] , \south_out_f[DATA][21] , 
        \south_out_f[DATA][20] , \south_out_f[DATA][19] , 
        \south_out_f[DATA][18] , \south_out_f[DATA][17] , 
        \south_out_f[DATA][16] , \south_out_f[DATA][15] , 
        \south_out_f[DATA][14] , \south_out_f[DATA][13] , 
        \south_out_f[DATA][12] , \south_out_f[DATA][11] , 
        \south_out_f[DATA][10] , \south_out_f[DATA][9] , 
        \south_out_f[DATA][8] , \south_out_f[DATA][7] , \south_out_f[DATA][6] , 
        \south_out_f[DATA][5] , \south_out_f[DATA][4] , \south_out_f[DATA][3] , 
        \south_out_f[DATA][2] , \south_out_f[DATA][1] , \south_out_f[DATA][0] }), .south_out_b(\south_out_b[ACK] ), .west_out_f({\west_out_f[REQ] , 
        \west_out_f[DATA][34] , \west_out_f[DATA][33] , \west_out_f[DATA][32] , 
        \west_out_f[DATA][31] , \west_out_f[DATA][30] , \west_out_f[DATA][29] , 
        \west_out_f[DATA][28] , \west_out_f[DATA][27] , \west_out_f[DATA][26] , 
        \west_out_f[DATA][25] , \west_out_f[DATA][24] , \west_out_f[DATA][23] , 
        \west_out_f[DATA][22] , \west_out_f[DATA][21] , \west_out_f[DATA][20] , 
        \west_out_f[DATA][19] , \west_out_f[DATA][18] , \west_out_f[DATA][17] , 
        \west_out_f[DATA][16] , \west_out_f[DATA][15] , \west_out_f[DATA][14] , 
        \west_out_f[DATA][13] , \west_out_f[DATA][12] , \west_out_f[DATA][11] , 
        \west_out_f[DATA][10] , \west_out_f[DATA][9] , \west_out_f[DATA][8] , 
        \west_out_f[DATA][7] , \west_out_f[DATA][6] , \west_out_f[DATA][5] , 
        \west_out_f[DATA][4] , \west_out_f[DATA][3] , \west_out_f[DATA][2] , 
        \west_out_f[DATA][1] , \west_out_f[DATA][0] }), .west_out_b(
        \west_out_b[ACK] ), .resource_out_f({SYNOPSYS_UNCONNECTED__17, 
        net_to_ip}), .resource_out_b(n9) );
  HS65_LS_DFPRQNX9 half_clk_reg ( .D(n11), .CP(n_clk), .RN(n8), .QN(n11) );
  HS65_LS_IVX9 I_2 ( .A(n4), .Z(\ip_to_net_f[REQ] ) );
  HS65_LH_IVX2 I_1 ( .A(n10), .Z(del_half_clk0) );
  HS65_LS_IVX9 U3 ( .A(n11), .Z(n10) );
  HS65_LH_IVX2 U4 ( .A(n1), .Z(n3) );
  HS65_LS_IVX106 U5 ( .A(del_half_clk0), .Z(n1) );
  HS65_LS_BFX9 U6 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U7 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U8 ( .A(n7), .Z(n6) );
  HS65_LS_BFX9 U9 ( .A(n3), .Z(n7) );
  HS65_LS_IVX9 U10 ( .A(reset), .Z(n8) );
  HS65_LS_IVX9 U11 ( .A(del_half_clk0), .Z(n9) );
endmodule


module noc ( p_clk, n_clk, reset, p_ports_in, p_ports_out, spm_ports_in, 
        spm_ports_out );
  input [263:0] p_ports_in;
  output [135:0] p_ports_out;
  input [263:0] spm_ports_in;
  output [391:0] spm_ports_out;
  input p_clk, n_clk, reset;
  wire   spm_ports_out_1__1__MADDR__31_, spm_ports_out_1__1__MADDR__30_,
         spm_ports_out_1__1__MADDR__29_, spm_ports_out_1__1__MADDR__28_,
         spm_ports_out_1__1__MADDR__27_, spm_ports_out_1__1__MADDR__26_,
         spm_ports_out_1__1__MADDR__25_, spm_ports_out_1__1__MADDR__24_,
         spm_ports_out_1__1__MADDR__23_, spm_ports_out_1__1__MADDR__22_,
         spm_ports_out_1__1__MADDR__21_, spm_ports_out_1__1__MADDR__20_,
         spm_ports_out_1__1__MADDR__19_, spm_ports_out_1__1__MADDR__18_,
         spm_ports_out_1__1__MADDR__17_, spm_ports_out_1__1__MADDR__16_, n258,
         spm_ports_out_1__0__MADDR__31_, spm_ports_out_1__0__MADDR__30_,
         spm_ports_out_1__0__MADDR__29_, spm_ports_out_1__0__MADDR__28_,
         spm_ports_out_1__0__MADDR__27_, spm_ports_out_1__0__MADDR__26_,
         spm_ports_out_1__0__MADDR__25_, spm_ports_out_1__0__MADDR__24_,
         spm_ports_out_1__0__MADDR__23_, spm_ports_out_1__0__MADDR__22_,
         spm_ports_out_1__0__MADDR__21_, spm_ports_out_1__0__MADDR__20_,
         spm_ports_out_1__0__MADDR__19_, spm_ports_out_1__0__MADDR__18_,
         spm_ports_out_1__0__MADDR__17_, spm_ports_out_1__0__MADDR__16_,
         spm_ports_out_1__0__MADDR__15_, spm_ports_out_0__1__MADDR__31_,
         spm_ports_out_0__1__MADDR__30_, spm_ports_out_0__1__MADDR__29_,
         spm_ports_out_0__1__MADDR__28_, spm_ports_out_0__1__MADDR__27_,
         spm_ports_out_0__1__MADDR__26_, spm_ports_out_0__1__MADDR__25_,
         spm_ports_out_0__1__MADDR__24_, spm_ports_out_0__1__MADDR__23_,
         spm_ports_out_0__1__MADDR__22_, spm_ports_out_0__1__MADDR__21_,
         spm_ports_out_0__1__MADDR__20_, spm_ports_out_0__1__MADDR__19_,
         spm_ports_out_0__1__MADDR__18_, spm_ports_out_0__1__MADDR__17_,
         spm_ports_out_0__1__MADDR__16_, spm_ports_out_0__1__MADDR__15_,
         spm_ports_out_0__0__MADDR__31_, spm_ports_out_0__0__MADDR__30_,
         spm_ports_out_0__0__MADDR__29_, spm_ports_out_0__0__MADDR__28_,
         spm_ports_out_0__0__MADDR__27_, spm_ports_out_0__0__MADDR__26_,
         spm_ports_out_0__0__MADDR__25_, spm_ports_out_0__0__MADDR__24_,
         spm_ports_out_0__0__MADDR__23_, spm_ports_out_0__0__MADDR__22_,
         spm_ports_out_0__0__MADDR__21_, spm_ports_out_0__0__MADDR__20_,
         spm_ports_out_0__0__MADDR__19_, spm_ports_out_0__0__MADDR__18_,
         spm_ports_out_0__0__MADDR__17_, spm_ports_out_0__0__MADDR__16_,
         spm_ports_out_0__0__MADDR__15_, west_out_0__0__FORWARD__REQ_,
         west_out_0__1__FORWARD__REQ_, west_out_0__1__FORWARD__DATA__34_,
         west_out_0__1__FORWARD__DATA__33_, west_out_0__1__FORWARD__DATA__32_,
         west_out_0__1__FORWARD__DATA__31_, west_out_0__1__FORWARD__DATA__30_,
         west_out_0__1__FORWARD__DATA__29_, west_out_0__1__FORWARD__DATA__28_,
         west_out_0__1__FORWARD__DATA__27_, west_out_0__1__FORWARD__DATA__26_,
         west_out_0__1__FORWARD__DATA__25_, west_out_0__1__FORWARD__DATA__24_,
         west_out_0__1__FORWARD__DATA__23_, west_out_0__1__FORWARD__DATA__22_,
         west_out_0__1__FORWARD__DATA__21_, west_out_0__1__FORWARD__DATA__20_,
         west_out_0__1__FORWARD__DATA__19_, west_out_0__1__FORWARD__DATA__18_,
         west_out_0__1__FORWARD__DATA__17_, west_out_0__1__FORWARD__DATA__16_,
         west_out_0__1__FORWARD__DATA__15_, west_out_0__1__FORWARD__DATA__14_,
         west_out_0__1__FORWARD__DATA__13_, west_out_0__1__FORWARD__DATA__12_,
         west_out_0__1__FORWARD__DATA__11_, west_out_0__1__FORWARD__DATA__10_,
         west_out_0__1__FORWARD__DATA__9_, west_out_0__1__FORWARD__DATA__8_,
         west_out_0__1__FORWARD__DATA__7_, west_out_0__1__FORWARD__DATA__6_,
         west_out_0__1__FORWARD__DATA__5_, west_out_0__1__FORWARD__DATA__4_,
         west_out_0__1__FORWARD__DATA__3_, west_out_0__1__FORWARD__DATA__2_,
         west_out_0__1__FORWARD__DATA__1_, west_out_0__1__FORWARD__DATA__0_,
         west_out_1__0__FORWARD__REQ_, west_out_1__0__FORWARD__DATA__34_,
         west_out_1__0__FORWARD__DATA__33_, west_out_1__0__FORWARD__DATA__32_,
         west_out_1__0__FORWARD__DATA__31_, west_out_1__0__FORWARD__DATA__30_,
         west_out_1__0__FORWARD__DATA__29_, west_out_1__0__FORWARD__DATA__28_,
         west_out_1__0__FORWARD__DATA__27_, west_out_1__0__FORWARD__DATA__26_,
         west_out_1__0__FORWARD__DATA__25_, west_out_1__0__FORWARD__DATA__24_,
         west_out_1__0__FORWARD__DATA__23_, west_out_1__0__FORWARD__DATA__22_,
         west_out_1__0__FORWARD__DATA__21_, west_out_1__0__FORWARD__DATA__20_,
         west_out_1__0__FORWARD__DATA__19_, west_out_1__0__FORWARD__DATA__18_,
         west_out_1__0__FORWARD__DATA__17_, west_out_1__0__FORWARD__DATA__16_,
         west_out_1__0__FORWARD__DATA__15_, west_out_1__0__FORWARD__DATA__14_,
         west_out_1__0__FORWARD__DATA__13_, west_out_1__0__FORWARD__DATA__12_,
         west_out_1__0__FORWARD__DATA__11_, west_out_1__0__FORWARD__DATA__10_,
         west_out_1__0__FORWARD__DATA__9_, west_out_1__0__FORWARD__DATA__8_,
         west_out_1__0__FORWARD__DATA__7_, west_out_1__0__FORWARD__DATA__6_,
         west_out_1__0__FORWARD__DATA__5_, west_out_1__0__FORWARD__DATA__4_,
         west_out_1__0__FORWARD__DATA__3_, west_out_1__0__FORWARD__DATA__2_,
         west_out_1__0__FORWARD__DATA__1_, west_out_1__0__FORWARD__DATA__0_,
         west_out_1__1__FORWARD__REQ_, west_out_1__1__FORWARD__DATA__34_,
         west_out_1__1__FORWARD__DATA__33_, west_out_1__1__FORWARD__DATA__32_,
         west_out_1__1__FORWARD__DATA__31_, west_out_1__1__FORWARD__DATA__30_,
         west_out_1__1__FORWARD__DATA__29_, west_out_1__1__FORWARD__DATA__28_,
         west_out_1__1__FORWARD__DATA__27_, west_out_1__1__FORWARD__DATA__26_,
         west_out_1__1__FORWARD__DATA__25_, west_out_1__1__FORWARD__DATA__24_,
         west_out_1__1__FORWARD__DATA__23_, west_out_1__1__FORWARD__DATA__22_,
         west_out_1__1__FORWARD__DATA__21_, west_out_1__1__FORWARD__DATA__20_,
         west_out_1__1__FORWARD__DATA__19_, west_out_1__1__FORWARD__DATA__18_,
         west_out_1__1__FORWARD__DATA__17_, west_out_1__1__FORWARD__DATA__16_,
         west_out_1__1__FORWARD__DATA__15_, west_out_1__1__FORWARD__DATA__14_,
         west_out_1__1__FORWARD__DATA__13_, west_out_1__1__FORWARD__DATA__12_,
         west_out_1__1__FORWARD__DATA__11_, west_out_1__1__FORWARD__DATA__10_,
         west_out_1__1__FORWARD__DATA__9_, west_out_1__1__FORWARD__DATA__8_,
         west_out_1__1__FORWARD__DATA__7_, west_out_1__1__FORWARD__DATA__6_,
         west_out_1__1__FORWARD__DATA__5_, west_out_1__1__FORWARD__DATA__4_,
         west_out_1__1__FORWARD__DATA__3_, west_out_1__1__FORWARD__DATA__2_,
         west_out_1__1__FORWARD__DATA__1_, west_out_1__1__FORWARD__DATA__0_,
         south_out_0__0__FORWARD__REQ_, south_out_0__0__FORWARD__DATA__34_,
         south_out_0__0__FORWARD__DATA__33_,
         south_out_0__0__FORWARD__DATA__32_,
         south_out_0__0__FORWARD__DATA__31_,
         south_out_0__0__FORWARD__DATA__30_,
         south_out_0__0__FORWARD__DATA__29_,
         south_out_0__0__FORWARD__DATA__28_,
         south_out_0__0__FORWARD__DATA__27_,
         south_out_0__0__FORWARD__DATA__26_,
         south_out_0__0__FORWARD__DATA__25_,
         south_out_0__0__FORWARD__DATA__24_,
         south_out_0__0__FORWARD__DATA__23_,
         south_out_0__0__FORWARD__DATA__22_,
         south_out_0__0__FORWARD__DATA__21_,
         south_out_0__0__FORWARD__DATA__20_,
         south_out_0__0__FORWARD__DATA__19_,
         south_out_0__0__FORWARD__DATA__18_,
         south_out_0__0__FORWARD__DATA__17_,
         south_out_0__0__FORWARD__DATA__16_,
         south_out_0__0__FORWARD__DATA__15_,
         south_out_0__0__FORWARD__DATA__14_,
         south_out_0__0__FORWARD__DATA__13_,
         south_out_0__0__FORWARD__DATA__12_,
         south_out_0__0__FORWARD__DATA__11_,
         south_out_0__0__FORWARD__DATA__10_, south_out_0__0__FORWARD__DATA__9_,
         south_out_0__0__FORWARD__DATA__8_, south_out_0__0__FORWARD__DATA__7_,
         south_out_0__0__FORWARD__DATA__6_, south_out_0__0__FORWARD__DATA__5_,
         south_out_0__0__FORWARD__DATA__4_, south_out_0__0__FORWARD__DATA__3_,
         south_out_0__0__FORWARD__DATA__2_, south_out_0__0__FORWARD__DATA__1_,
         south_out_0__0__FORWARD__DATA__0_, south_out_0__1__FORWARD__REQ_,
         south_out_0__1__FORWARD__DATA__34_,
         south_out_0__1__FORWARD__DATA__33_,
         south_out_0__1__FORWARD__DATA__32_,
         south_out_0__1__FORWARD__DATA__31_,
         south_out_0__1__FORWARD__DATA__30_,
         south_out_0__1__FORWARD__DATA__29_,
         south_out_0__1__FORWARD__DATA__28_,
         south_out_0__1__FORWARD__DATA__27_,
         south_out_0__1__FORWARD__DATA__26_,
         south_out_0__1__FORWARD__DATA__25_,
         south_out_0__1__FORWARD__DATA__24_,
         south_out_0__1__FORWARD__DATA__23_,
         south_out_0__1__FORWARD__DATA__22_,
         south_out_0__1__FORWARD__DATA__21_,
         south_out_0__1__FORWARD__DATA__20_,
         south_out_0__1__FORWARD__DATA__19_,
         south_out_0__1__FORWARD__DATA__18_,
         south_out_0__1__FORWARD__DATA__17_,
         south_out_0__1__FORWARD__DATA__16_,
         south_out_0__1__FORWARD__DATA__15_,
         south_out_0__1__FORWARD__DATA__14_,
         south_out_0__1__FORWARD__DATA__13_,
         south_out_0__1__FORWARD__DATA__12_,
         south_out_0__1__FORWARD__DATA__11_,
         south_out_0__1__FORWARD__DATA__10_, south_out_0__1__FORWARD__DATA__9_,
         south_out_0__1__FORWARD__DATA__8_, south_out_0__1__FORWARD__DATA__7_,
         south_out_0__1__FORWARD__DATA__6_, south_out_0__1__FORWARD__DATA__5_,
         south_out_0__1__FORWARD__DATA__4_, south_out_0__1__FORWARD__DATA__3_,
         south_out_0__1__FORWARD__DATA__2_, south_out_0__1__FORWARD__DATA__1_,
         south_out_0__1__FORWARD__DATA__0_, south_out_1__0__FORWARD__REQ_,
         south_out_1__1__FORWARD__REQ_, south_out_1__1__FORWARD__DATA__34_,
         south_out_1__1__FORWARD__DATA__33_,
         south_out_1__1__FORWARD__DATA__32_,
         south_out_1__1__FORWARD__DATA__31_,
         south_out_1__1__FORWARD__DATA__30_,
         south_out_1__1__FORWARD__DATA__29_,
         south_out_1__1__FORWARD__DATA__28_,
         south_out_1__1__FORWARD__DATA__27_,
         south_out_1__1__FORWARD__DATA__26_,
         south_out_1__1__FORWARD__DATA__25_,
         south_out_1__1__FORWARD__DATA__24_,
         south_out_1__1__FORWARD__DATA__23_,
         south_out_1__1__FORWARD__DATA__22_,
         south_out_1__1__FORWARD__DATA__21_,
         south_out_1__1__FORWARD__DATA__20_,
         south_out_1__1__FORWARD__DATA__19_,
         south_out_1__1__FORWARD__DATA__18_,
         south_out_1__1__FORWARD__DATA__17_,
         south_out_1__1__FORWARD__DATA__16_,
         south_out_1__1__FORWARD__DATA__15_,
         south_out_1__1__FORWARD__DATA__14_,
         south_out_1__1__FORWARD__DATA__13_,
         south_out_1__1__FORWARD__DATA__12_,
         south_out_1__1__FORWARD__DATA__11_,
         south_out_1__1__FORWARD__DATA__10_, south_out_1__1__FORWARD__DATA__9_,
         south_out_1__1__FORWARD__DATA__8_, south_out_1__1__FORWARD__DATA__7_,
         south_out_1__1__FORWARD__DATA__6_, south_out_1__1__FORWARD__DATA__5_,
         south_out_1__1__FORWARD__DATA__4_, south_out_1__1__FORWARD__DATA__3_,
         south_out_1__1__FORWARD__DATA__2_, south_out_1__1__FORWARD__DATA__1_,
         south_out_1__1__FORWARD__DATA__0_, east_out_0__0__FORWARD__REQ_,
         east_out_0__0__FORWARD__DATA__34_, east_out_0__0__FORWARD__DATA__33_,
         east_out_0__0__FORWARD__DATA__32_, east_out_0__0__FORWARD__DATA__31_,
         east_out_0__0__FORWARD__DATA__30_, east_out_0__0__FORWARD__DATA__29_,
         east_out_0__0__FORWARD__DATA__28_, east_out_0__0__FORWARD__DATA__27_,
         east_out_0__0__FORWARD__DATA__26_, east_out_0__0__FORWARD__DATA__25_,
         east_out_0__0__FORWARD__DATA__24_, east_out_0__0__FORWARD__DATA__23_,
         east_out_0__0__FORWARD__DATA__22_, east_out_0__0__FORWARD__DATA__21_,
         east_out_0__0__FORWARD__DATA__20_, east_out_0__0__FORWARD__DATA__19_,
         east_out_0__0__FORWARD__DATA__18_, east_out_0__0__FORWARD__DATA__17_,
         east_out_0__0__FORWARD__DATA__16_, east_out_0__0__FORWARD__DATA__15_,
         east_out_0__0__FORWARD__DATA__14_, east_out_0__0__FORWARD__DATA__13_,
         east_out_0__0__FORWARD__DATA__12_, east_out_0__0__FORWARD__DATA__11_,
         east_out_0__0__FORWARD__DATA__10_, east_out_0__0__FORWARD__DATA__9_,
         east_out_0__0__FORWARD__DATA__8_, east_out_0__0__FORWARD__DATA__7_,
         east_out_0__0__FORWARD__DATA__6_, east_out_0__0__FORWARD__DATA__5_,
         east_out_0__0__FORWARD__DATA__4_, east_out_0__0__FORWARD__DATA__3_,
         east_out_0__0__FORWARD__DATA__2_, east_out_0__0__FORWARD__DATA__1_,
         east_out_0__0__FORWARD__DATA__0_, east_out_0__1__FORWARD__REQ_,
         east_out_1__0__FORWARD__REQ_, east_out_1__0__FORWARD__DATA__34_,
         east_out_1__0__FORWARD__DATA__33_, east_out_1__0__FORWARD__DATA__32_,
         east_out_1__0__FORWARD__DATA__31_, east_out_1__0__FORWARD__DATA__30_,
         east_out_1__0__FORWARD__DATA__29_, east_out_1__0__FORWARD__DATA__28_,
         east_out_1__0__FORWARD__DATA__27_, east_out_1__0__FORWARD__DATA__26_,
         east_out_1__0__FORWARD__DATA__25_, east_out_1__0__FORWARD__DATA__24_,
         east_out_1__0__FORWARD__DATA__23_, east_out_1__0__FORWARD__DATA__22_,
         east_out_1__0__FORWARD__DATA__21_, east_out_1__0__FORWARD__DATA__20_,
         east_out_1__0__FORWARD__DATA__19_, east_out_1__0__FORWARD__DATA__18_,
         east_out_1__0__FORWARD__DATA__17_, east_out_1__0__FORWARD__DATA__16_,
         east_out_1__0__FORWARD__DATA__15_, east_out_1__0__FORWARD__DATA__14_,
         east_out_1__0__FORWARD__DATA__13_, east_out_1__0__FORWARD__DATA__12_,
         east_out_1__0__FORWARD__DATA__11_, east_out_1__0__FORWARD__DATA__10_,
         east_out_1__0__FORWARD__DATA__9_, east_out_1__0__FORWARD__DATA__8_,
         east_out_1__0__FORWARD__DATA__7_, east_out_1__0__FORWARD__DATA__6_,
         east_out_1__0__FORWARD__DATA__5_, east_out_1__0__FORWARD__DATA__4_,
         east_out_1__0__FORWARD__DATA__3_, east_out_1__0__FORWARD__DATA__2_,
         east_out_1__0__FORWARD__DATA__1_, east_out_1__0__FORWARD__DATA__0_,
         east_out_1__1__FORWARD__REQ_, east_out_1__1__FORWARD__DATA__34_,
         east_out_1__1__FORWARD__DATA__33_, east_out_1__1__FORWARD__DATA__32_,
         east_out_1__1__FORWARD__DATA__31_, east_out_1__1__FORWARD__DATA__30_,
         east_out_1__1__FORWARD__DATA__29_, east_out_1__1__FORWARD__DATA__28_,
         east_out_1__1__FORWARD__DATA__27_, east_out_1__1__FORWARD__DATA__26_,
         east_out_1__1__FORWARD__DATA__25_, east_out_1__1__FORWARD__DATA__24_,
         east_out_1__1__FORWARD__DATA__23_, east_out_1__1__FORWARD__DATA__22_,
         east_out_1__1__FORWARD__DATA__21_, east_out_1__1__FORWARD__DATA__20_,
         east_out_1__1__FORWARD__DATA__19_, east_out_1__1__FORWARD__DATA__18_,
         east_out_1__1__FORWARD__DATA__17_, east_out_1__1__FORWARD__DATA__16_,
         east_out_1__1__FORWARD__DATA__15_, east_out_1__1__FORWARD__DATA__14_,
         east_out_1__1__FORWARD__DATA__13_, east_out_1__1__FORWARD__DATA__12_,
         east_out_1__1__FORWARD__DATA__11_, east_out_1__1__FORWARD__DATA__10_,
         east_out_1__1__FORWARD__DATA__9_, east_out_1__1__FORWARD__DATA__8_,
         east_out_1__1__FORWARD__DATA__7_, east_out_1__1__FORWARD__DATA__6_,
         east_out_1__1__FORWARD__DATA__5_, east_out_1__1__FORWARD__DATA__4_,
         east_out_1__1__FORWARD__DATA__3_, east_out_1__1__FORWARD__DATA__2_,
         east_out_1__1__FORWARD__DATA__1_, east_out_1__1__FORWARD__DATA__0_,
         north_out_0__0__FORWARD__REQ_, north_out_0__1__FORWARD__REQ_,
         north_out_0__1__FORWARD__DATA__34_,
         north_out_0__1__FORWARD__DATA__33_,
         north_out_0__1__FORWARD__DATA__32_,
         north_out_0__1__FORWARD__DATA__31_,
         north_out_0__1__FORWARD__DATA__30_,
         north_out_0__1__FORWARD__DATA__29_,
         north_out_0__1__FORWARD__DATA__28_,
         north_out_0__1__FORWARD__DATA__27_,
         north_out_0__1__FORWARD__DATA__26_,
         north_out_0__1__FORWARD__DATA__25_,
         north_out_0__1__FORWARD__DATA__24_,
         north_out_0__1__FORWARD__DATA__23_,
         north_out_0__1__FORWARD__DATA__22_,
         north_out_0__1__FORWARD__DATA__21_,
         north_out_0__1__FORWARD__DATA__20_,
         north_out_0__1__FORWARD__DATA__19_,
         north_out_0__1__FORWARD__DATA__18_,
         north_out_0__1__FORWARD__DATA__17_,
         north_out_0__1__FORWARD__DATA__16_,
         north_out_0__1__FORWARD__DATA__15_,
         north_out_0__1__FORWARD__DATA__14_,
         north_out_0__1__FORWARD__DATA__13_,
         north_out_0__1__FORWARD__DATA__12_,
         north_out_0__1__FORWARD__DATA__11_,
         north_out_0__1__FORWARD__DATA__10_, north_out_0__1__FORWARD__DATA__9_,
         north_out_0__1__FORWARD__DATA__8_, north_out_0__1__FORWARD__DATA__7_,
         north_out_0__1__FORWARD__DATA__6_, north_out_0__1__FORWARD__DATA__5_,
         north_out_0__1__FORWARD__DATA__4_, north_out_0__1__FORWARD__DATA__3_,
         north_out_0__1__FORWARD__DATA__2_, north_out_0__1__FORWARD__DATA__1_,
         north_out_0__1__FORWARD__DATA__0_, north_out_1__0__FORWARD__REQ_,
         north_out_1__0__FORWARD__DATA__34_,
         north_out_1__0__FORWARD__DATA__33_,
         north_out_1__0__FORWARD__DATA__32_,
         north_out_1__0__FORWARD__DATA__31_,
         north_out_1__0__FORWARD__DATA__30_,
         north_out_1__0__FORWARD__DATA__29_,
         north_out_1__0__FORWARD__DATA__28_,
         north_out_1__0__FORWARD__DATA__27_,
         north_out_1__0__FORWARD__DATA__26_,
         north_out_1__0__FORWARD__DATA__25_,
         north_out_1__0__FORWARD__DATA__24_,
         north_out_1__0__FORWARD__DATA__23_,
         north_out_1__0__FORWARD__DATA__22_,
         north_out_1__0__FORWARD__DATA__21_,
         north_out_1__0__FORWARD__DATA__20_,
         north_out_1__0__FORWARD__DATA__19_,
         north_out_1__0__FORWARD__DATA__18_,
         north_out_1__0__FORWARD__DATA__17_,
         north_out_1__0__FORWARD__DATA__16_,
         north_out_1__0__FORWARD__DATA__15_,
         north_out_1__0__FORWARD__DATA__14_,
         north_out_1__0__FORWARD__DATA__13_,
         north_out_1__0__FORWARD__DATA__12_,
         north_out_1__0__FORWARD__DATA__11_,
         north_out_1__0__FORWARD__DATA__10_, north_out_1__0__FORWARD__DATA__9_,
         north_out_1__0__FORWARD__DATA__8_, north_out_1__0__FORWARD__DATA__7_,
         north_out_1__0__FORWARD__DATA__6_, north_out_1__0__FORWARD__DATA__5_,
         north_out_1__0__FORWARD__DATA__4_, north_out_1__0__FORWARD__DATA__3_,
         north_out_1__0__FORWARD__DATA__2_, north_out_1__0__FORWARD__DATA__1_,
         north_out_1__0__FORWARD__DATA__0_, north_out_1__1__FORWARD__REQ_,
         north_out_1__1__FORWARD__DATA__34_,
         north_out_1__1__FORWARD__DATA__33_,
         north_out_1__1__FORWARD__DATA__32_,
         north_out_1__1__FORWARD__DATA__31_,
         north_out_1__1__FORWARD__DATA__30_,
         north_out_1__1__FORWARD__DATA__29_,
         north_out_1__1__FORWARD__DATA__28_,
         north_out_1__1__FORWARD__DATA__27_,
         north_out_1__1__FORWARD__DATA__26_,
         north_out_1__1__FORWARD__DATA__25_,
         north_out_1__1__FORWARD__DATA__24_,
         north_out_1__1__FORWARD__DATA__23_,
         north_out_1__1__FORWARD__DATA__22_,
         north_out_1__1__FORWARD__DATA__21_,
         north_out_1__1__FORWARD__DATA__20_,
         north_out_1__1__FORWARD__DATA__19_,
         north_out_1__1__FORWARD__DATA__18_,
         north_out_1__1__FORWARD__DATA__17_,
         north_out_1__1__FORWARD__DATA__16_,
         north_out_1__1__FORWARD__DATA__15_,
         north_out_1__1__FORWARD__DATA__14_,
         north_out_1__1__FORWARD__DATA__13_,
         north_out_1__1__FORWARD__DATA__12_,
         north_out_1__1__FORWARD__DATA__11_,
         north_out_1__1__FORWARD__DATA__10_, north_out_1__1__FORWARD__DATA__9_,
         north_out_1__1__FORWARD__DATA__8_, north_out_1__1__FORWARD__DATA__7_,
         north_out_1__1__FORWARD__DATA__6_, north_out_1__1__FORWARD__DATA__5_,
         north_out_1__1__FORWARD__DATA__4_, north_out_1__1__FORWARD__DATA__3_,
         north_out_1__1__FORWARD__DATA__2_, north_out_1__1__FORWARD__DATA__1_,
         north_out_1__1__FORWARD__DATA__0_, west_in_0__0__FORWARD__DATA__34_,
         west_in_0__0__FORWARD__DATA__33_, west_in_0__0__FORWARD__DATA__32_,
         west_in_0__0__FORWARD__DATA__31_, west_in_0__0__FORWARD__DATA__30_,
         west_in_0__0__FORWARD__DATA__29_, west_in_0__0__FORWARD__DATA__28_,
         west_in_0__0__FORWARD__DATA__27_, west_in_0__0__FORWARD__DATA__26_,
         west_in_0__0__FORWARD__DATA__25_, west_in_0__0__FORWARD__DATA__24_,
         west_in_0__0__FORWARD__DATA__23_, west_in_0__0__FORWARD__DATA__22_,
         west_in_0__0__FORWARD__DATA__21_, west_in_0__0__FORWARD__DATA__20_,
         west_in_0__0__FORWARD__DATA__19_, west_in_0__0__FORWARD__DATA__18_,
         west_in_0__0__FORWARD__DATA__17_, west_in_0__0__FORWARD__DATA__16_,
         west_in_0__0__FORWARD__DATA__15_, west_in_0__0__FORWARD__DATA__14_,
         west_in_0__0__FORWARD__DATA__13_, west_in_0__0__FORWARD__DATA__12_,
         west_in_0__0__FORWARD__DATA__11_, west_in_0__0__FORWARD__DATA__10_,
         west_in_0__0__FORWARD__DATA__9_, west_in_0__0__FORWARD__DATA__8_,
         west_in_0__0__FORWARD__DATA__7_, west_in_0__0__FORWARD__DATA__6_,
         west_in_0__0__FORWARD__DATA__5_, west_in_0__0__FORWARD__DATA__4_,
         west_in_0__0__FORWARD__DATA__3_, west_in_0__0__FORWARD__DATA__2_,
         west_in_0__0__FORWARD__DATA__1_, west_in_0__0__FORWARD__DATA__0_,
         west_in_0__0__BACKWARD__ACK, west_in_0__1__BACKWARD__ACK,
         west_in_1__0__BACKWARD__ACK, west_in_1__1__BACKWARD__ACK,
         south_in_0__0__BACKWARD__ACK, south_in_0__1__BACKWARD__ACK,
         south_in_1__0__FORWARD__DATA__34_, south_in_1__0__FORWARD__DATA__33_,
         south_in_1__0__FORWARD__DATA__32_, south_in_1__0__FORWARD__DATA__31_,
         south_in_1__0__FORWARD__DATA__30_, south_in_1__0__FORWARD__DATA__29_,
         south_in_1__0__FORWARD__DATA__28_, south_in_1__0__FORWARD__DATA__27_,
         south_in_1__0__FORWARD__DATA__26_, south_in_1__0__FORWARD__DATA__25_,
         south_in_1__0__FORWARD__DATA__24_, south_in_1__0__FORWARD__DATA__23_,
         south_in_1__0__FORWARD__DATA__22_, south_in_1__0__FORWARD__DATA__21_,
         south_in_1__0__FORWARD__DATA__20_, south_in_1__0__FORWARD__DATA__19_,
         south_in_1__0__FORWARD__DATA__18_, south_in_1__0__FORWARD__DATA__17_,
         south_in_1__0__FORWARD__DATA__16_, south_in_1__0__FORWARD__DATA__15_,
         south_in_1__0__FORWARD__DATA__14_, south_in_1__0__FORWARD__DATA__13_,
         south_in_1__0__FORWARD__DATA__12_, south_in_1__0__FORWARD__DATA__11_,
         south_in_1__0__FORWARD__DATA__10_, south_in_1__0__FORWARD__DATA__9_,
         south_in_1__0__FORWARD__DATA__8_, south_in_1__0__FORWARD__DATA__7_,
         south_in_1__0__FORWARD__DATA__6_, south_in_1__0__FORWARD__DATA__5_,
         south_in_1__0__FORWARD__DATA__4_, south_in_1__0__FORWARD__DATA__3_,
         south_in_1__0__FORWARD__DATA__2_, south_in_1__0__FORWARD__DATA__1_,
         south_in_1__0__FORWARD__DATA__0_, south_in_1__0__BACKWARD__ACK,
         south_in_1__1__BACKWARD__ACK, east_in_0__0__BACKWARD__ACK,
         east_in_0__1__FORWARD__DATA__34_, east_in_0__1__FORWARD__DATA__33_,
         east_in_0__1__FORWARD__DATA__32_, east_in_0__1__FORWARD__DATA__31_,
         east_in_0__1__FORWARD__DATA__30_, east_in_0__1__FORWARD__DATA__29_,
         east_in_0__1__FORWARD__DATA__28_, east_in_0__1__FORWARD__DATA__27_,
         east_in_0__1__FORWARD__DATA__26_, east_in_0__1__FORWARD__DATA__25_,
         east_in_0__1__FORWARD__DATA__24_, east_in_0__1__FORWARD__DATA__23_,
         east_in_0__1__FORWARD__DATA__22_, east_in_0__1__FORWARD__DATA__21_,
         east_in_0__1__FORWARD__DATA__20_, east_in_0__1__FORWARD__DATA__19_,
         east_in_0__1__FORWARD__DATA__18_, east_in_0__1__FORWARD__DATA__17_,
         east_in_0__1__FORWARD__DATA__16_, east_in_0__1__FORWARD__DATA__15_,
         east_in_0__1__FORWARD__DATA__14_, east_in_0__1__FORWARD__DATA__13_,
         east_in_0__1__FORWARD__DATA__12_, east_in_0__1__FORWARD__DATA__11_,
         east_in_0__1__FORWARD__DATA__10_, east_in_0__1__FORWARD__DATA__9_,
         east_in_0__1__FORWARD__DATA__8_, east_in_0__1__FORWARD__DATA__7_,
         east_in_0__1__FORWARD__DATA__6_, east_in_0__1__FORWARD__DATA__5_,
         east_in_0__1__FORWARD__DATA__4_, east_in_0__1__FORWARD__DATA__3_,
         east_in_0__1__FORWARD__DATA__2_, east_in_0__1__FORWARD__DATA__1_,
         east_in_0__1__FORWARD__DATA__0_, east_in_0__1__BACKWARD__ACK,
         east_in_1__0__BACKWARD__ACK, east_in_1__1__BACKWARD__ACK,
         north_in_0__0__FORWARD__DATA__34_, north_in_0__0__FORWARD__DATA__33_,
         north_in_0__0__FORWARD__DATA__32_, north_in_0__0__FORWARD__DATA__31_,
         north_in_0__0__FORWARD__DATA__30_, north_in_0__0__FORWARD__DATA__29_,
         north_in_0__0__FORWARD__DATA__28_, north_in_0__0__FORWARD__DATA__27_,
         north_in_0__0__FORWARD__DATA__26_, north_in_0__0__FORWARD__DATA__25_,
         north_in_0__0__FORWARD__DATA__24_, north_in_0__0__FORWARD__DATA__23_,
         north_in_0__0__FORWARD__DATA__22_, north_in_0__0__FORWARD__DATA__21_,
         north_in_0__0__FORWARD__DATA__20_, north_in_0__0__FORWARD__DATA__19_,
         north_in_0__0__FORWARD__DATA__18_, north_in_0__0__FORWARD__DATA__17_,
         north_in_0__0__FORWARD__DATA__16_, north_in_0__0__FORWARD__DATA__15_,
         north_in_0__0__FORWARD__DATA__14_, north_in_0__0__FORWARD__DATA__13_,
         north_in_0__0__FORWARD__DATA__12_, north_in_0__0__FORWARD__DATA__11_,
         north_in_0__0__FORWARD__DATA__10_, north_in_0__0__FORWARD__DATA__9_,
         north_in_0__0__FORWARD__DATA__8_, north_in_0__0__FORWARD__DATA__7_,
         north_in_0__0__FORWARD__DATA__6_, north_in_0__0__FORWARD__DATA__5_,
         north_in_0__0__FORWARD__DATA__4_, north_in_0__0__FORWARD__DATA__3_,
         north_in_0__0__FORWARD__DATA__2_, north_in_0__0__FORWARD__DATA__1_,
         north_in_0__0__FORWARD__DATA__0_, north_in_0__0__BACKWARD__ACK,
         north_in_0__1__BACKWARD__ACK, north_in_1__0__BACKWARD__ACK,
         north_in_1__1__BACKWARD__ACK, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256;
  wire   [3:0] north_out_req0;
  wire   [3:0] north_out_req1;
  wire   [3:0] east_out_req0;
  wire   [3:0] east_out_req1;
  wire   [3:0] south_out_req0;
  wire   [3:0] south_out_req1;
  wire   [3:0] west_out_req0;
  wire   [3:0] west_out_req1;
  wire   [3:0] north_in_ack0;
  wire   [3:0] north_in_ack1;
  wire   [3:0] east_in_ack0;
  wire   [3:0] east_in_ack1;
  wire   [3:0] south_in_ack0;
  wire   [3:0] south_in_ack1;
  wire   [3:0] west_in_ack0;
  wire   [3:0] west_in_ack1;
  assign spm_ports_out[291] = 1'b0;
  assign spm_ports_out[290] = 1'b0;
  assign spm_ports_out[289] = 1'b0;
  assign spm_ports_out[288] = 1'b0;
  assign spm_ports_out[287] = 1'b0;
  assign spm_ports_out[286] = 1'b0;
  assign spm_ports_out[285] = 1'b0;
  assign spm_ports_out[284] = 1'b0;
  assign spm_ports_out[283] = 1'b0;
  assign spm_ports_out[282] = 1'b0;
  assign spm_ports_out[281] = 1'b0;
  assign spm_ports_out[280] = 1'b0;
  assign spm_ports_out[279] = 1'b0;
  assign spm_ports_out[278] = 1'b0;
  assign spm_ports_out[277] = 1'b0;
  assign spm_ports_out[276] = 1'b0;
  assign spm_ports_out[275] = 1'b0;
  assign spm_ports_out[193] = 1'b0;
  assign spm_ports_out[192] = 1'b0;
  assign spm_ports_out[191] = 1'b0;
  assign spm_ports_out[190] = 1'b0;
  assign spm_ports_out[189] = 1'b0;
  assign spm_ports_out[188] = 1'b0;
  assign spm_ports_out[187] = 1'b0;
  assign spm_ports_out[186] = 1'b0;
  assign spm_ports_out[185] = 1'b0;
  assign spm_ports_out[184] = 1'b0;
  assign spm_ports_out[183] = 1'b0;
  assign spm_ports_out[182] = 1'b0;
  assign spm_ports_out[181] = 1'b0;
  assign spm_ports_out[180] = 1'b0;
  assign spm_ports_out[179] = 1'b0;
  assign spm_ports_out[178] = 1'b0;
  assign spm_ports_out[177] = 1'b0;
  assign spm_ports_out[95] = 1'b0;
  assign spm_ports_out[94] = 1'b0;
  assign spm_ports_out[93] = 1'b0;
  assign spm_ports_out[92] = 1'b0;
  assign spm_ports_out[91] = 1'b0;
  assign spm_ports_out[90] = 1'b0;
  assign spm_ports_out[89] = 1'b0;
  assign spm_ports_out[88] = 1'b0;
  assign spm_ports_out[87] = 1'b0;
  assign spm_ports_out[86] = 1'b0;
  assign spm_ports_out[85] = 1'b0;
  assign spm_ports_out[84] = 1'b0;
  assign spm_ports_out[83] = 1'b0;
  assign spm_ports_out[82] = 1'b0;
  assign spm_ports_out[81] = 1'b0;
  assign spm_ports_out[80] = 1'b0;
  assign spm_ports_out[79] = 1'b0;
  assign spm_ports_out[389] = 1'b0;
  assign spm_ports_out[388] = 1'b0;
  assign spm_ports_out[387] = 1'b0;
  assign spm_ports_out[386] = 1'b0;
  assign spm_ports_out[385] = 1'b0;
  assign spm_ports_out[384] = 1'b0;
  assign spm_ports_out[383] = 1'b0;
  assign spm_ports_out[382] = 1'b0;
  assign spm_ports_out[381] = 1'b0;
  assign spm_ports_out[380] = 1'b0;
  assign spm_ports_out[379] = 1'b0;
  assign spm_ports_out[378] = 1'b0;
  assign spm_ports_out[377] = 1'b0;
  assign spm_ports_out[376] = 1'b0;
  assign spm_ports_out[375] = 1'b0;
  assign spm_ports_out[374] = 1'b0;
  assign spm_ports_out[373] = 1'b0;

  noc_node_0 node_1_1 ( .p_clk(p_clk), .n_clk(n_clk), .reset(reset), .proc_in(
        p_ports_in[263:198]), .proc_out(p_ports_out[135:102]), .spm_in(
        spm_ports_in[263:198]), .spm_out({spm_ports_out[391:390], 
        spm_ports_out_1__1__MADDR__31_, spm_ports_out_1__1__MADDR__30_, 
        spm_ports_out_1__1__MADDR__29_, spm_ports_out_1__1__MADDR__28_, 
        spm_ports_out_1__1__MADDR__27_, spm_ports_out_1__1__MADDR__26_, 
        spm_ports_out_1__1__MADDR__25_, spm_ports_out_1__1__MADDR__24_, 
        spm_ports_out_1__1__MADDR__23_, spm_ports_out_1__1__MADDR__22_, 
        spm_ports_out_1__1__MADDR__21_, spm_ports_out_1__1__MADDR__20_, 
        spm_ports_out_1__1__MADDR__19_, spm_ports_out_1__1__MADDR__18_, 
        spm_ports_out_1__1__MADDR__17_, spm_ports_out_1__1__MADDR__16_, n258, 
        spm_ports_out[372:294]}), .north_in_f({south_out_req1[2], 
        south_out_0__1__FORWARD__DATA__34_, south_out_0__1__FORWARD__DATA__33_, 
        south_out_0__1__FORWARD__DATA__32_, south_out_0__1__FORWARD__DATA__31_, 
        south_out_0__1__FORWARD__DATA__30_, south_out_0__1__FORWARD__DATA__29_, 
        south_out_0__1__FORWARD__DATA__28_, south_out_0__1__FORWARD__DATA__27_, 
        south_out_0__1__FORWARD__DATA__26_, south_out_0__1__FORWARD__DATA__25_, 
        south_out_0__1__FORWARD__DATA__24_, south_out_0__1__FORWARD__DATA__23_, 
        south_out_0__1__FORWARD__DATA__22_, south_out_0__1__FORWARD__DATA__21_, 
        south_out_0__1__FORWARD__DATA__20_, south_out_0__1__FORWARD__DATA__19_, 
        south_out_0__1__FORWARD__DATA__18_, south_out_0__1__FORWARD__DATA__17_, 
        south_out_0__1__FORWARD__DATA__16_, south_out_0__1__FORWARD__DATA__15_, 
        south_out_0__1__FORWARD__DATA__14_, south_out_0__1__FORWARD__DATA__13_, 
        south_out_0__1__FORWARD__DATA__12_, south_out_0__1__FORWARD__DATA__11_, 
        south_out_0__1__FORWARD__DATA__10_, south_out_0__1__FORWARD__DATA__9_, 
        south_out_0__1__FORWARD__DATA__8_, south_out_0__1__FORWARD__DATA__7_, 
        south_out_0__1__FORWARD__DATA__6_, south_out_0__1__FORWARD__DATA__5_, 
        south_out_0__1__FORWARD__DATA__4_, south_out_0__1__FORWARD__DATA__3_, 
        south_out_0__1__FORWARD__DATA__2_, south_out_0__1__FORWARD__DATA__1_, 
        south_out_0__1__FORWARD__DATA__0_}), .north_in_b(
        north_in_1__1__BACKWARD__ACK), .east_in_f({west_out_req1[1], 
        west_out_1__0__FORWARD__DATA__34_, west_out_1__0__FORWARD__DATA__33_, 
        west_out_1__0__FORWARD__DATA__32_, west_out_1__0__FORWARD__DATA__31_, 
        west_out_1__0__FORWARD__DATA__30_, west_out_1__0__FORWARD__DATA__29_, 
        west_out_1__0__FORWARD__DATA__28_, west_out_1__0__FORWARD__DATA__27_, 
        west_out_1__0__FORWARD__DATA__26_, west_out_1__0__FORWARD__DATA__25_, 
        west_out_1__0__FORWARD__DATA__24_, west_out_1__0__FORWARD__DATA__23_, 
        west_out_1__0__FORWARD__DATA__22_, west_out_1__0__FORWARD__DATA__21_, 
        west_out_1__0__FORWARD__DATA__20_, west_out_1__0__FORWARD__DATA__19_, 
        west_out_1__0__FORWARD__DATA__18_, west_out_1__0__FORWARD__DATA__17_, 
        west_out_1__0__FORWARD__DATA__16_, west_out_1__0__FORWARD__DATA__15_, 
        west_out_1__0__FORWARD__DATA__14_, west_out_1__0__FORWARD__DATA__13_, 
        west_out_1__0__FORWARD__DATA__12_, west_out_1__0__FORWARD__DATA__11_, 
        west_out_1__0__FORWARD__DATA__10_, west_out_1__0__FORWARD__DATA__9_, 
        west_out_1__0__FORWARD__DATA__8_, west_out_1__0__FORWARD__DATA__7_, 
        west_out_1__0__FORWARD__DATA__6_, west_out_1__0__FORWARD__DATA__5_, 
        west_out_1__0__FORWARD__DATA__4_, west_out_1__0__FORWARD__DATA__3_, 
        west_out_1__0__FORWARD__DATA__2_, west_out_1__0__FORWARD__DATA__1_, 
        west_out_1__0__FORWARD__DATA__0_}), .east_in_b(
        east_in_1__1__BACKWARD__ACK), .south_in_f({north_out_req1[2], 
        north_out_0__1__FORWARD__DATA__34_, north_out_0__1__FORWARD__DATA__33_, 
        north_out_0__1__FORWARD__DATA__32_, north_out_0__1__FORWARD__DATA__31_, 
        north_out_0__1__FORWARD__DATA__30_, north_out_0__1__FORWARD__DATA__29_, 
        north_out_0__1__FORWARD__DATA__28_, north_out_0__1__FORWARD__DATA__27_, 
        north_out_0__1__FORWARD__DATA__26_, north_out_0__1__FORWARD__DATA__25_, 
        north_out_0__1__FORWARD__DATA__24_, north_out_0__1__FORWARD__DATA__23_, 
        north_out_0__1__FORWARD__DATA__22_, north_out_0__1__FORWARD__DATA__21_, 
        north_out_0__1__FORWARD__DATA__20_, north_out_0__1__FORWARD__DATA__19_, 
        north_out_0__1__FORWARD__DATA__18_, north_out_0__1__FORWARD__DATA__17_, 
        north_out_0__1__FORWARD__DATA__16_, north_out_0__1__FORWARD__DATA__15_, 
        north_out_0__1__FORWARD__DATA__14_, north_out_0__1__FORWARD__DATA__13_, 
        north_out_0__1__FORWARD__DATA__12_, north_out_0__1__FORWARD__DATA__11_, 
        north_out_0__1__FORWARD__DATA__10_, north_out_0__1__FORWARD__DATA__9_, 
        north_out_0__1__FORWARD__DATA__8_, north_out_0__1__FORWARD__DATA__7_, 
        north_out_0__1__FORWARD__DATA__6_, north_out_0__1__FORWARD__DATA__5_, 
        north_out_0__1__FORWARD__DATA__4_, north_out_0__1__FORWARD__DATA__3_, 
        north_out_0__1__FORWARD__DATA__2_, north_out_0__1__FORWARD__DATA__1_, 
        north_out_0__1__FORWARD__DATA__0_}), .south_in_b(
        south_in_1__1__BACKWARD__ACK), .west_in_f({east_out_req1[1], 
        east_out_1__0__FORWARD__DATA__34_, east_out_1__0__FORWARD__DATA__33_, 
        east_out_1__0__FORWARD__DATA__32_, east_out_1__0__FORWARD__DATA__31_, 
        east_out_1__0__FORWARD__DATA__30_, east_out_1__0__FORWARD__DATA__29_, 
        east_out_1__0__FORWARD__DATA__28_, east_out_1__0__FORWARD__DATA__27_, 
        east_out_1__0__FORWARD__DATA__26_, east_out_1__0__FORWARD__DATA__25_, 
        east_out_1__0__FORWARD__DATA__24_, east_out_1__0__FORWARD__DATA__23_, 
        east_out_1__0__FORWARD__DATA__22_, east_out_1__0__FORWARD__DATA__21_, 
        east_out_1__0__FORWARD__DATA__20_, east_out_1__0__FORWARD__DATA__19_, 
        east_out_1__0__FORWARD__DATA__18_, east_out_1__0__FORWARD__DATA__17_, 
        east_out_1__0__FORWARD__DATA__16_, east_out_1__0__FORWARD__DATA__15_, 
        east_out_1__0__FORWARD__DATA__14_, east_out_1__0__FORWARD__DATA__13_, 
        east_out_1__0__FORWARD__DATA__12_, east_out_1__0__FORWARD__DATA__11_, 
        east_out_1__0__FORWARD__DATA__10_, east_out_1__0__FORWARD__DATA__9_, 
        east_out_1__0__FORWARD__DATA__8_, east_out_1__0__FORWARD__DATA__7_, 
        east_out_1__0__FORWARD__DATA__6_, east_out_1__0__FORWARD__DATA__5_, 
        east_out_1__0__FORWARD__DATA__4_, east_out_1__0__FORWARD__DATA__3_, 
        east_out_1__0__FORWARD__DATA__2_, east_out_1__0__FORWARD__DATA__1_, 
        east_out_1__0__FORWARD__DATA__0_}), .west_in_b(
        west_in_1__1__BACKWARD__ACK), .north_out_f({
        north_out_1__1__FORWARD__REQ_, north_out_1__1__FORWARD__DATA__34_, 
        north_out_1__1__FORWARD__DATA__33_, north_out_1__1__FORWARD__DATA__32_, 
        north_out_1__1__FORWARD__DATA__31_, north_out_1__1__FORWARD__DATA__30_, 
        north_out_1__1__FORWARD__DATA__29_, north_out_1__1__FORWARD__DATA__28_, 
        north_out_1__1__FORWARD__DATA__27_, north_out_1__1__FORWARD__DATA__26_, 
        north_out_1__1__FORWARD__DATA__25_, north_out_1__1__FORWARD__DATA__24_, 
        north_out_1__1__FORWARD__DATA__23_, north_out_1__1__FORWARD__DATA__22_, 
        north_out_1__1__FORWARD__DATA__21_, north_out_1__1__FORWARD__DATA__20_, 
        north_out_1__1__FORWARD__DATA__19_, north_out_1__1__FORWARD__DATA__18_, 
        north_out_1__1__FORWARD__DATA__17_, north_out_1__1__FORWARD__DATA__16_, 
        north_out_1__1__FORWARD__DATA__15_, north_out_1__1__FORWARD__DATA__14_, 
        north_out_1__1__FORWARD__DATA__13_, north_out_1__1__FORWARD__DATA__12_, 
        north_out_1__1__FORWARD__DATA__11_, north_out_1__1__FORWARD__DATA__10_, 
        north_out_1__1__FORWARD__DATA__9_, north_out_1__1__FORWARD__DATA__8_, 
        north_out_1__1__FORWARD__DATA__7_, north_out_1__1__FORWARD__DATA__6_, 
        north_out_1__1__FORWARD__DATA__5_, north_out_1__1__FORWARD__DATA__4_, 
        north_out_1__1__FORWARD__DATA__3_, north_out_1__1__FORWARD__DATA__2_, 
        north_out_1__1__FORWARD__DATA__1_, north_out_1__1__FORWARD__DATA__0_}), 
        .north_out_b(south_in_ack1[2]), .east_out_f({
        east_out_1__1__FORWARD__REQ_, east_out_1__1__FORWARD__DATA__34_, 
        east_out_1__1__FORWARD__DATA__33_, east_out_1__1__FORWARD__DATA__32_, 
        east_out_1__1__FORWARD__DATA__31_, east_out_1__1__FORWARD__DATA__30_, 
        east_out_1__1__FORWARD__DATA__29_, east_out_1__1__FORWARD__DATA__28_, 
        east_out_1__1__FORWARD__DATA__27_, east_out_1__1__FORWARD__DATA__26_, 
        east_out_1__1__FORWARD__DATA__25_, east_out_1__1__FORWARD__DATA__24_, 
        east_out_1__1__FORWARD__DATA__23_, east_out_1__1__FORWARD__DATA__22_, 
        east_out_1__1__FORWARD__DATA__21_, east_out_1__1__FORWARD__DATA__20_, 
        east_out_1__1__FORWARD__DATA__19_, east_out_1__1__FORWARD__DATA__18_, 
        east_out_1__1__FORWARD__DATA__17_, east_out_1__1__FORWARD__DATA__16_, 
        east_out_1__1__FORWARD__DATA__15_, east_out_1__1__FORWARD__DATA__14_, 
        east_out_1__1__FORWARD__DATA__13_, east_out_1__1__FORWARD__DATA__12_, 
        east_out_1__1__FORWARD__DATA__11_, east_out_1__1__FORWARD__DATA__10_, 
        east_out_1__1__FORWARD__DATA__9_, east_out_1__1__FORWARD__DATA__8_, 
        east_out_1__1__FORWARD__DATA__7_, east_out_1__1__FORWARD__DATA__6_, 
        east_out_1__1__FORWARD__DATA__5_, east_out_1__1__FORWARD__DATA__4_, 
        east_out_1__1__FORWARD__DATA__3_, east_out_1__1__FORWARD__DATA__2_, 
        east_out_1__1__FORWARD__DATA__1_, east_out_1__1__FORWARD__DATA__0_}), 
        .east_out_b(west_in_ack1[1]), .south_out_f({
        south_out_1__1__FORWARD__REQ_, south_out_1__1__FORWARD__DATA__34_, 
        south_out_1__1__FORWARD__DATA__33_, south_out_1__1__FORWARD__DATA__32_, 
        south_out_1__1__FORWARD__DATA__31_, south_out_1__1__FORWARD__DATA__30_, 
        south_out_1__1__FORWARD__DATA__29_, south_out_1__1__FORWARD__DATA__28_, 
        south_out_1__1__FORWARD__DATA__27_, south_out_1__1__FORWARD__DATA__26_, 
        south_out_1__1__FORWARD__DATA__25_, south_out_1__1__FORWARD__DATA__24_, 
        south_out_1__1__FORWARD__DATA__23_, south_out_1__1__FORWARD__DATA__22_, 
        south_out_1__1__FORWARD__DATA__21_, south_out_1__1__FORWARD__DATA__20_, 
        south_out_1__1__FORWARD__DATA__19_, south_out_1__1__FORWARD__DATA__18_, 
        south_out_1__1__FORWARD__DATA__17_, south_out_1__1__FORWARD__DATA__16_, 
        south_out_1__1__FORWARD__DATA__15_, south_out_1__1__FORWARD__DATA__14_, 
        south_out_1__1__FORWARD__DATA__13_, south_out_1__1__FORWARD__DATA__12_, 
        south_out_1__1__FORWARD__DATA__11_, south_out_1__1__FORWARD__DATA__10_, 
        south_out_1__1__FORWARD__DATA__9_, south_out_1__1__FORWARD__DATA__8_, 
        south_out_1__1__FORWARD__DATA__7_, south_out_1__1__FORWARD__DATA__6_, 
        south_out_1__1__FORWARD__DATA__5_, south_out_1__1__FORWARD__DATA__4_, 
        south_out_1__1__FORWARD__DATA__3_, south_out_1__1__FORWARD__DATA__2_, 
        south_out_1__1__FORWARD__DATA__1_, south_out_1__1__FORWARD__DATA__0_}), 
        .south_out_b(north_in_ack1[2]), .west_out_f({
        west_out_1__1__FORWARD__REQ_, west_out_1__1__FORWARD__DATA__34_, 
        west_out_1__1__FORWARD__DATA__33_, west_out_1__1__FORWARD__DATA__32_, 
        west_out_1__1__FORWARD__DATA__31_, west_out_1__1__FORWARD__DATA__30_, 
        west_out_1__1__FORWARD__DATA__29_, west_out_1__1__FORWARD__DATA__28_, 
        west_out_1__1__FORWARD__DATA__27_, west_out_1__1__FORWARD__DATA__26_, 
        west_out_1__1__FORWARD__DATA__25_, west_out_1__1__FORWARD__DATA__24_, 
        west_out_1__1__FORWARD__DATA__23_, west_out_1__1__FORWARD__DATA__22_, 
        west_out_1__1__FORWARD__DATA__21_, west_out_1__1__FORWARD__DATA__20_, 
        west_out_1__1__FORWARD__DATA__19_, west_out_1__1__FORWARD__DATA__18_, 
        west_out_1__1__FORWARD__DATA__17_, west_out_1__1__FORWARD__DATA__16_, 
        west_out_1__1__FORWARD__DATA__15_, west_out_1__1__FORWARD__DATA__14_, 
        west_out_1__1__FORWARD__DATA__13_, west_out_1__1__FORWARD__DATA__12_, 
        west_out_1__1__FORWARD__DATA__11_, west_out_1__1__FORWARD__DATA__10_, 
        west_out_1__1__FORWARD__DATA__9_, west_out_1__1__FORWARD__DATA__8_, 
        west_out_1__1__FORWARD__DATA__7_, west_out_1__1__FORWARD__DATA__6_, 
        west_out_1__1__FORWARD__DATA__5_, west_out_1__1__FORWARD__DATA__4_, 
        west_out_1__1__FORWARD__DATA__3_, west_out_1__1__FORWARD__DATA__2_, 
        west_out_1__1__FORWARD__DATA__1_, west_out_1__1__FORWARD__DATA__0_}), 
        .west_out_b(east_in_ack1[1]) );
  noc_node_3 node_1_0 ( .p_clk(p_clk), .n_clk(n_clk), .reset(reset), .proc_in(
        p_ports_in[197:132]), .proc_out(p_ports_out[101:68]), .spm_in(
        spm_ports_in[197:132]), .spm_out({spm_ports_out[293:292], 
        spm_ports_out_1__0__MADDR__31_, spm_ports_out_1__0__MADDR__30_, 
        spm_ports_out_1__0__MADDR__29_, spm_ports_out_1__0__MADDR__28_, 
        spm_ports_out_1__0__MADDR__27_, spm_ports_out_1__0__MADDR__26_, 
        spm_ports_out_1__0__MADDR__25_, spm_ports_out_1__0__MADDR__24_, 
        spm_ports_out_1__0__MADDR__23_, spm_ports_out_1__0__MADDR__22_, 
        spm_ports_out_1__0__MADDR__21_, spm_ports_out_1__0__MADDR__20_, 
        spm_ports_out_1__0__MADDR__19_, spm_ports_out_1__0__MADDR__18_, 
        spm_ports_out_1__0__MADDR__17_, spm_ports_out_1__0__MADDR__16_, 
        spm_ports_out_1__0__MADDR__15_, spm_ports_out[274:196]}), .north_in_f(
        {south_out_req1[3], south_out_0__0__FORWARD__DATA__34_, 
        south_out_0__0__FORWARD__DATA__33_, south_out_0__0__FORWARD__DATA__32_, 
        south_out_0__0__FORWARD__DATA__31_, south_out_0__0__FORWARD__DATA__30_, 
        south_out_0__0__FORWARD__DATA__29_, south_out_0__0__FORWARD__DATA__28_, 
        south_out_0__0__FORWARD__DATA__27_, south_out_0__0__FORWARD__DATA__26_, 
        south_out_0__0__FORWARD__DATA__25_, south_out_0__0__FORWARD__DATA__24_, 
        south_out_0__0__FORWARD__DATA__23_, south_out_0__0__FORWARD__DATA__22_, 
        south_out_0__0__FORWARD__DATA__21_, south_out_0__0__FORWARD__DATA__20_, 
        south_out_0__0__FORWARD__DATA__19_, south_out_0__0__FORWARD__DATA__18_, 
        south_out_0__0__FORWARD__DATA__17_, south_out_0__0__FORWARD__DATA__16_, 
        south_out_0__0__FORWARD__DATA__15_, south_out_0__0__FORWARD__DATA__14_, 
        south_out_0__0__FORWARD__DATA__13_, south_out_0__0__FORWARD__DATA__12_, 
        south_out_0__0__FORWARD__DATA__11_, south_out_0__0__FORWARD__DATA__10_, 
        south_out_0__0__FORWARD__DATA__9_, south_out_0__0__FORWARD__DATA__8_, 
        south_out_0__0__FORWARD__DATA__7_, south_out_0__0__FORWARD__DATA__6_, 
        south_out_0__0__FORWARD__DATA__5_, south_out_0__0__FORWARD__DATA__4_, 
        south_out_0__0__FORWARD__DATA__3_, south_out_0__0__FORWARD__DATA__2_, 
        south_out_0__0__FORWARD__DATA__1_, south_out_0__0__FORWARD__DATA__0_}), 
        .north_in_b(north_in_1__0__BACKWARD__ACK), .east_in_f({
        west_out_req1[0], west_out_1__1__FORWARD__DATA__34_, 
        west_out_1__1__FORWARD__DATA__33_, west_out_1__1__FORWARD__DATA__32_, 
        west_out_1__1__FORWARD__DATA__31_, west_out_1__1__FORWARD__DATA__30_, 
        west_out_1__1__FORWARD__DATA__29_, west_out_1__1__FORWARD__DATA__28_, 
        west_out_1__1__FORWARD__DATA__27_, west_out_1__1__FORWARD__DATA__26_, 
        west_out_1__1__FORWARD__DATA__25_, west_out_1__1__FORWARD__DATA__24_, 
        west_out_1__1__FORWARD__DATA__23_, west_out_1__1__FORWARD__DATA__22_, 
        west_out_1__1__FORWARD__DATA__21_, west_out_1__1__FORWARD__DATA__20_, 
        west_out_1__1__FORWARD__DATA__19_, west_out_1__1__FORWARD__DATA__18_, 
        west_out_1__1__FORWARD__DATA__17_, west_out_1__1__FORWARD__DATA__16_, 
        west_out_1__1__FORWARD__DATA__15_, west_out_1__1__FORWARD__DATA__14_, 
        west_out_1__1__FORWARD__DATA__13_, west_out_1__1__FORWARD__DATA__12_, 
        west_out_1__1__FORWARD__DATA__11_, west_out_1__1__FORWARD__DATA__10_, 
        west_out_1__1__FORWARD__DATA__9_, west_out_1__1__FORWARD__DATA__8_, 
        west_out_1__1__FORWARD__DATA__7_, west_out_1__1__FORWARD__DATA__6_, 
        west_out_1__1__FORWARD__DATA__5_, west_out_1__1__FORWARD__DATA__4_, 
        west_out_1__1__FORWARD__DATA__3_, west_out_1__1__FORWARD__DATA__2_, 
        west_out_1__1__FORWARD__DATA__1_, west_out_1__1__FORWARD__DATA__0_}), 
        .east_in_b(east_in_1__0__BACKWARD__ACK), .south_in_f({
        north_out_req1[3], south_in_1__0__FORWARD__DATA__34_, 
        south_in_1__0__FORWARD__DATA__33_, south_in_1__0__FORWARD__DATA__32_, 
        south_in_1__0__FORWARD__DATA__31_, south_in_1__0__FORWARD__DATA__30_, 
        south_in_1__0__FORWARD__DATA__29_, south_in_1__0__FORWARD__DATA__28_, 
        south_in_1__0__FORWARD__DATA__27_, south_in_1__0__FORWARD__DATA__26_, 
        south_in_1__0__FORWARD__DATA__25_, south_in_1__0__FORWARD__DATA__24_, 
        south_in_1__0__FORWARD__DATA__23_, south_in_1__0__FORWARD__DATA__22_, 
        south_in_1__0__FORWARD__DATA__21_, south_in_1__0__FORWARD__DATA__20_, 
        south_in_1__0__FORWARD__DATA__19_, south_in_1__0__FORWARD__DATA__18_, 
        south_in_1__0__FORWARD__DATA__17_, south_in_1__0__FORWARD__DATA__16_, 
        south_in_1__0__FORWARD__DATA__15_, south_in_1__0__FORWARD__DATA__14_, 
        south_in_1__0__FORWARD__DATA__13_, south_in_1__0__FORWARD__DATA__12_, 
        south_in_1__0__FORWARD__DATA__11_, south_in_1__0__FORWARD__DATA__10_, 
        south_in_1__0__FORWARD__DATA__9_, south_in_1__0__FORWARD__DATA__8_, 
        south_in_1__0__FORWARD__DATA__7_, south_in_1__0__FORWARD__DATA__6_, 
        south_in_1__0__FORWARD__DATA__5_, south_in_1__0__FORWARD__DATA__4_, 
        south_in_1__0__FORWARD__DATA__3_, south_in_1__0__FORWARD__DATA__2_, 
        south_in_1__0__FORWARD__DATA__1_, south_in_1__0__FORWARD__DATA__0_}), 
        .south_in_b(south_in_1__0__BACKWARD__ACK), .west_in_f({
        east_out_req1[0], east_out_1__1__FORWARD__DATA__34_, 
        east_out_1__1__FORWARD__DATA__33_, east_out_1__1__FORWARD__DATA__32_, 
        east_out_1__1__FORWARD__DATA__31_, east_out_1__1__FORWARD__DATA__30_, 
        east_out_1__1__FORWARD__DATA__29_, east_out_1__1__FORWARD__DATA__28_, 
        east_out_1__1__FORWARD__DATA__27_, east_out_1__1__FORWARD__DATA__26_, 
        east_out_1__1__FORWARD__DATA__25_, east_out_1__1__FORWARD__DATA__24_, 
        east_out_1__1__FORWARD__DATA__23_, east_out_1__1__FORWARD__DATA__22_, 
        east_out_1__1__FORWARD__DATA__21_, east_out_1__1__FORWARD__DATA__20_, 
        east_out_1__1__FORWARD__DATA__19_, east_out_1__1__FORWARD__DATA__18_, 
        east_out_1__1__FORWARD__DATA__17_, east_out_1__1__FORWARD__DATA__16_, 
        east_out_1__1__FORWARD__DATA__15_, east_out_1__1__FORWARD__DATA__14_, 
        east_out_1__1__FORWARD__DATA__13_, east_out_1__1__FORWARD__DATA__12_, 
        east_out_1__1__FORWARD__DATA__11_, east_out_1__1__FORWARD__DATA__10_, 
        east_out_1__1__FORWARD__DATA__9_, east_out_1__1__FORWARD__DATA__8_, 
        east_out_1__1__FORWARD__DATA__7_, east_out_1__1__FORWARD__DATA__6_, 
        east_out_1__1__FORWARD__DATA__5_, east_out_1__1__FORWARD__DATA__4_, 
        east_out_1__1__FORWARD__DATA__3_, east_out_1__1__FORWARD__DATA__2_, 
        east_out_1__1__FORWARD__DATA__1_, east_out_1__1__FORWARD__DATA__0_}), 
        .west_in_b(west_in_1__0__BACKWARD__ACK), .north_out_f({
        north_out_1__0__FORWARD__REQ_, north_out_1__0__FORWARD__DATA__34_, 
        north_out_1__0__FORWARD__DATA__33_, north_out_1__0__FORWARD__DATA__32_, 
        north_out_1__0__FORWARD__DATA__31_, north_out_1__0__FORWARD__DATA__30_, 
        north_out_1__0__FORWARD__DATA__29_, north_out_1__0__FORWARD__DATA__28_, 
        north_out_1__0__FORWARD__DATA__27_, north_out_1__0__FORWARD__DATA__26_, 
        north_out_1__0__FORWARD__DATA__25_, north_out_1__0__FORWARD__DATA__24_, 
        north_out_1__0__FORWARD__DATA__23_, north_out_1__0__FORWARD__DATA__22_, 
        north_out_1__0__FORWARD__DATA__21_, north_out_1__0__FORWARD__DATA__20_, 
        north_out_1__0__FORWARD__DATA__19_, north_out_1__0__FORWARD__DATA__18_, 
        north_out_1__0__FORWARD__DATA__17_, north_out_1__0__FORWARD__DATA__16_, 
        north_out_1__0__FORWARD__DATA__15_, north_out_1__0__FORWARD__DATA__14_, 
        north_out_1__0__FORWARD__DATA__13_, north_out_1__0__FORWARD__DATA__12_, 
        north_out_1__0__FORWARD__DATA__11_, north_out_1__0__FORWARD__DATA__10_, 
        north_out_1__0__FORWARD__DATA__9_, north_out_1__0__FORWARD__DATA__8_, 
        north_out_1__0__FORWARD__DATA__7_, north_out_1__0__FORWARD__DATA__6_, 
        north_out_1__0__FORWARD__DATA__5_, north_out_1__0__FORWARD__DATA__4_, 
        north_out_1__0__FORWARD__DATA__3_, north_out_1__0__FORWARD__DATA__2_, 
        north_out_1__0__FORWARD__DATA__1_, north_out_1__0__FORWARD__DATA__0_}), 
        .north_out_b(south_in_ack1[3]), .east_out_f({
        east_out_1__0__FORWARD__REQ_, east_out_1__0__FORWARD__DATA__34_, 
        east_out_1__0__FORWARD__DATA__33_, east_out_1__0__FORWARD__DATA__32_, 
        east_out_1__0__FORWARD__DATA__31_, east_out_1__0__FORWARD__DATA__30_, 
        east_out_1__0__FORWARD__DATA__29_, east_out_1__0__FORWARD__DATA__28_, 
        east_out_1__0__FORWARD__DATA__27_, east_out_1__0__FORWARD__DATA__26_, 
        east_out_1__0__FORWARD__DATA__25_, east_out_1__0__FORWARD__DATA__24_, 
        east_out_1__0__FORWARD__DATA__23_, east_out_1__0__FORWARD__DATA__22_, 
        east_out_1__0__FORWARD__DATA__21_, east_out_1__0__FORWARD__DATA__20_, 
        east_out_1__0__FORWARD__DATA__19_, east_out_1__0__FORWARD__DATA__18_, 
        east_out_1__0__FORWARD__DATA__17_, east_out_1__0__FORWARD__DATA__16_, 
        east_out_1__0__FORWARD__DATA__15_, east_out_1__0__FORWARD__DATA__14_, 
        east_out_1__0__FORWARD__DATA__13_, east_out_1__0__FORWARD__DATA__12_, 
        east_out_1__0__FORWARD__DATA__11_, east_out_1__0__FORWARD__DATA__10_, 
        east_out_1__0__FORWARD__DATA__9_, east_out_1__0__FORWARD__DATA__8_, 
        east_out_1__0__FORWARD__DATA__7_, east_out_1__0__FORWARD__DATA__6_, 
        east_out_1__0__FORWARD__DATA__5_, east_out_1__0__FORWARD__DATA__4_, 
        east_out_1__0__FORWARD__DATA__3_, east_out_1__0__FORWARD__DATA__2_, 
        east_out_1__0__FORWARD__DATA__1_, east_out_1__0__FORWARD__DATA__0_}), 
        .east_out_b(west_in_ack1[0]), .south_out_f({
        south_out_1__0__FORWARD__REQ_, north_in_0__0__FORWARD__DATA__34_, 
        north_in_0__0__FORWARD__DATA__33_, north_in_0__0__FORWARD__DATA__32_, 
        north_in_0__0__FORWARD__DATA__31_, north_in_0__0__FORWARD__DATA__30_, 
        north_in_0__0__FORWARD__DATA__29_, north_in_0__0__FORWARD__DATA__28_, 
        north_in_0__0__FORWARD__DATA__27_, north_in_0__0__FORWARD__DATA__26_, 
        north_in_0__0__FORWARD__DATA__25_, north_in_0__0__FORWARD__DATA__24_, 
        north_in_0__0__FORWARD__DATA__23_, north_in_0__0__FORWARD__DATA__22_, 
        north_in_0__0__FORWARD__DATA__21_, north_in_0__0__FORWARD__DATA__20_, 
        north_in_0__0__FORWARD__DATA__19_, north_in_0__0__FORWARD__DATA__18_, 
        north_in_0__0__FORWARD__DATA__17_, north_in_0__0__FORWARD__DATA__16_, 
        north_in_0__0__FORWARD__DATA__15_, north_in_0__0__FORWARD__DATA__14_, 
        north_in_0__0__FORWARD__DATA__13_, north_in_0__0__FORWARD__DATA__12_, 
        north_in_0__0__FORWARD__DATA__11_, north_in_0__0__FORWARD__DATA__10_, 
        north_in_0__0__FORWARD__DATA__9_, north_in_0__0__FORWARD__DATA__8_, 
        north_in_0__0__FORWARD__DATA__7_, north_in_0__0__FORWARD__DATA__6_, 
        north_in_0__0__FORWARD__DATA__5_, north_in_0__0__FORWARD__DATA__4_, 
        north_in_0__0__FORWARD__DATA__3_, north_in_0__0__FORWARD__DATA__2_, 
        north_in_0__0__FORWARD__DATA__1_, north_in_0__0__FORWARD__DATA__0_}), 
        .south_out_b(north_in_ack1[3]), .west_out_f({
        west_out_1__0__FORWARD__REQ_, west_out_1__0__FORWARD__DATA__34_, 
        west_out_1__0__FORWARD__DATA__33_, west_out_1__0__FORWARD__DATA__32_, 
        west_out_1__0__FORWARD__DATA__31_, west_out_1__0__FORWARD__DATA__30_, 
        west_out_1__0__FORWARD__DATA__29_, west_out_1__0__FORWARD__DATA__28_, 
        west_out_1__0__FORWARD__DATA__27_, west_out_1__0__FORWARD__DATA__26_, 
        west_out_1__0__FORWARD__DATA__25_, west_out_1__0__FORWARD__DATA__24_, 
        west_out_1__0__FORWARD__DATA__23_, west_out_1__0__FORWARD__DATA__22_, 
        west_out_1__0__FORWARD__DATA__21_, west_out_1__0__FORWARD__DATA__20_, 
        west_out_1__0__FORWARD__DATA__19_, west_out_1__0__FORWARD__DATA__18_, 
        west_out_1__0__FORWARD__DATA__17_, west_out_1__0__FORWARD__DATA__16_, 
        west_out_1__0__FORWARD__DATA__15_, west_out_1__0__FORWARD__DATA__14_, 
        west_out_1__0__FORWARD__DATA__13_, west_out_1__0__FORWARD__DATA__12_, 
        west_out_1__0__FORWARD__DATA__11_, west_out_1__0__FORWARD__DATA__10_, 
        west_out_1__0__FORWARD__DATA__9_, west_out_1__0__FORWARD__DATA__8_, 
        west_out_1__0__FORWARD__DATA__7_, west_out_1__0__FORWARD__DATA__6_, 
        west_out_1__0__FORWARD__DATA__5_, west_out_1__0__FORWARD__DATA__4_, 
        west_out_1__0__FORWARD__DATA__3_, west_out_1__0__FORWARD__DATA__2_, 
        west_out_1__0__FORWARD__DATA__1_, west_out_1__0__FORWARD__DATA__0_}), 
        .west_out_b(east_in_ack1[0]) );
  noc_node_2 node_0_1 ( .p_clk(p_clk), .n_clk(n_clk), .reset(reset), .proc_in(
        p_ports_in[131:66]), .proc_out(p_ports_out[67:34]), .spm_in(
        spm_ports_in[131:66]), .spm_out({spm_ports_out[195:194], 
        spm_ports_out_0__1__MADDR__31_, spm_ports_out_0__1__MADDR__30_, 
        spm_ports_out_0__1__MADDR__29_, spm_ports_out_0__1__MADDR__28_, 
        spm_ports_out_0__1__MADDR__27_, spm_ports_out_0__1__MADDR__26_, 
        spm_ports_out_0__1__MADDR__25_, spm_ports_out_0__1__MADDR__24_, 
        spm_ports_out_0__1__MADDR__23_, spm_ports_out_0__1__MADDR__22_, 
        spm_ports_out_0__1__MADDR__21_, spm_ports_out_0__1__MADDR__20_, 
        spm_ports_out_0__1__MADDR__19_, spm_ports_out_0__1__MADDR__18_, 
        spm_ports_out_0__1__MADDR__17_, spm_ports_out_0__1__MADDR__16_, 
        spm_ports_out_0__1__MADDR__15_, spm_ports_out[176:98]}), .north_in_f({
        south_out_req1[0], south_out_1__1__FORWARD__DATA__34_, 
        south_out_1__1__FORWARD__DATA__33_, south_out_1__1__FORWARD__DATA__32_, 
        south_out_1__1__FORWARD__DATA__31_, south_out_1__1__FORWARD__DATA__30_, 
        south_out_1__1__FORWARD__DATA__29_, south_out_1__1__FORWARD__DATA__28_, 
        south_out_1__1__FORWARD__DATA__27_, south_out_1__1__FORWARD__DATA__26_, 
        south_out_1__1__FORWARD__DATA__25_, south_out_1__1__FORWARD__DATA__24_, 
        south_out_1__1__FORWARD__DATA__23_, south_out_1__1__FORWARD__DATA__22_, 
        south_out_1__1__FORWARD__DATA__21_, south_out_1__1__FORWARD__DATA__20_, 
        south_out_1__1__FORWARD__DATA__19_, south_out_1__1__FORWARD__DATA__18_, 
        south_out_1__1__FORWARD__DATA__17_, south_out_1__1__FORWARD__DATA__16_, 
        south_out_1__1__FORWARD__DATA__15_, south_out_1__1__FORWARD__DATA__14_, 
        south_out_1__1__FORWARD__DATA__13_, south_out_1__1__FORWARD__DATA__12_, 
        south_out_1__1__FORWARD__DATA__11_, south_out_1__1__FORWARD__DATA__10_, 
        south_out_1__1__FORWARD__DATA__9_, south_out_1__1__FORWARD__DATA__8_, 
        south_out_1__1__FORWARD__DATA__7_, south_out_1__1__FORWARD__DATA__6_, 
        south_out_1__1__FORWARD__DATA__5_, south_out_1__1__FORWARD__DATA__4_, 
        south_out_1__1__FORWARD__DATA__3_, south_out_1__1__FORWARD__DATA__2_, 
        south_out_1__1__FORWARD__DATA__1_, south_out_1__1__FORWARD__DATA__0_}), 
        .north_in_b(north_in_0__1__BACKWARD__ACK), .east_in_f({
        west_out_req1[3], east_in_0__1__FORWARD__DATA__34_, 
        east_in_0__1__FORWARD__DATA__33_, east_in_0__1__FORWARD__DATA__32_, 
        east_in_0__1__FORWARD__DATA__31_, east_in_0__1__FORWARD__DATA__30_, 
        east_in_0__1__FORWARD__DATA__29_, east_in_0__1__FORWARD__DATA__28_, 
        east_in_0__1__FORWARD__DATA__27_, east_in_0__1__FORWARD__DATA__26_, 
        east_in_0__1__FORWARD__DATA__25_, east_in_0__1__FORWARD__DATA__24_, 
        east_in_0__1__FORWARD__DATA__23_, east_in_0__1__FORWARD__DATA__22_, 
        east_in_0__1__FORWARD__DATA__21_, east_in_0__1__FORWARD__DATA__20_, 
        east_in_0__1__FORWARD__DATA__19_, east_in_0__1__FORWARD__DATA__18_, 
        east_in_0__1__FORWARD__DATA__17_, east_in_0__1__FORWARD__DATA__16_, 
        east_in_0__1__FORWARD__DATA__15_, east_in_0__1__FORWARD__DATA__14_, 
        east_in_0__1__FORWARD__DATA__13_, east_in_0__1__FORWARD__DATA__12_, 
        east_in_0__1__FORWARD__DATA__11_, east_in_0__1__FORWARD__DATA__10_, 
        east_in_0__1__FORWARD__DATA__9_, east_in_0__1__FORWARD__DATA__8_, 
        east_in_0__1__FORWARD__DATA__7_, east_in_0__1__FORWARD__DATA__6_, 
        east_in_0__1__FORWARD__DATA__5_, east_in_0__1__FORWARD__DATA__4_, 
        east_in_0__1__FORWARD__DATA__3_, east_in_0__1__FORWARD__DATA__2_, 
        east_in_0__1__FORWARD__DATA__1_, east_in_0__1__FORWARD__DATA__0_}), 
        .east_in_b(east_in_0__1__BACKWARD__ACK), .south_in_f({
        north_out_req1[0], north_out_1__1__FORWARD__DATA__34_, 
        north_out_1__1__FORWARD__DATA__33_, north_out_1__1__FORWARD__DATA__32_, 
        north_out_1__1__FORWARD__DATA__31_, north_out_1__1__FORWARD__DATA__30_, 
        north_out_1__1__FORWARD__DATA__29_, north_out_1__1__FORWARD__DATA__28_, 
        north_out_1__1__FORWARD__DATA__27_, north_out_1__1__FORWARD__DATA__26_, 
        north_out_1__1__FORWARD__DATA__25_, north_out_1__1__FORWARD__DATA__24_, 
        north_out_1__1__FORWARD__DATA__23_, north_out_1__1__FORWARD__DATA__22_, 
        north_out_1__1__FORWARD__DATA__21_, north_out_1__1__FORWARD__DATA__20_, 
        north_out_1__1__FORWARD__DATA__19_, north_out_1__1__FORWARD__DATA__18_, 
        north_out_1__1__FORWARD__DATA__17_, north_out_1__1__FORWARD__DATA__16_, 
        north_out_1__1__FORWARD__DATA__15_, north_out_1__1__FORWARD__DATA__14_, 
        north_out_1__1__FORWARD__DATA__13_, north_out_1__1__FORWARD__DATA__12_, 
        north_out_1__1__FORWARD__DATA__11_, north_out_1__1__FORWARD__DATA__10_, 
        north_out_1__1__FORWARD__DATA__9_, north_out_1__1__FORWARD__DATA__8_, 
        north_out_1__1__FORWARD__DATA__7_, north_out_1__1__FORWARD__DATA__6_, 
        north_out_1__1__FORWARD__DATA__5_, north_out_1__1__FORWARD__DATA__4_, 
        north_out_1__1__FORWARD__DATA__3_, north_out_1__1__FORWARD__DATA__2_, 
        north_out_1__1__FORWARD__DATA__1_, north_out_1__1__FORWARD__DATA__0_}), 
        .south_in_b(south_in_0__1__BACKWARD__ACK), .west_in_f({
        east_out_req1[3], east_out_0__0__FORWARD__DATA__34_, 
        east_out_0__0__FORWARD__DATA__33_, east_out_0__0__FORWARD__DATA__32_, 
        east_out_0__0__FORWARD__DATA__31_, east_out_0__0__FORWARD__DATA__30_, 
        east_out_0__0__FORWARD__DATA__29_, east_out_0__0__FORWARD__DATA__28_, 
        east_out_0__0__FORWARD__DATA__27_, east_out_0__0__FORWARD__DATA__26_, 
        east_out_0__0__FORWARD__DATA__25_, east_out_0__0__FORWARD__DATA__24_, 
        east_out_0__0__FORWARD__DATA__23_, east_out_0__0__FORWARD__DATA__22_, 
        east_out_0__0__FORWARD__DATA__21_, east_out_0__0__FORWARD__DATA__20_, 
        east_out_0__0__FORWARD__DATA__19_, east_out_0__0__FORWARD__DATA__18_, 
        east_out_0__0__FORWARD__DATA__17_, east_out_0__0__FORWARD__DATA__16_, 
        east_out_0__0__FORWARD__DATA__15_, east_out_0__0__FORWARD__DATA__14_, 
        east_out_0__0__FORWARD__DATA__13_, east_out_0__0__FORWARD__DATA__12_, 
        east_out_0__0__FORWARD__DATA__11_, east_out_0__0__FORWARD__DATA__10_, 
        east_out_0__0__FORWARD__DATA__9_, east_out_0__0__FORWARD__DATA__8_, 
        east_out_0__0__FORWARD__DATA__7_, east_out_0__0__FORWARD__DATA__6_, 
        east_out_0__0__FORWARD__DATA__5_, east_out_0__0__FORWARD__DATA__4_, 
        east_out_0__0__FORWARD__DATA__3_, east_out_0__0__FORWARD__DATA__2_, 
        east_out_0__0__FORWARD__DATA__1_, east_out_0__0__FORWARD__DATA__0_}), 
        .west_in_b(west_in_0__1__BACKWARD__ACK), .north_out_f({
        north_out_0__1__FORWARD__REQ_, north_out_0__1__FORWARD__DATA__34_, 
        north_out_0__1__FORWARD__DATA__33_, north_out_0__1__FORWARD__DATA__32_, 
        north_out_0__1__FORWARD__DATA__31_, north_out_0__1__FORWARD__DATA__30_, 
        north_out_0__1__FORWARD__DATA__29_, north_out_0__1__FORWARD__DATA__28_, 
        north_out_0__1__FORWARD__DATA__27_, north_out_0__1__FORWARD__DATA__26_, 
        north_out_0__1__FORWARD__DATA__25_, north_out_0__1__FORWARD__DATA__24_, 
        north_out_0__1__FORWARD__DATA__23_, north_out_0__1__FORWARD__DATA__22_, 
        north_out_0__1__FORWARD__DATA__21_, north_out_0__1__FORWARD__DATA__20_, 
        north_out_0__1__FORWARD__DATA__19_, north_out_0__1__FORWARD__DATA__18_, 
        north_out_0__1__FORWARD__DATA__17_, north_out_0__1__FORWARD__DATA__16_, 
        north_out_0__1__FORWARD__DATA__15_, north_out_0__1__FORWARD__DATA__14_, 
        north_out_0__1__FORWARD__DATA__13_, north_out_0__1__FORWARD__DATA__12_, 
        north_out_0__1__FORWARD__DATA__11_, north_out_0__1__FORWARD__DATA__10_, 
        north_out_0__1__FORWARD__DATA__9_, north_out_0__1__FORWARD__DATA__8_, 
        north_out_0__1__FORWARD__DATA__7_, north_out_0__1__FORWARD__DATA__6_, 
        north_out_0__1__FORWARD__DATA__5_, north_out_0__1__FORWARD__DATA__4_, 
        north_out_0__1__FORWARD__DATA__3_, north_out_0__1__FORWARD__DATA__2_, 
        north_out_0__1__FORWARD__DATA__1_, north_out_0__1__FORWARD__DATA__0_}), 
        .north_out_b(south_in_ack1[0]), .east_out_f({
        east_out_0__1__FORWARD__REQ_, west_in_0__0__FORWARD__DATA__34_, 
        west_in_0__0__FORWARD__DATA__33_, west_in_0__0__FORWARD__DATA__32_, 
        west_in_0__0__FORWARD__DATA__31_, west_in_0__0__FORWARD__DATA__30_, 
        west_in_0__0__FORWARD__DATA__29_, west_in_0__0__FORWARD__DATA__28_, 
        west_in_0__0__FORWARD__DATA__27_, west_in_0__0__FORWARD__DATA__26_, 
        west_in_0__0__FORWARD__DATA__25_, west_in_0__0__FORWARD__DATA__24_, 
        west_in_0__0__FORWARD__DATA__23_, west_in_0__0__FORWARD__DATA__22_, 
        west_in_0__0__FORWARD__DATA__21_, west_in_0__0__FORWARD__DATA__20_, 
        west_in_0__0__FORWARD__DATA__19_, west_in_0__0__FORWARD__DATA__18_, 
        west_in_0__0__FORWARD__DATA__17_, west_in_0__0__FORWARD__DATA__16_, 
        west_in_0__0__FORWARD__DATA__15_, west_in_0__0__FORWARD__DATA__14_, 
        west_in_0__0__FORWARD__DATA__13_, west_in_0__0__FORWARD__DATA__12_, 
        west_in_0__0__FORWARD__DATA__11_, west_in_0__0__FORWARD__DATA__10_, 
        west_in_0__0__FORWARD__DATA__9_, west_in_0__0__FORWARD__DATA__8_, 
        west_in_0__0__FORWARD__DATA__7_, west_in_0__0__FORWARD__DATA__6_, 
        west_in_0__0__FORWARD__DATA__5_, west_in_0__0__FORWARD__DATA__4_, 
        west_in_0__0__FORWARD__DATA__3_, west_in_0__0__FORWARD__DATA__2_, 
        west_in_0__0__FORWARD__DATA__1_, west_in_0__0__FORWARD__DATA__0_}), 
        .east_out_b(west_in_ack1[3]), .south_out_f({
        south_out_0__1__FORWARD__REQ_, south_out_0__1__FORWARD__DATA__34_, 
        south_out_0__1__FORWARD__DATA__33_, south_out_0__1__FORWARD__DATA__32_, 
        south_out_0__1__FORWARD__DATA__31_, south_out_0__1__FORWARD__DATA__30_, 
        south_out_0__1__FORWARD__DATA__29_, south_out_0__1__FORWARD__DATA__28_, 
        south_out_0__1__FORWARD__DATA__27_, south_out_0__1__FORWARD__DATA__26_, 
        south_out_0__1__FORWARD__DATA__25_, south_out_0__1__FORWARD__DATA__24_, 
        south_out_0__1__FORWARD__DATA__23_, south_out_0__1__FORWARD__DATA__22_, 
        south_out_0__1__FORWARD__DATA__21_, south_out_0__1__FORWARD__DATA__20_, 
        south_out_0__1__FORWARD__DATA__19_, south_out_0__1__FORWARD__DATA__18_, 
        south_out_0__1__FORWARD__DATA__17_, south_out_0__1__FORWARD__DATA__16_, 
        south_out_0__1__FORWARD__DATA__15_, south_out_0__1__FORWARD__DATA__14_, 
        south_out_0__1__FORWARD__DATA__13_, south_out_0__1__FORWARD__DATA__12_, 
        south_out_0__1__FORWARD__DATA__11_, south_out_0__1__FORWARD__DATA__10_, 
        south_out_0__1__FORWARD__DATA__9_, south_out_0__1__FORWARD__DATA__8_, 
        south_out_0__1__FORWARD__DATA__7_, south_out_0__1__FORWARD__DATA__6_, 
        south_out_0__1__FORWARD__DATA__5_, south_out_0__1__FORWARD__DATA__4_, 
        south_out_0__1__FORWARD__DATA__3_, south_out_0__1__FORWARD__DATA__2_, 
        south_out_0__1__FORWARD__DATA__1_, south_out_0__1__FORWARD__DATA__0_}), 
        .south_out_b(north_in_ack1[0]), .west_out_f({
        west_out_0__1__FORWARD__REQ_, west_out_0__1__FORWARD__DATA__34_, 
        west_out_0__1__FORWARD__DATA__33_, west_out_0__1__FORWARD__DATA__32_, 
        west_out_0__1__FORWARD__DATA__31_, west_out_0__1__FORWARD__DATA__30_, 
        west_out_0__1__FORWARD__DATA__29_, west_out_0__1__FORWARD__DATA__28_, 
        west_out_0__1__FORWARD__DATA__27_, west_out_0__1__FORWARD__DATA__26_, 
        west_out_0__1__FORWARD__DATA__25_, west_out_0__1__FORWARD__DATA__24_, 
        west_out_0__1__FORWARD__DATA__23_, west_out_0__1__FORWARD__DATA__22_, 
        west_out_0__1__FORWARD__DATA__21_, west_out_0__1__FORWARD__DATA__20_, 
        west_out_0__1__FORWARD__DATA__19_, west_out_0__1__FORWARD__DATA__18_, 
        west_out_0__1__FORWARD__DATA__17_, west_out_0__1__FORWARD__DATA__16_, 
        west_out_0__1__FORWARD__DATA__15_, west_out_0__1__FORWARD__DATA__14_, 
        west_out_0__1__FORWARD__DATA__13_, west_out_0__1__FORWARD__DATA__12_, 
        west_out_0__1__FORWARD__DATA__11_, west_out_0__1__FORWARD__DATA__10_, 
        west_out_0__1__FORWARD__DATA__9_, west_out_0__1__FORWARD__DATA__8_, 
        west_out_0__1__FORWARD__DATA__7_, west_out_0__1__FORWARD__DATA__6_, 
        west_out_0__1__FORWARD__DATA__5_, west_out_0__1__FORWARD__DATA__4_, 
        west_out_0__1__FORWARD__DATA__3_, west_out_0__1__FORWARD__DATA__2_, 
        west_out_0__1__FORWARD__DATA__1_, west_out_0__1__FORWARD__DATA__0_}), 
        .west_out_b(east_in_ack1[3]) );
  noc_node_1 node_0_0 ( .p_clk(p_clk), .n_clk(n_clk), .reset(reset), .proc_in(
        p_ports_in[65:0]), .proc_out(p_ports_out[33:0]), .spm_in(
        spm_ports_in[65:0]), .spm_out({spm_ports_out[97:96], 
        spm_ports_out_0__0__MADDR__31_, spm_ports_out_0__0__MADDR__30_, 
        spm_ports_out_0__0__MADDR__29_, spm_ports_out_0__0__MADDR__28_, 
        spm_ports_out_0__0__MADDR__27_, spm_ports_out_0__0__MADDR__26_, 
        spm_ports_out_0__0__MADDR__25_, spm_ports_out_0__0__MADDR__24_, 
        spm_ports_out_0__0__MADDR__23_, spm_ports_out_0__0__MADDR__22_, 
        spm_ports_out_0__0__MADDR__21_, spm_ports_out_0__0__MADDR__20_, 
        spm_ports_out_0__0__MADDR__19_, spm_ports_out_0__0__MADDR__18_, 
        spm_ports_out_0__0__MADDR__17_, spm_ports_out_0__0__MADDR__16_, 
        spm_ports_out_0__0__MADDR__15_, spm_ports_out[78:0]}), .north_in_f({
        south_out_req1[1], north_in_0__0__FORWARD__DATA__34_, 
        north_in_0__0__FORWARD__DATA__33_, north_in_0__0__FORWARD__DATA__32_, 
        north_in_0__0__FORWARD__DATA__31_, north_in_0__0__FORWARD__DATA__30_, 
        north_in_0__0__FORWARD__DATA__29_, north_in_0__0__FORWARD__DATA__28_, 
        north_in_0__0__FORWARD__DATA__27_, north_in_0__0__FORWARD__DATA__26_, 
        north_in_0__0__FORWARD__DATA__25_, north_in_0__0__FORWARD__DATA__24_, 
        north_in_0__0__FORWARD__DATA__23_, north_in_0__0__FORWARD__DATA__22_, 
        north_in_0__0__FORWARD__DATA__21_, north_in_0__0__FORWARD__DATA__20_, 
        north_in_0__0__FORWARD__DATA__19_, north_in_0__0__FORWARD__DATA__18_, 
        north_in_0__0__FORWARD__DATA__17_, north_in_0__0__FORWARD__DATA__16_, 
        north_in_0__0__FORWARD__DATA__15_, north_in_0__0__FORWARD__DATA__14_, 
        north_in_0__0__FORWARD__DATA__13_, north_in_0__0__FORWARD__DATA__12_, 
        north_in_0__0__FORWARD__DATA__11_, north_in_0__0__FORWARD__DATA__10_, 
        north_in_0__0__FORWARD__DATA__9_, north_in_0__0__FORWARD__DATA__8_, 
        north_in_0__0__FORWARD__DATA__7_, north_in_0__0__FORWARD__DATA__6_, 
        north_in_0__0__FORWARD__DATA__5_, north_in_0__0__FORWARD__DATA__4_, 
        north_in_0__0__FORWARD__DATA__3_, north_in_0__0__FORWARD__DATA__2_, 
        north_in_0__0__FORWARD__DATA__1_, north_in_0__0__FORWARD__DATA__0_}), 
        .north_in_b(north_in_0__0__BACKWARD__ACK), .east_in_f({
        west_out_req1[2], west_out_0__1__FORWARD__DATA__34_, 
        west_out_0__1__FORWARD__DATA__33_, west_out_0__1__FORWARD__DATA__32_, 
        west_out_0__1__FORWARD__DATA__31_, west_out_0__1__FORWARD__DATA__30_, 
        west_out_0__1__FORWARD__DATA__29_, west_out_0__1__FORWARD__DATA__28_, 
        west_out_0__1__FORWARD__DATA__27_, west_out_0__1__FORWARD__DATA__26_, 
        west_out_0__1__FORWARD__DATA__25_, west_out_0__1__FORWARD__DATA__24_, 
        west_out_0__1__FORWARD__DATA__23_, west_out_0__1__FORWARD__DATA__22_, 
        west_out_0__1__FORWARD__DATA__21_, west_out_0__1__FORWARD__DATA__20_, 
        west_out_0__1__FORWARD__DATA__19_, west_out_0__1__FORWARD__DATA__18_, 
        west_out_0__1__FORWARD__DATA__17_, west_out_0__1__FORWARD__DATA__16_, 
        west_out_0__1__FORWARD__DATA__15_, west_out_0__1__FORWARD__DATA__14_, 
        west_out_0__1__FORWARD__DATA__13_, west_out_0__1__FORWARD__DATA__12_, 
        west_out_0__1__FORWARD__DATA__11_, west_out_0__1__FORWARD__DATA__10_, 
        west_out_0__1__FORWARD__DATA__9_, west_out_0__1__FORWARD__DATA__8_, 
        west_out_0__1__FORWARD__DATA__7_, west_out_0__1__FORWARD__DATA__6_, 
        west_out_0__1__FORWARD__DATA__5_, west_out_0__1__FORWARD__DATA__4_, 
        west_out_0__1__FORWARD__DATA__3_, west_out_0__1__FORWARD__DATA__2_, 
        west_out_0__1__FORWARD__DATA__1_, west_out_0__1__FORWARD__DATA__0_}), 
        .east_in_b(east_in_0__0__BACKWARD__ACK), .south_in_f({
        north_out_req1[1], north_out_1__0__FORWARD__DATA__34_, 
        north_out_1__0__FORWARD__DATA__33_, north_out_1__0__FORWARD__DATA__32_, 
        north_out_1__0__FORWARD__DATA__31_, north_out_1__0__FORWARD__DATA__30_, 
        north_out_1__0__FORWARD__DATA__29_, north_out_1__0__FORWARD__DATA__28_, 
        north_out_1__0__FORWARD__DATA__27_, north_out_1__0__FORWARD__DATA__26_, 
        north_out_1__0__FORWARD__DATA__25_, north_out_1__0__FORWARD__DATA__24_, 
        north_out_1__0__FORWARD__DATA__23_, north_out_1__0__FORWARD__DATA__22_, 
        north_out_1__0__FORWARD__DATA__21_, north_out_1__0__FORWARD__DATA__20_, 
        north_out_1__0__FORWARD__DATA__19_, north_out_1__0__FORWARD__DATA__18_, 
        north_out_1__0__FORWARD__DATA__17_, north_out_1__0__FORWARD__DATA__16_, 
        north_out_1__0__FORWARD__DATA__15_, north_out_1__0__FORWARD__DATA__14_, 
        north_out_1__0__FORWARD__DATA__13_, north_out_1__0__FORWARD__DATA__12_, 
        north_out_1__0__FORWARD__DATA__11_, north_out_1__0__FORWARD__DATA__10_, 
        north_out_1__0__FORWARD__DATA__9_, north_out_1__0__FORWARD__DATA__8_, 
        north_out_1__0__FORWARD__DATA__7_, north_out_1__0__FORWARD__DATA__6_, 
        north_out_1__0__FORWARD__DATA__5_, north_out_1__0__FORWARD__DATA__4_, 
        north_out_1__0__FORWARD__DATA__3_, north_out_1__0__FORWARD__DATA__2_, 
        north_out_1__0__FORWARD__DATA__1_, north_out_1__0__FORWARD__DATA__0_}), 
        .south_in_b(south_in_0__0__BACKWARD__ACK), .west_in_f({
        east_out_req1[2], west_in_0__0__FORWARD__DATA__34_, 
        west_in_0__0__FORWARD__DATA__33_, west_in_0__0__FORWARD__DATA__32_, 
        west_in_0__0__FORWARD__DATA__31_, west_in_0__0__FORWARD__DATA__30_, 
        west_in_0__0__FORWARD__DATA__29_, west_in_0__0__FORWARD__DATA__28_, 
        west_in_0__0__FORWARD__DATA__27_, west_in_0__0__FORWARD__DATA__26_, 
        west_in_0__0__FORWARD__DATA__25_, west_in_0__0__FORWARD__DATA__24_, 
        west_in_0__0__FORWARD__DATA__23_, west_in_0__0__FORWARD__DATA__22_, 
        west_in_0__0__FORWARD__DATA__21_, west_in_0__0__FORWARD__DATA__20_, 
        west_in_0__0__FORWARD__DATA__19_, west_in_0__0__FORWARD__DATA__18_, 
        west_in_0__0__FORWARD__DATA__17_, west_in_0__0__FORWARD__DATA__16_, 
        west_in_0__0__FORWARD__DATA__15_, west_in_0__0__FORWARD__DATA__14_, 
        west_in_0__0__FORWARD__DATA__13_, west_in_0__0__FORWARD__DATA__12_, 
        west_in_0__0__FORWARD__DATA__11_, west_in_0__0__FORWARD__DATA__10_, 
        west_in_0__0__FORWARD__DATA__9_, west_in_0__0__FORWARD__DATA__8_, 
        west_in_0__0__FORWARD__DATA__7_, west_in_0__0__FORWARD__DATA__6_, 
        west_in_0__0__FORWARD__DATA__5_, west_in_0__0__FORWARD__DATA__4_, 
        west_in_0__0__FORWARD__DATA__3_, west_in_0__0__FORWARD__DATA__2_, 
        west_in_0__0__FORWARD__DATA__1_, west_in_0__0__FORWARD__DATA__0_}), 
        .west_in_b(west_in_0__0__BACKWARD__ACK), .north_out_f({
        north_out_0__0__FORWARD__REQ_, south_in_1__0__FORWARD__DATA__34_, 
        south_in_1__0__FORWARD__DATA__33_, south_in_1__0__FORWARD__DATA__32_, 
        south_in_1__0__FORWARD__DATA__31_, south_in_1__0__FORWARD__DATA__30_, 
        south_in_1__0__FORWARD__DATA__29_, south_in_1__0__FORWARD__DATA__28_, 
        south_in_1__0__FORWARD__DATA__27_, south_in_1__0__FORWARD__DATA__26_, 
        south_in_1__0__FORWARD__DATA__25_, south_in_1__0__FORWARD__DATA__24_, 
        south_in_1__0__FORWARD__DATA__23_, south_in_1__0__FORWARD__DATA__22_, 
        south_in_1__0__FORWARD__DATA__21_, south_in_1__0__FORWARD__DATA__20_, 
        south_in_1__0__FORWARD__DATA__19_, south_in_1__0__FORWARD__DATA__18_, 
        south_in_1__0__FORWARD__DATA__17_, south_in_1__0__FORWARD__DATA__16_, 
        south_in_1__0__FORWARD__DATA__15_, south_in_1__0__FORWARD__DATA__14_, 
        south_in_1__0__FORWARD__DATA__13_, south_in_1__0__FORWARD__DATA__12_, 
        south_in_1__0__FORWARD__DATA__11_, south_in_1__0__FORWARD__DATA__10_, 
        south_in_1__0__FORWARD__DATA__9_, south_in_1__0__FORWARD__DATA__8_, 
        south_in_1__0__FORWARD__DATA__7_, south_in_1__0__FORWARD__DATA__6_, 
        south_in_1__0__FORWARD__DATA__5_, south_in_1__0__FORWARD__DATA__4_, 
        south_in_1__0__FORWARD__DATA__3_, south_in_1__0__FORWARD__DATA__2_, 
        south_in_1__0__FORWARD__DATA__1_, south_in_1__0__FORWARD__DATA__0_}), 
        .north_out_b(south_in_ack1[1]), .east_out_f({
        east_out_0__0__FORWARD__REQ_, east_out_0__0__FORWARD__DATA__34_, 
        east_out_0__0__FORWARD__DATA__33_, east_out_0__0__FORWARD__DATA__32_, 
        east_out_0__0__FORWARD__DATA__31_, east_out_0__0__FORWARD__DATA__30_, 
        east_out_0__0__FORWARD__DATA__29_, east_out_0__0__FORWARD__DATA__28_, 
        east_out_0__0__FORWARD__DATA__27_, east_out_0__0__FORWARD__DATA__26_, 
        east_out_0__0__FORWARD__DATA__25_, east_out_0__0__FORWARD__DATA__24_, 
        east_out_0__0__FORWARD__DATA__23_, east_out_0__0__FORWARD__DATA__22_, 
        east_out_0__0__FORWARD__DATA__21_, east_out_0__0__FORWARD__DATA__20_, 
        east_out_0__0__FORWARD__DATA__19_, east_out_0__0__FORWARD__DATA__18_, 
        east_out_0__0__FORWARD__DATA__17_, east_out_0__0__FORWARD__DATA__16_, 
        east_out_0__0__FORWARD__DATA__15_, east_out_0__0__FORWARD__DATA__14_, 
        east_out_0__0__FORWARD__DATA__13_, east_out_0__0__FORWARD__DATA__12_, 
        east_out_0__0__FORWARD__DATA__11_, east_out_0__0__FORWARD__DATA__10_, 
        east_out_0__0__FORWARD__DATA__9_, east_out_0__0__FORWARD__DATA__8_, 
        east_out_0__0__FORWARD__DATA__7_, east_out_0__0__FORWARD__DATA__6_, 
        east_out_0__0__FORWARD__DATA__5_, east_out_0__0__FORWARD__DATA__4_, 
        east_out_0__0__FORWARD__DATA__3_, east_out_0__0__FORWARD__DATA__2_, 
        east_out_0__0__FORWARD__DATA__1_, east_out_0__0__FORWARD__DATA__0_}), 
        .east_out_b(west_in_ack1[2]), .south_out_f({
        south_out_0__0__FORWARD__REQ_, south_out_0__0__FORWARD__DATA__34_, 
        south_out_0__0__FORWARD__DATA__33_, south_out_0__0__FORWARD__DATA__32_, 
        south_out_0__0__FORWARD__DATA__31_, south_out_0__0__FORWARD__DATA__30_, 
        south_out_0__0__FORWARD__DATA__29_, south_out_0__0__FORWARD__DATA__28_, 
        south_out_0__0__FORWARD__DATA__27_, south_out_0__0__FORWARD__DATA__26_, 
        south_out_0__0__FORWARD__DATA__25_, south_out_0__0__FORWARD__DATA__24_, 
        south_out_0__0__FORWARD__DATA__23_, south_out_0__0__FORWARD__DATA__22_, 
        south_out_0__0__FORWARD__DATA__21_, south_out_0__0__FORWARD__DATA__20_, 
        south_out_0__0__FORWARD__DATA__19_, south_out_0__0__FORWARD__DATA__18_, 
        south_out_0__0__FORWARD__DATA__17_, south_out_0__0__FORWARD__DATA__16_, 
        south_out_0__0__FORWARD__DATA__15_, south_out_0__0__FORWARD__DATA__14_, 
        south_out_0__0__FORWARD__DATA__13_, south_out_0__0__FORWARD__DATA__12_, 
        south_out_0__0__FORWARD__DATA__11_, south_out_0__0__FORWARD__DATA__10_, 
        south_out_0__0__FORWARD__DATA__9_, south_out_0__0__FORWARD__DATA__8_, 
        south_out_0__0__FORWARD__DATA__7_, south_out_0__0__FORWARD__DATA__6_, 
        south_out_0__0__FORWARD__DATA__5_, south_out_0__0__FORWARD__DATA__4_, 
        south_out_0__0__FORWARD__DATA__3_, south_out_0__0__FORWARD__DATA__2_, 
        south_out_0__0__FORWARD__DATA__1_, south_out_0__0__FORWARD__DATA__0_}), 
        .south_out_b(north_in_ack1[1]), .west_out_f({
        west_out_0__0__FORWARD__REQ_, east_in_0__1__FORWARD__DATA__34_, 
        east_in_0__1__FORWARD__DATA__33_, east_in_0__1__FORWARD__DATA__32_, 
        east_in_0__1__FORWARD__DATA__31_, east_in_0__1__FORWARD__DATA__30_, 
        east_in_0__1__FORWARD__DATA__29_, east_in_0__1__FORWARD__DATA__28_, 
        east_in_0__1__FORWARD__DATA__27_, east_in_0__1__FORWARD__DATA__26_, 
        east_in_0__1__FORWARD__DATA__25_, east_in_0__1__FORWARD__DATA__24_, 
        east_in_0__1__FORWARD__DATA__23_, east_in_0__1__FORWARD__DATA__22_, 
        east_in_0__1__FORWARD__DATA__21_, east_in_0__1__FORWARD__DATA__20_, 
        east_in_0__1__FORWARD__DATA__19_, east_in_0__1__FORWARD__DATA__18_, 
        east_in_0__1__FORWARD__DATA__17_, east_in_0__1__FORWARD__DATA__16_, 
        east_in_0__1__FORWARD__DATA__15_, east_in_0__1__FORWARD__DATA__14_, 
        east_in_0__1__FORWARD__DATA__13_, east_in_0__1__FORWARD__DATA__12_, 
        east_in_0__1__FORWARD__DATA__11_, east_in_0__1__FORWARD__DATA__10_, 
        east_in_0__1__FORWARD__DATA__9_, east_in_0__1__FORWARD__DATA__8_, 
        east_in_0__1__FORWARD__DATA__7_, east_in_0__1__FORWARD__DATA__6_, 
        east_in_0__1__FORWARD__DATA__5_, east_in_0__1__FORWARD__DATA__4_, 
        east_in_0__1__FORWARD__DATA__3_, east_in_0__1__FORWARD__DATA__2_, 
        east_in_0__1__FORWARD__DATA__1_, east_in_0__1__FORWARD__DATA__0_}), 
        .west_out_b(east_in_ack1[2]) );
  HS65_LS_IVX9 I_29 ( .A(n161), .Z(south_in_ack1[1]) );
  HS65_LS_IVX9 I_47 ( .A(n169), .Z(west_in_ack1[2]) );
  HS65_LS_IVX9 I_25 ( .A(n177), .Z(north_in_ack1[1]) );
  HS65_LS_IVX9 I_43 ( .A(n57), .Z(east_in_ack1[2]) );
  HS65_LS_IVX9 I_13 ( .A(n65), .Z(south_in_ack1[0]) );
  HS65_LS_IVX9 I_63 ( .A(n73), .Z(west_in_ack1[3]) );
  HS65_LS_IVX9 I_9 ( .A(n81), .Z(north_in_ack1[0]) );
  HS65_LS_IVX9 I_59 ( .A(n89), .Z(east_in_ack1[3]) );
  HS65_LS_IVX9 I_61 ( .A(n217), .Z(south_in_ack1[3]) );
  HS65_LS_IVX9 I_15 ( .A(n225), .Z(west_in_ack1[0]) );
  HS65_LS_IVX9 I_57 ( .A(n233), .Z(north_in_ack1[3]) );
  HS65_LS_IVX9 I_11 ( .A(n241), .Z(east_in_ack1[0]) );
  HS65_LS_IVX9 I_45 ( .A(n249), .Z(south_in_ack1[2]) );
  HS65_LS_IVX9 I_31 ( .A(n185), .Z(west_in_ack1[1]) );
  HS65_LS_IVX9 I_41 ( .A(n193), .Z(north_in_ack1[2]) );
  HS65_LS_IVX9 I_27 ( .A(n201), .Z(east_in_ack1[1]) );
  HS65_LS_IVX9 I_37 ( .A(n209), .Z(south_out_req1[2]) );
  HS65_LS_IVX9 I_35 ( .A(n97), .Z(east_out_req1[2]) );
  HS65_LS_IVX9 I_39 ( .A(n105), .Z(west_out_req1[2]) );
  HS65_LS_IVX9 I_17 ( .A(n113), .Z(north_out_req1[1]) );
  HS65_LS_IVX9 I_21 ( .A(n121), .Z(south_out_req1[1]) );
  HS65_LS_IVX9 I_51 ( .A(n129), .Z(east_out_req1[3]) );
  HS65_LS_IVX9 I_55 ( .A(n137), .Z(west_out_req1[3]) );
  HS65_LS_IVX9 I_1 ( .A(n145), .Z(north_out_req1[0]) );
  HS65_LS_IVX9 I_5 ( .A(n153), .Z(south_out_req1[0]) );
  HS65_LS_IVX9 I_3 ( .A(n1), .Z(east_out_req1[0]) );
  HS65_LS_IVX9 I_7 ( .A(n9), .Z(west_out_req1[0]) );
  HS65_LS_IVX9 I_49 ( .A(n17), .Z(north_out_req1[3]) );
  HS65_LS_IVX9 I_53 ( .A(n25), .Z(south_out_req1[3]) );
  HS65_LS_IVX9 I_19 ( .A(n33), .Z(east_out_req1[1]) );
  HS65_LS_IVX9 I_23 ( .A(n41), .Z(west_out_req1[1]) );
  HS65_LS_IVX9 I_33 ( .A(n49), .Z(north_out_req1[2]) );
  HS65_LH_IVX2 I_44 ( .A(south_in_0__1__BACKWARD__ACK), .Z(south_in_ack0[2])
         );
  HS65_LH_IVX2 I_10 ( .A(east_in_1__1__BACKWARD__ACK), .Z(east_in_ack0[0]) );
  HS65_LH_IVX2 I_56 ( .A(north_in_0__0__BACKWARD__ACK), .Z(north_in_ack0[3])
         );
  HS65_LH_IVX2 I_14 ( .A(west_in_1__1__BACKWARD__ACK), .Z(west_in_ack0[0]) );
  HS65_LH_IVX2 I_60 ( .A(south_in_0__0__BACKWARD__ACK), .Z(south_in_ack0[3])
         );
  HS65_LH_IVX2 I_36 ( .A(south_out_0__1__FORWARD__REQ_), .Z(south_out_req0[2])
         );
  HS65_LH_IVX2 I_26 ( .A(east_in_1__0__BACKWARD__ACK), .Z(east_in_ack0[1]) );
  HS65_LH_IVX2 I_40 ( .A(north_in_0__1__BACKWARD__ACK), .Z(north_in_ack0[2])
         );
  HS65_LH_IVX2 I_30 ( .A(west_in_1__0__BACKWARD__ACK), .Z(west_in_ack0[1]) );
  HS65_LH_IVX2 I_24 ( .A(north_in_1__0__BACKWARD__ACK), .Z(north_in_ack0[1])
         );
  HS65_LH_IVX2 I_46 ( .A(west_in_0__1__BACKWARD__ACK), .Z(west_in_ack0[2]) );
  HS65_LH_IVX2 I_28 ( .A(south_in_1__0__BACKWARD__ACK), .Z(south_in_ack0[1])
         );
  HS65_LH_IVX2 I_4 ( .A(south_out_1__1__FORWARD__REQ_), .Z(south_out_req0[0])
         );
  HS65_LH_IVX2 I_0 ( .A(north_out_1__1__FORWARD__REQ_), .Z(north_out_req0[0])
         );
  HS65_LH_IVX2 I_54 ( .A(west_out_0__0__FORWARD__REQ_), .Z(west_out_req0[3])
         );
  HS65_LH_IVX2 I_50 ( .A(east_out_0__0__FORWARD__REQ_), .Z(east_out_req0[3])
         );
  HS65_LH_IVX2 I_20 ( .A(south_out_1__0__FORWARD__REQ_), .Z(south_out_req0[1])
         );
  HS65_LH_IVX2 I_16 ( .A(north_out_1__0__FORWARD__REQ_), .Z(north_out_req0[1])
         );
  HS65_LH_IVX2 I_38 ( .A(west_out_0__1__FORWARD__REQ_), .Z(west_out_req0[2])
         );
  HS65_LH_IVX2 I_34 ( .A(east_out_0__1__FORWARD__REQ_), .Z(east_out_req0[2])
         );
  HS65_LH_IVX2 I_58 ( .A(east_in_0__0__BACKWARD__ACK), .Z(east_in_ack0[3]) );
  HS65_LH_IVX2 I_8 ( .A(north_in_1__1__BACKWARD__ACK), .Z(north_in_ack0[0])
         );
  HS65_LH_IVX2 I_62 ( .A(west_in_0__0__BACKWARD__ACK), .Z(west_in_ack0[3]) );
  HS65_LH_IVX2 I_12 ( .A(south_in_1__1__BACKWARD__ACK), .Z(south_in_ack0[0])
         );
  HS65_LH_IVX2 I_42 ( .A(east_in_0__1__BACKWARD__ACK), .Z(east_in_ack0[2]) );
  HS65_LH_IVX2 I_32 ( .A(north_out_0__1__FORWARD__REQ_), .Z(north_out_req0[2])
         );
  HS65_LH_IVX2 I_22 ( .A(west_out_1__0__FORWARD__REQ_), .Z(west_out_req0[1])
         );
  HS65_LH_IVX2 I_18 ( .A(east_out_1__0__FORWARD__REQ_), .Z(east_out_req0[1])
         );
  HS65_LH_IVX2 I_52 ( .A(south_out_0__0__FORWARD__REQ_), .Z(south_out_req0[3])
         );
  HS65_LH_IVX2 I_48 ( .A(north_out_0__0__FORWARD__REQ_), .Z(north_out_req0[3])
         );
  HS65_LH_IVX2 I_6 ( .A(west_out_1__1__FORWARD__REQ_), .Z(west_out_req0[0]) );
  HS65_LH_IVX2 I_2 ( .A(east_out_1__1__FORWARD__REQ_), .Z(east_out_req0[0]) );
  HS65_LS_BFX9 U1 ( .A(n2), .Z(n1) );
  HS65_LS_BFX9 U2 ( .A(n3), .Z(n2) );
  HS65_LS_BFX9 U3 ( .A(n4), .Z(n3) );
  HS65_LS_BFX9 U4 ( .A(n5), .Z(n4) );
  HS65_LS_BFX9 U5 ( .A(n6), .Z(n5) );
  HS65_LS_BFX9 U6 ( .A(n7), .Z(n6) );
  HS65_LS_BFX9 U7 ( .A(n8), .Z(n7) );
  HS65_LS_BFX9 U8 ( .A(east_out_req0[0]), .Z(n8) );
  HS65_LS_BFX9 U9 ( .A(n10), .Z(n9) );
  HS65_LS_BFX9 U10 ( .A(n11), .Z(n10) );
  HS65_LS_BFX9 U11 ( .A(n12), .Z(n11) );
  HS65_LS_BFX9 U12 ( .A(n13), .Z(n12) );
  HS65_LS_BFX9 U13 ( .A(n14), .Z(n13) );
  HS65_LS_BFX9 U14 ( .A(n15), .Z(n14) );
  HS65_LS_BFX9 U15 ( .A(n16), .Z(n15) );
  HS65_LS_BFX9 U16 ( .A(west_out_req0[0]), .Z(n16) );
  HS65_LS_BFX9 U17 ( .A(n18), .Z(n17) );
  HS65_LS_BFX9 U18 ( .A(n19), .Z(n18) );
  HS65_LS_BFX9 U19 ( .A(n20), .Z(n19) );
  HS65_LS_BFX9 U20 ( .A(n21), .Z(n20) );
  HS65_LS_BFX9 U21 ( .A(n22), .Z(n21) );
  HS65_LS_BFX9 U22 ( .A(n23), .Z(n22) );
  HS65_LS_BFX9 U23 ( .A(n24), .Z(n23) );
  HS65_LS_BFX9 U24 ( .A(north_out_req0[3]), .Z(n24) );
  HS65_LS_BFX9 U25 ( .A(n26), .Z(n25) );
  HS65_LS_BFX9 U26 ( .A(n27), .Z(n26) );
  HS65_LS_BFX9 U27 ( .A(n28), .Z(n27) );
  HS65_LS_BFX9 U28 ( .A(n29), .Z(n28) );
  HS65_LS_BFX9 U29 ( .A(n30), .Z(n29) );
  HS65_LS_BFX9 U30 ( .A(n31), .Z(n30) );
  HS65_LS_BFX9 U31 ( .A(n32), .Z(n31) );
  HS65_LS_BFX9 U32 ( .A(south_out_req0[3]), .Z(n32) );
  HS65_LS_BFX9 U33 ( .A(n34), .Z(n33) );
  HS65_LS_BFX9 U34 ( .A(n35), .Z(n34) );
  HS65_LS_BFX9 U35 ( .A(n36), .Z(n35) );
  HS65_LS_BFX9 U36 ( .A(n37), .Z(n36) );
  HS65_LS_BFX9 U37 ( .A(n38), .Z(n37) );
  HS65_LS_BFX9 U38 ( .A(n39), .Z(n38) );
  HS65_LS_BFX9 U39 ( .A(n40), .Z(n39) );
  HS65_LS_BFX9 U40 ( .A(east_out_req0[1]), .Z(n40) );
  HS65_LS_BFX9 U41 ( .A(n42), .Z(n41) );
  HS65_LS_BFX9 U42 ( .A(n43), .Z(n42) );
  HS65_LS_BFX9 U43 ( .A(n44), .Z(n43) );
  HS65_LS_BFX9 U44 ( .A(n45), .Z(n44) );
  HS65_LS_BFX9 U45 ( .A(n46), .Z(n45) );
  HS65_LS_BFX9 U46 ( .A(n47), .Z(n46) );
  HS65_LS_BFX9 U47 ( .A(n48), .Z(n47) );
  HS65_LS_BFX9 U48 ( .A(west_out_req0[1]), .Z(n48) );
  HS65_LS_BFX9 U49 ( .A(n50), .Z(n49) );
  HS65_LS_BFX9 U50 ( .A(n51), .Z(n50) );
  HS65_LS_BFX9 U51 ( .A(n52), .Z(n51) );
  HS65_LS_BFX9 U52 ( .A(n53), .Z(n52) );
  HS65_LS_BFX9 U53 ( .A(n54), .Z(n53) );
  HS65_LS_BFX9 U54 ( .A(n55), .Z(n54) );
  HS65_LS_BFX9 U55 ( .A(n56), .Z(n55) );
  HS65_LS_BFX9 U56 ( .A(north_out_req0[2]), .Z(n56) );
  HS65_LS_BFX9 U57 ( .A(n58), .Z(n57) );
  HS65_LS_BFX9 U58 ( .A(n59), .Z(n58) );
  HS65_LS_BFX9 U59 ( .A(n60), .Z(n59) );
  HS65_LS_BFX9 U60 ( .A(n61), .Z(n60) );
  HS65_LS_BFX9 U61 ( .A(n62), .Z(n61) );
  HS65_LS_BFX9 U62 ( .A(n63), .Z(n62) );
  HS65_LS_BFX9 U63 ( .A(n64), .Z(n63) );
  HS65_LS_BFX9 U64 ( .A(east_in_ack0[2]), .Z(n64) );
  HS65_LS_BFX9 U65 ( .A(n66), .Z(n65) );
  HS65_LS_BFX9 U66 ( .A(n67), .Z(n66) );
  HS65_LS_BFX9 U67 ( .A(n68), .Z(n67) );
  HS65_LS_BFX9 U68 ( .A(n69), .Z(n68) );
  HS65_LS_BFX9 U69 ( .A(n70), .Z(n69) );
  HS65_LS_BFX9 U70 ( .A(n71), .Z(n70) );
  HS65_LS_BFX9 U71 ( .A(n72), .Z(n71) );
  HS65_LS_BFX9 U72 ( .A(south_in_ack0[0]), .Z(n72) );
  HS65_LS_BFX9 U73 ( .A(n74), .Z(n73) );
  HS65_LS_BFX9 U74 ( .A(n75), .Z(n74) );
  HS65_LS_BFX9 U75 ( .A(n76), .Z(n75) );
  HS65_LS_BFX9 U76 ( .A(n77), .Z(n76) );
  HS65_LS_BFX9 U77 ( .A(n78), .Z(n77) );
  HS65_LS_BFX9 U78 ( .A(n79), .Z(n78) );
  HS65_LS_BFX9 U79 ( .A(n80), .Z(n79) );
  HS65_LS_BFX9 U80 ( .A(west_in_ack0[3]), .Z(n80) );
  HS65_LS_BFX9 U81 ( .A(n82), .Z(n81) );
  HS65_LS_BFX9 U82 ( .A(n83), .Z(n82) );
  HS65_LS_BFX9 U83 ( .A(n84), .Z(n83) );
  HS65_LS_BFX9 U84 ( .A(n85), .Z(n84) );
  HS65_LS_BFX9 U85 ( .A(n86), .Z(n85) );
  HS65_LS_BFX9 U86 ( .A(n87), .Z(n86) );
  HS65_LS_BFX9 U87 ( .A(n88), .Z(n87) );
  HS65_LS_BFX9 U88 ( .A(north_in_ack0[0]), .Z(n88) );
  HS65_LS_BFX9 U89 ( .A(n90), .Z(n89) );
  HS65_LS_BFX9 U90 ( .A(n91), .Z(n90) );
  HS65_LS_BFX9 U91 ( .A(n92), .Z(n91) );
  HS65_LS_BFX9 U92 ( .A(n93), .Z(n92) );
  HS65_LS_BFX9 U93 ( .A(n94), .Z(n93) );
  HS65_LS_BFX9 U94 ( .A(n95), .Z(n94) );
  HS65_LS_BFX9 U95 ( .A(n96), .Z(n95) );
  HS65_LS_BFX9 U96 ( .A(east_in_ack0[3]), .Z(n96) );
  HS65_LS_BFX9 U97 ( .A(n98), .Z(n97) );
  HS65_LS_BFX9 U98 ( .A(n99), .Z(n98) );
  HS65_LS_BFX9 U99 ( .A(n100), .Z(n99) );
  HS65_LS_BFX9 U100 ( .A(n101), .Z(n100) );
  HS65_LS_BFX9 U101 ( .A(n102), .Z(n101) );
  HS65_LS_BFX9 U102 ( .A(n103), .Z(n102) );
  HS65_LS_BFX9 U103 ( .A(n104), .Z(n103) );
  HS65_LS_BFX9 U104 ( .A(east_out_req0[2]), .Z(n104) );
  HS65_LS_BFX9 U105 ( .A(n106), .Z(n105) );
  HS65_LS_BFX9 U106 ( .A(n107), .Z(n106) );
  HS65_LS_BFX9 U107 ( .A(n108), .Z(n107) );
  HS65_LS_BFX9 U108 ( .A(n109), .Z(n108) );
  HS65_LS_BFX9 U109 ( .A(n110), .Z(n109) );
  HS65_LS_BFX9 U110 ( .A(n111), .Z(n110) );
  HS65_LS_BFX9 U111 ( .A(n112), .Z(n111) );
  HS65_LS_BFX9 U112 ( .A(west_out_req0[2]), .Z(n112) );
  HS65_LS_BFX9 U113 ( .A(n114), .Z(n113) );
  HS65_LS_BFX9 U114 ( .A(n115), .Z(n114) );
  HS65_LS_BFX9 U115 ( .A(n116), .Z(n115) );
  HS65_LS_BFX9 U116 ( .A(n117), .Z(n116) );
  HS65_LS_BFX9 U117 ( .A(n118), .Z(n117) );
  HS65_LS_BFX9 U118 ( .A(n119), .Z(n118) );
  HS65_LS_BFX9 U119 ( .A(n120), .Z(n119) );
  HS65_LS_BFX9 U120 ( .A(north_out_req0[1]), .Z(n120) );
  HS65_LS_BFX9 U121 ( .A(n122), .Z(n121) );
  HS65_LS_BFX9 U122 ( .A(n123), .Z(n122) );
  HS65_LS_BFX9 U123 ( .A(n124), .Z(n123) );
  HS65_LS_BFX9 U124 ( .A(n125), .Z(n124) );
  HS65_LS_BFX9 U125 ( .A(n126), .Z(n125) );
  HS65_LS_BFX9 U126 ( .A(n127), .Z(n126) );
  HS65_LS_BFX9 U127 ( .A(n128), .Z(n127) );
  HS65_LS_BFX9 U128 ( .A(south_out_req0[1]), .Z(n128) );
  HS65_LS_BFX9 U129 ( .A(n130), .Z(n129) );
  HS65_LS_BFX9 U130 ( .A(n131), .Z(n130) );
  HS65_LS_BFX9 U131 ( .A(n132), .Z(n131) );
  HS65_LS_BFX9 U132 ( .A(n133), .Z(n132) );
  HS65_LS_BFX9 U133 ( .A(n134), .Z(n133) );
  HS65_LS_BFX9 U134 ( .A(n135), .Z(n134) );
  HS65_LS_BFX9 U135 ( .A(n136), .Z(n135) );
  HS65_LS_BFX9 U136 ( .A(east_out_req0[3]), .Z(n136) );
  HS65_LS_BFX9 U137 ( .A(n138), .Z(n137) );
  HS65_LS_BFX9 U138 ( .A(n139), .Z(n138) );
  HS65_LS_BFX9 U139 ( .A(n140), .Z(n139) );
  HS65_LS_BFX9 U140 ( .A(n141), .Z(n140) );
  HS65_LS_BFX9 U141 ( .A(n142), .Z(n141) );
  HS65_LS_BFX9 U142 ( .A(n143), .Z(n142) );
  HS65_LS_BFX9 U143 ( .A(n144), .Z(n143) );
  HS65_LS_BFX9 U144 ( .A(west_out_req0[3]), .Z(n144) );
  HS65_LS_BFX9 U145 ( .A(n146), .Z(n145) );
  HS65_LS_BFX9 U146 ( .A(n147), .Z(n146) );
  HS65_LS_BFX9 U147 ( .A(n148), .Z(n147) );
  HS65_LS_BFX9 U148 ( .A(n149), .Z(n148) );
  HS65_LS_BFX9 U149 ( .A(n150), .Z(n149) );
  HS65_LS_BFX9 U150 ( .A(n151), .Z(n150) );
  HS65_LS_BFX9 U151 ( .A(n152), .Z(n151) );
  HS65_LS_BFX9 U152 ( .A(north_out_req0[0]), .Z(n152) );
  HS65_LS_BFX9 U153 ( .A(n154), .Z(n153) );
  HS65_LS_BFX9 U154 ( .A(n155), .Z(n154) );
  HS65_LS_BFX9 U155 ( .A(n156), .Z(n155) );
  HS65_LS_BFX9 U156 ( .A(n157), .Z(n156) );
  HS65_LS_BFX9 U157 ( .A(n158), .Z(n157) );
  HS65_LS_BFX9 U158 ( .A(n159), .Z(n158) );
  HS65_LS_BFX9 U159 ( .A(n160), .Z(n159) );
  HS65_LS_BFX9 U160 ( .A(south_out_req0[0]), .Z(n160) );
  HS65_LS_BFX9 U161 ( .A(n162), .Z(n161) );
  HS65_LS_BFX9 U162 ( .A(n163), .Z(n162) );
  HS65_LS_BFX9 U163 ( .A(n164), .Z(n163) );
  HS65_LS_BFX9 U164 ( .A(n165), .Z(n164) );
  HS65_LS_BFX9 U165 ( .A(n166), .Z(n165) );
  HS65_LS_BFX9 U166 ( .A(n167), .Z(n166) );
  HS65_LS_BFX9 U167 ( .A(n168), .Z(n167) );
  HS65_LS_BFX9 U168 ( .A(south_in_ack0[1]), .Z(n168) );
  HS65_LS_BFX9 U169 ( .A(n170), .Z(n169) );
  HS65_LS_BFX9 U170 ( .A(n171), .Z(n170) );
  HS65_LS_BFX9 U171 ( .A(n172), .Z(n171) );
  HS65_LS_BFX9 U172 ( .A(n173), .Z(n172) );
  HS65_LS_BFX9 U173 ( .A(n174), .Z(n173) );
  HS65_LS_BFX9 U174 ( .A(n175), .Z(n174) );
  HS65_LS_BFX9 U175 ( .A(n176), .Z(n175) );
  HS65_LS_BFX9 U176 ( .A(west_in_ack0[2]), .Z(n176) );
  HS65_LS_BFX9 U177 ( .A(n178), .Z(n177) );
  HS65_LS_BFX9 U178 ( .A(n179), .Z(n178) );
  HS65_LS_BFX9 U179 ( .A(n180), .Z(n179) );
  HS65_LS_BFX9 U180 ( .A(n181), .Z(n180) );
  HS65_LS_BFX9 U181 ( .A(n182), .Z(n181) );
  HS65_LS_BFX9 U182 ( .A(n183), .Z(n182) );
  HS65_LS_BFX9 U183 ( .A(n184), .Z(n183) );
  HS65_LS_BFX9 U184 ( .A(north_in_ack0[1]), .Z(n184) );
  HS65_LS_BFX9 U185 ( .A(n186), .Z(n185) );
  HS65_LS_BFX9 U186 ( .A(n187), .Z(n186) );
  HS65_LS_BFX9 U187 ( .A(n188), .Z(n187) );
  HS65_LS_BFX9 U188 ( .A(n189), .Z(n188) );
  HS65_LS_BFX9 U189 ( .A(n190), .Z(n189) );
  HS65_LS_BFX9 U190 ( .A(n191), .Z(n190) );
  HS65_LS_BFX9 U191 ( .A(n192), .Z(n191) );
  HS65_LS_BFX9 U192 ( .A(west_in_ack0[1]), .Z(n192) );
  HS65_LS_BFX9 U193 ( .A(n194), .Z(n193) );
  HS65_LS_BFX9 U194 ( .A(n195), .Z(n194) );
  HS65_LS_BFX9 U195 ( .A(n196), .Z(n195) );
  HS65_LS_BFX9 U196 ( .A(n197), .Z(n196) );
  HS65_LS_BFX9 U197 ( .A(n198), .Z(n197) );
  HS65_LS_BFX9 U198 ( .A(n199), .Z(n198) );
  HS65_LS_BFX9 U199 ( .A(n200), .Z(n199) );
  HS65_LS_BFX9 U200 ( .A(north_in_ack0[2]), .Z(n200) );
  HS65_LS_BFX9 U201 ( .A(n202), .Z(n201) );
  HS65_LS_BFX9 U202 ( .A(n203), .Z(n202) );
  HS65_LS_BFX9 U203 ( .A(n204), .Z(n203) );
  HS65_LS_BFX9 U204 ( .A(n205), .Z(n204) );
  HS65_LS_BFX9 U205 ( .A(n206), .Z(n205) );
  HS65_LS_BFX9 U206 ( .A(n207), .Z(n206) );
  HS65_LS_BFX9 U207 ( .A(n208), .Z(n207) );
  HS65_LS_BFX9 U208 ( .A(east_in_ack0[1]), .Z(n208) );
  HS65_LS_BFX9 U209 ( .A(n210), .Z(n209) );
  HS65_LS_BFX9 U210 ( .A(n211), .Z(n210) );
  HS65_LS_BFX9 U211 ( .A(n212), .Z(n211) );
  HS65_LS_BFX9 U212 ( .A(n213), .Z(n212) );
  HS65_LS_BFX9 U213 ( .A(n214), .Z(n213) );
  HS65_LS_BFX9 U214 ( .A(n215), .Z(n214) );
  HS65_LS_BFX9 U215 ( .A(n216), .Z(n215) );
  HS65_LS_BFX9 U216 ( .A(south_out_req0[2]), .Z(n216) );
  HS65_LS_BFX9 U217 ( .A(n218), .Z(n217) );
  HS65_LS_BFX9 U218 ( .A(n219), .Z(n218) );
  HS65_LS_BFX9 U219 ( .A(n220), .Z(n219) );
  HS65_LS_BFX9 U220 ( .A(n221), .Z(n220) );
  HS65_LS_BFX9 U221 ( .A(n222), .Z(n221) );
  HS65_LS_BFX9 U222 ( .A(n223), .Z(n222) );
  HS65_LS_BFX9 U223 ( .A(n224), .Z(n223) );
  HS65_LS_BFX9 U224 ( .A(south_in_ack0[3]), .Z(n224) );
  HS65_LS_BFX9 U225 ( .A(n226), .Z(n225) );
  HS65_LS_BFX9 U226 ( .A(n227), .Z(n226) );
  HS65_LS_BFX9 U227 ( .A(n228), .Z(n227) );
  HS65_LS_BFX9 U228 ( .A(n229), .Z(n228) );
  HS65_LS_BFX9 U229 ( .A(n230), .Z(n229) );
  HS65_LS_BFX9 U230 ( .A(n231), .Z(n230) );
  HS65_LS_BFX9 U231 ( .A(n232), .Z(n231) );
  HS65_LS_BFX9 U232 ( .A(west_in_ack0[0]), .Z(n232) );
  HS65_LS_BFX9 U233 ( .A(n234), .Z(n233) );
  HS65_LS_BFX9 U234 ( .A(n235), .Z(n234) );
  HS65_LS_BFX9 U235 ( .A(n236), .Z(n235) );
  HS65_LS_BFX9 U236 ( .A(n237), .Z(n236) );
  HS65_LS_BFX9 U237 ( .A(n238), .Z(n237) );
  HS65_LS_BFX9 U238 ( .A(n239), .Z(n238) );
  HS65_LS_BFX9 U239 ( .A(n240), .Z(n239) );
  HS65_LS_BFX9 U240 ( .A(north_in_ack0[3]), .Z(n240) );
  HS65_LS_BFX9 U241 ( .A(n242), .Z(n241) );
  HS65_LS_BFX9 U242 ( .A(n243), .Z(n242) );
  HS65_LS_BFX9 U243 ( .A(n244), .Z(n243) );
  HS65_LS_BFX9 U244 ( .A(n245), .Z(n244) );
  HS65_LS_BFX9 U245 ( .A(n246), .Z(n245) );
  HS65_LS_BFX9 U246 ( .A(n247), .Z(n246) );
  HS65_LS_BFX9 U247 ( .A(n248), .Z(n247) );
  HS65_LS_BFX9 U248 ( .A(east_in_ack0[0]), .Z(n248) );
  HS65_LS_BFX9 U249 ( .A(n250), .Z(n249) );
  HS65_LS_BFX9 U250 ( .A(n251), .Z(n250) );
  HS65_LS_BFX9 U251 ( .A(n252), .Z(n251) );
  HS65_LS_BFX9 U252 ( .A(n253), .Z(n252) );
  HS65_LS_BFX9 U253 ( .A(n254), .Z(n253) );
  HS65_LS_BFX9 U254 ( .A(n255), .Z(n254) );
  HS65_LS_BFX9 U255 ( .A(n256), .Z(n255) );
  HS65_LS_BFX9 U256 ( .A(south_in_ack0[2]), .Z(n256) );
endmodule

