##
## LEF for PtnCells ;
## created by Encounter v13.13-s017_1 on Thu Mar 20 12:06:46 2014
##

VERSION 5.6 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO spm
  CLASS BLOCK ;
  FOREIGN spm 0 0 ;
  ORIGIN 0.0000 0.0000 ;
  SIZE 500.0000 BY 208.0000 ;
  SYMMETRY X Y R90 ;
  PIN a_spm_slave[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 156.7500 207.4800 156.8500 208.0000 ;
    END
  END a_spm_slave[63]
  PIN a_spm_slave[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 155.7500 207.4800 155.8500 208.0000 ;
    END
  END a_spm_slave[62]
  PIN a_spm_slave[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.7500 207.4800 154.8500 208.0000 ;
    END
  END a_spm_slave[61]
  PIN a_spm_slave[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.7500 207.4800 153.8500 208.0000 ;
    END
  END a_spm_slave[60]
  PIN a_spm_slave[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.7500 207.4800 152.8500 208.0000 ;
    END
  END a_spm_slave[59]
  PIN a_spm_slave[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 151.7500 207.4800 151.8500 208.0000 ;
    END
  END a_spm_slave[58]
  PIN a_spm_slave[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.7500 207.4800 150.8500 208.0000 ;
    END
  END a_spm_slave[57]
  PIN a_spm_slave[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 149.7500 207.4800 149.8500 208.0000 ;
    END
  END a_spm_slave[56]
  PIN a_spm_slave[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.7500 207.4800 148.8500 208.0000 ;
    END
  END a_spm_slave[55]
  PIN a_spm_slave[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 147.7500 207.4800 147.8500 208.0000 ;
    END
  END a_spm_slave[54]
  PIN a_spm_slave[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.7500 207.4800 146.8500 208.0000 ;
    END
  END a_spm_slave[53]
  PIN a_spm_slave[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.7500 207.4800 145.8500 208.0000 ;
    END
  END a_spm_slave[52]
  PIN a_spm_slave[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.7500 207.4800 144.8500 208.0000 ;
    END
  END a_spm_slave[51]
  PIN a_spm_slave[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 143.7500 207.4800 143.8500 208.0000 ;
    END
  END a_spm_slave[50]
  PIN a_spm_slave[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.7500 207.4800 142.8500 208.0000 ;
    END
  END a_spm_slave[49]
  PIN a_spm_slave[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.7500 207.4800 141.8500 208.0000 ;
    END
  END a_spm_slave[48]
  PIN a_spm_slave[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 140.7500 207.4800 140.8500 208.0000 ;
    END
  END a_spm_slave[47]
  PIN a_spm_slave[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.7500 207.4800 139.8500 208.0000 ;
    END
  END a_spm_slave[46]
  PIN a_spm_slave[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.7500 207.4800 138.8500 208.0000 ;
    END
  END a_spm_slave[45]
  PIN a_spm_slave[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.7500 207.4800 137.8500 208.0000 ;
    END
  END a_spm_slave[44]
  PIN a_spm_slave[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 136.7500 207.4800 136.8500 208.0000 ;
    END
  END a_spm_slave[43]
  PIN a_spm_slave[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 135.7500 207.4800 135.8500 208.0000 ;
    END
  END a_spm_slave[42]
  PIN a_spm_slave[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.7500 207.4800 134.8500 208.0000 ;
    END
  END a_spm_slave[41]
  PIN a_spm_slave[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 133.7500 207.4800 133.8500 208.0000 ;
    END
  END a_spm_slave[40]
  PIN a_spm_slave[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.7500 207.4800 132.8500 208.0000 ;
    END
  END a_spm_slave[39]
  PIN a_spm_slave[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.7500 207.4800 131.8500 208.0000 ;
    END
  END a_spm_slave[38]
  PIN a_spm_slave[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.7500 207.4800 130.8500 208.0000 ;
    END
  END a_spm_slave[37]
  PIN a_spm_slave[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.7500 207.4800 129.8500 208.0000 ;
    END
  END a_spm_slave[36]
  PIN a_spm_slave[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.7500 207.4800 128.8500 208.0000 ;
    END
  END a_spm_slave[35]
  PIN a_spm_slave[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 127.7500 207.4800 127.8500 208.0000 ;
    END
  END a_spm_slave[34]
  PIN a_spm_slave[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.7500 207.4800 126.8500 208.0000 ;
    END
  END a_spm_slave[33]
  PIN a_spm_slave[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.7500 207.4800 125.8500 208.0000 ;
    END
  END a_spm_slave[32]
  PIN a_spm_slave[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.7500 207.4800 124.8500 208.0000 ;
    END
  END a_spm_slave[31]
  PIN a_spm_slave[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.7500 207.4800 123.8500 208.0000 ;
    END
  END a_spm_slave[30]
  PIN a_spm_slave[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.7500 207.4800 122.8500 208.0000 ;
    END
  END a_spm_slave[29]
  PIN a_spm_slave[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 121.7500 207.4800 121.8500 208.0000 ;
    END
  END a_spm_slave[28]
  PIN a_spm_slave[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.7500 207.4800 120.8500 208.0000 ;
    END
  END a_spm_slave[27]
  PIN a_spm_slave[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.7500 207.4800 119.8500 208.0000 ;
    END
  END a_spm_slave[26]
  PIN a_spm_slave[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 118.7500 207.4800 118.8500 208.0000 ;
    END
  END a_spm_slave[25]
  PIN a_spm_slave[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.7500 207.4800 117.8500 208.0000 ;
    END
  END a_spm_slave[24]
  PIN a_spm_slave[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 116.7500 207.4800 116.8500 208.0000 ;
    END
  END a_spm_slave[23]
  PIN a_spm_slave[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.7500 207.4800 115.8500 208.0000 ;
    END
  END a_spm_slave[22]
  PIN a_spm_slave[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.7500 207.4800 114.8500 208.0000 ;
    END
  END a_spm_slave[21]
  PIN a_spm_slave[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 113.7500 207.4800 113.8500 208.0000 ;
    END
  END a_spm_slave[20]
  PIN a_spm_slave[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.7500 207.4800 112.8500 208.0000 ;
    END
  END a_spm_slave[19]
  PIN a_spm_slave[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.7500 207.4800 111.8500 208.0000 ;
    END
  END a_spm_slave[18]
  PIN a_spm_slave[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.7500 207.4800 110.8500 208.0000 ;
    END
  END a_spm_slave[17]
  PIN a_spm_slave[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.7500 207.4800 109.8500 208.0000 ;
    END
  END a_spm_slave[16]
  PIN a_spm_slave[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.7500 207.4800 108.8500 208.0000 ;
    END
  END a_spm_slave[15]
  PIN a_spm_slave[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.7500 207.4800 107.8500 208.0000 ;
    END
  END a_spm_slave[14]
  PIN a_spm_slave[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.7500 207.4800 106.8500 208.0000 ;
    END
  END a_spm_slave[13]
  PIN a_spm_slave[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.7500 207.4800 105.8500 208.0000 ;
    END
  END a_spm_slave[12]
  PIN a_spm_slave[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.7500 207.4800 104.8500 208.0000 ;
    END
  END a_spm_slave[11]
  PIN a_spm_slave[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.7500 207.4800 103.8500 208.0000 ;
    END
  END a_spm_slave[10]
  PIN a_spm_slave[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.7500 207.4800 102.8500 208.0000 ;
    END
  END a_spm_slave[9]
  PIN a_spm_slave[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.7500 207.4800 101.8500 208.0000 ;
    END
  END a_spm_slave[8]
  PIN a_spm_slave[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.7500 207.4800 100.8500 208.0000 ;
    END
  END a_spm_slave[7]
  PIN a_spm_slave[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.7500 207.4800 99.8500 208.0000 ;
    END
  END a_spm_slave[6]
  PIN a_spm_slave[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.7500 207.4800 98.8500 208.0000 ;
    END
  END a_spm_slave[5]
  PIN a_spm_slave[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.7500 207.4800 97.8500 208.0000 ;
    END
  END a_spm_slave[4]
  PIN a_spm_slave[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.7500 207.4800 96.8500 208.0000 ;
    END
  END a_spm_slave[3]
  PIN a_spm_slave[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.7500 207.4800 95.8500 208.0000 ;
    END
  END a_spm_slave[2]
  PIN a_spm_slave[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.7500 207.4800 94.8500 208.0000 ;
    END
  END a_spm_slave[1]
  PIN a_spm_slave[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.7500 207.4800 93.8500 208.0000 ;
    END
  END a_spm_slave[0]
  PIN a_spm_master[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92.7500 207.4800 92.8500 208.0000 ;
    END
  END a_spm_master[72]
  PIN a_spm_master[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 91.7500 207.4800 91.8500 208.0000 ;
    END
  END a_spm_master[71]
  PIN a_spm_master[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.7500 207.4800 90.8500 208.0000 ;
    END
  END a_spm_master[70]
  PIN a_spm_master[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.7500 207.4800 89.8500 208.0000 ;
    END
  END a_spm_master[69]
  PIN a_spm_master[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.7500 207.4800 88.8500 208.0000 ;
    END
  END a_spm_master[68]
  PIN a_spm_master[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.7500 207.4800 87.8500 208.0000 ;
    END
  END a_spm_master[67]
  PIN a_spm_master[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.7500 207.4800 86.8500 208.0000 ;
    END
  END a_spm_master[66]
  PIN a_spm_master[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.7500 207.4800 85.8500 208.0000 ;
    END
  END a_spm_master[65]
  PIN a_spm_master[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 84.7500 207.4800 84.8500 208.0000 ;
    END
  END a_spm_master[64]
  PIN a_spm_master[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.7500 207.4800 83.8500 208.0000 ;
    END
  END a_spm_master[63]
  PIN a_spm_master[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.7500 207.4800 82.8500 208.0000 ;
    END
  END a_spm_master[62]
  PIN a_spm_master[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.7500 207.4800 81.8500 208.0000 ;
    END
  END a_spm_master[61]
  PIN a_spm_master[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.7500 207.4800 80.8500 208.0000 ;
    END
  END a_spm_master[60]
  PIN a_spm_master[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.7500 207.4800 79.8500 208.0000 ;
    END
  END a_spm_master[59]
  PIN a_spm_master[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.7500 207.4800 78.8500 208.0000 ;
    END
  END a_spm_master[58]
  PIN a_spm_master[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.7500 207.4800 77.8500 208.0000 ;
    END
  END a_spm_master[57]
  PIN a_spm_master[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.7500 207.4800 76.8500 208.0000 ;
    END
  END a_spm_master[56]
  PIN a_spm_master[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.7500 207.4800 75.8500 208.0000 ;
    END
  END a_spm_master[55]
  PIN a_spm_master[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.7500 207.4800 74.8500 208.0000 ;
    END
  END a_spm_master[54]
  PIN a_spm_master[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.7500 207.4800 73.8500 208.0000 ;
    END
  END a_spm_master[53]
  PIN a_spm_master[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.7500 207.4800 72.8500 208.0000 ;
    END
  END a_spm_master[52]
  PIN a_spm_master[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.7500 207.4800 71.8500 208.0000 ;
    END
  END a_spm_master[51]
  PIN a_spm_master[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.7500 207.4800 70.8500 208.0000 ;
    END
  END a_spm_master[50]
  PIN a_spm_master[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.7500 207.4800 69.8500 208.0000 ;
    END
  END a_spm_master[49]
  PIN a_spm_master[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.7500 207.4800 68.8500 208.0000 ;
    END
  END a_spm_master[48]
  PIN a_spm_master[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.7500 207.4800 67.8500 208.0000 ;
    END
  END a_spm_master[47]
  PIN a_spm_master[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.7500 207.4800 66.8500 208.0000 ;
    END
  END a_spm_master[46]
  PIN a_spm_master[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.7500 207.4800 65.8500 208.0000 ;
    END
  END a_spm_master[45]
  PIN a_spm_master[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.7500 207.4800 64.8500 208.0000 ;
    END
  END a_spm_master[44]
  PIN a_spm_master[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.7500 207.4800 63.8500 208.0000 ;
    END
  END a_spm_master[43]
  PIN a_spm_master[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.7500 207.4800 62.8500 208.0000 ;
    END
  END a_spm_master[42]
  PIN a_spm_master[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.7500 207.4800 61.8500 208.0000 ;
    END
  END a_spm_master[41]
  PIN a_spm_master[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.7500 207.4800 60.8500 208.0000 ;
    END
  END a_spm_master[40]
  PIN a_spm_master[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.7500 207.4800 59.8500 208.0000 ;
    END
  END a_spm_master[39]
  PIN a_spm_master[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.7500 207.4800 58.8500 208.0000 ;
    END
  END a_spm_master[38]
  PIN a_spm_master[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.7500 207.4800 57.8500 208.0000 ;
    END
  END a_spm_master[37]
  PIN a_spm_master[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.7500 207.4800 56.8500 208.0000 ;
    END
  END a_spm_master[36]
  PIN a_spm_master[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.7500 207.4800 55.8500 208.0000 ;
    END
  END a_spm_master[35]
  PIN a_spm_master[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.7500 207.4800 54.8500 208.0000 ;
    END
  END a_spm_master[34]
  PIN a_spm_master[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.7500 207.4800 53.8500 208.0000 ;
    END
  END a_spm_master[33]
  PIN a_spm_master[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.7500 207.4800 52.8500 208.0000 ;
    END
  END a_spm_master[32]
  PIN a_spm_master[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.7500 207.4800 51.8500 208.0000 ;
    END
  END a_spm_master[31]
  PIN a_spm_master[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.7500 207.4800 50.8500 208.0000 ;
    END
  END a_spm_master[30]
  PIN a_spm_master[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.7500 207.4800 49.8500 208.0000 ;
    END
  END a_spm_master[29]
  PIN a_spm_master[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.7500 207.4800 48.8500 208.0000 ;
    END
  END a_spm_master[28]
  PIN a_spm_master[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.7500 207.4800 47.8500 208.0000 ;
    END
  END a_spm_master[27]
  PIN a_spm_master[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.7500 207.4800 46.8500 208.0000 ;
    END
  END a_spm_master[26]
  PIN a_spm_master[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.7500 207.4800 45.8500 208.0000 ;
    END
  END a_spm_master[25]
  PIN a_spm_master[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.7500 207.4800 44.8500 208.0000 ;
    END
  END a_spm_master[24]
  PIN a_spm_master[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.7500 207.4800 43.8500 208.0000 ;
    END
  END a_spm_master[23]
  PIN a_spm_master[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.7500 207.4800 42.8500 208.0000 ;
    END
  END a_spm_master[22]
  PIN a_spm_master[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.7500 207.4800 41.8500 208.0000 ;
    END
  END a_spm_master[21]
  PIN a_spm_master[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.7500 207.4800 40.8500 208.0000 ;
    END
  END a_spm_master[20]
  PIN a_spm_master[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.7500 207.4800 39.8500 208.0000 ;
    END
  END a_spm_master[19]
  PIN a_spm_master[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.7500 207.4800 38.8500 208.0000 ;
    END
  END a_spm_master[18]
  PIN a_spm_master[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.7500 207.4800 37.8500 208.0000 ;
    END
  END a_spm_master[17]
  PIN a_spm_master[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.7500 207.4800 36.8500 208.0000 ;
    END
  END a_spm_master[16]
  PIN a_spm_master[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.7500 207.4800 35.8500 208.0000 ;
    END
  END a_spm_master[15]
  PIN a_spm_master[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.7500 207.4800 34.8500 208.0000 ;
    END
  END a_spm_master[14]
  PIN a_spm_master[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.7500 207.4800 33.8500 208.0000 ;
    END
  END a_spm_master[13]
  PIN a_spm_master[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.7500 207.4800 32.8500 208.0000 ;
    END
  END a_spm_master[12]
  PIN a_spm_master[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.7500 207.4800 31.8500 208.0000 ;
    END
  END a_spm_master[11]
  PIN a_spm_master[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.7500 207.4800 30.8500 208.0000 ;
    END
  END a_spm_master[10]
  PIN a_spm_master[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.7500 207.4800 29.8500 208.0000 ;
    END
  END a_spm_master[9]
  PIN a_spm_master[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.7500 207.4800 28.8500 208.0000 ;
    END
  END a_spm_master[8]
  PIN a_spm_master[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.7500 207.4800 27.8500 208.0000 ;
    END
  END a_spm_master[7]
  PIN a_spm_master[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.7500 207.4800 26.8500 208.0000 ;
    END
  END a_spm_master[6]
  PIN a_spm_master[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.7500 207.4800 25.8500 208.0000 ;
    END
  END a_spm_master[5]
  PIN a_spm_master[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.7500 207.4800 24.8500 208.0000 ;
    END
  END a_spm_master[4]
  PIN a_spm_master[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.7500 207.4800 23.8500 208.0000 ;
    END
  END a_spm_master[3]
  PIN a_spm_master[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.7500 207.4800 22.8500 208.0000 ;
    END
  END a_spm_master[2]
  PIN a_spm_master[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.7500 207.4800 21.8500 208.0000 ;
    END
  END a_spm_master[1]
  PIN a_spm_master[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.7500 207.4800 20.8500 208.0000 ;
    END
  END a_spm_master[0]
  PIN b_spm_slave[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 138.3500 0.5200 138.4500 ;
    END
  END b_spm_slave[63]
  PIN b_spm_slave[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 137.3500 0.5200 137.4500 ;
    END
  END b_spm_slave[62]
  PIN b_spm_slave[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 136.3500 0.5200 136.4500 ;
    END
  END b_spm_slave[61]
  PIN b_spm_slave[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 135.3500 0.5200 135.4500 ;
    END
  END b_spm_slave[60]
  PIN b_spm_slave[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 134.3500 0.5200 134.4500 ;
    END
  END b_spm_slave[59]
  PIN b_spm_slave[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 133.3500 0.5200 133.4500 ;
    END
  END b_spm_slave[58]
  PIN b_spm_slave[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 132.3500 0.5200 132.4500 ;
    END
  END b_spm_slave[57]
  PIN b_spm_slave[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 131.3500 0.5200 131.4500 ;
    END
  END b_spm_slave[56]
  PIN b_spm_slave[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 130.3500 0.5200 130.4500 ;
    END
  END b_spm_slave[55]
  PIN b_spm_slave[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 129.3500 0.5200 129.4500 ;
    END
  END b_spm_slave[54]
  PIN b_spm_slave[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 128.3500 0.5200 128.4500 ;
    END
  END b_spm_slave[53]
  PIN b_spm_slave[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 127.3500 0.5200 127.4500 ;
    END
  END b_spm_slave[52]
  PIN b_spm_slave[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 126.3500 0.5200 126.4500 ;
    END
  END b_spm_slave[51]
  PIN b_spm_slave[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 125.3500 0.5200 125.4500 ;
    END
  END b_spm_slave[50]
  PIN b_spm_slave[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 124.3500 0.5200 124.4500 ;
    END
  END b_spm_slave[49]
  PIN b_spm_slave[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 123.3500 0.5200 123.4500 ;
    END
  END b_spm_slave[48]
  PIN b_spm_slave[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 122.3500 0.5200 122.4500 ;
    END
  END b_spm_slave[47]
  PIN b_spm_slave[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 121.3500 0.5200 121.4500 ;
    END
  END b_spm_slave[46]
  PIN b_spm_slave[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 120.3500 0.5200 120.4500 ;
    END
  END b_spm_slave[45]
  PIN b_spm_slave[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 119.3500 0.5200 119.4500 ;
    END
  END b_spm_slave[44]
  PIN b_spm_slave[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 118.3500 0.5200 118.4500 ;
    END
  END b_spm_slave[43]
  PIN b_spm_slave[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 117.3500 0.5200 117.4500 ;
    END
  END b_spm_slave[42]
  PIN b_spm_slave[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 116.3500 0.5200 116.4500 ;
    END
  END b_spm_slave[41]
  PIN b_spm_slave[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 115.3500 0.5200 115.4500 ;
    END
  END b_spm_slave[40]
  PIN b_spm_slave[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 114.3500 0.5200 114.4500 ;
    END
  END b_spm_slave[39]
  PIN b_spm_slave[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 113.3500 0.5200 113.4500 ;
    END
  END b_spm_slave[38]
  PIN b_spm_slave[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 112.3500 0.5200 112.4500 ;
    END
  END b_spm_slave[37]
  PIN b_spm_slave[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 111.3500 0.5200 111.4500 ;
    END
  END b_spm_slave[36]
  PIN b_spm_slave[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 110.3500 0.5200 110.4500 ;
    END
  END b_spm_slave[35]
  PIN b_spm_slave[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 109.3500 0.5200 109.4500 ;
    END
  END b_spm_slave[34]
  PIN b_spm_slave[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 108.3500 0.5200 108.4500 ;
    END
  END b_spm_slave[33]
  PIN b_spm_slave[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 107.3500 0.5200 107.4500 ;
    END
  END b_spm_slave[32]
  PIN b_spm_slave[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 106.3500 0.5200 106.4500 ;
    END
  END b_spm_slave[31]
  PIN b_spm_slave[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 105.3500 0.5200 105.4500 ;
    END
  END b_spm_slave[30]
  PIN b_spm_slave[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 104.3500 0.5200 104.4500 ;
    END
  END b_spm_slave[29]
  PIN b_spm_slave[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 103.3500 0.5200 103.4500 ;
    END
  END b_spm_slave[28]
  PIN b_spm_slave[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 102.3500 0.5200 102.4500 ;
    END
  END b_spm_slave[27]
  PIN b_spm_slave[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 101.3500 0.5200 101.4500 ;
    END
  END b_spm_slave[26]
  PIN b_spm_slave[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 100.3500 0.5200 100.4500 ;
    END
  END b_spm_slave[25]
  PIN b_spm_slave[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 99.3500 0.5200 99.4500 ;
    END
  END b_spm_slave[24]
  PIN b_spm_slave[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 98.3500 0.5200 98.4500 ;
    END
  END b_spm_slave[23]
  PIN b_spm_slave[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 97.3500 0.5200 97.4500 ;
    END
  END b_spm_slave[22]
  PIN b_spm_slave[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 96.3500 0.5200 96.4500 ;
    END
  END b_spm_slave[21]
  PIN b_spm_slave[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 95.3500 0.5200 95.4500 ;
    END
  END b_spm_slave[20]
  PIN b_spm_slave[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 94.3500 0.5200 94.4500 ;
    END
  END b_spm_slave[19]
  PIN b_spm_slave[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 93.3500 0.5200 93.4500 ;
    END
  END b_spm_slave[18]
  PIN b_spm_slave[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 92.3500 0.5200 92.4500 ;
    END
  END b_spm_slave[17]
  PIN b_spm_slave[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 91.3500 0.5200 91.4500 ;
    END
  END b_spm_slave[16]
  PIN b_spm_slave[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 90.3500 0.5200 90.4500 ;
    END
  END b_spm_slave[15]
  PIN b_spm_slave[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 89.3500 0.5200 89.4500 ;
    END
  END b_spm_slave[14]
  PIN b_spm_slave[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 88.3500 0.5200 88.4500 ;
    END
  END b_spm_slave[13]
  PIN b_spm_slave[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 87.3500 0.5200 87.4500 ;
    END
  END b_spm_slave[12]
  PIN b_spm_slave[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 86.3500 0.5200 86.4500 ;
    END
  END b_spm_slave[11]
  PIN b_spm_slave[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 85.3500 0.5200 85.4500 ;
    END
  END b_spm_slave[10]
  PIN b_spm_slave[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 84.3500 0.5200 84.4500 ;
    END
  END b_spm_slave[9]
  PIN b_spm_slave[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 83.3500 0.5200 83.4500 ;
    END
  END b_spm_slave[8]
  PIN b_spm_slave[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 82.3500 0.5200 82.4500 ;
    END
  END b_spm_slave[7]
  PIN b_spm_slave[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 81.3500 0.5200 81.4500 ;
    END
  END b_spm_slave[6]
  PIN b_spm_slave[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 80.3500 0.5200 80.4500 ;
    END
  END b_spm_slave[5]
  PIN b_spm_slave[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 79.3500 0.5200 79.4500 ;
    END
  END b_spm_slave[4]
  PIN b_spm_slave[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 78.3500 0.5200 78.4500 ;
    END
  END b_spm_slave[3]
  PIN b_spm_slave[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 77.3500 0.5200 77.4500 ;
    END
  END b_spm_slave[2]
  PIN b_spm_slave[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 76.3500 0.5200 76.4500 ;
    END
  END b_spm_slave[1]
  PIN b_spm_slave[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 75.3500 0.5200 75.4500 ;
    END
  END b_spm_slave[0]
  PIN b_spm_master[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 74.3500 0.5200 74.4500 ;
    END
  END b_spm_master[72]
  PIN b_spm_master[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 73.3500 0.5200 73.4500 ;
    END
  END b_spm_master[71]
  PIN b_spm_master[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 72.3500 0.5200 72.4500 ;
    END
  END b_spm_master[70]
  PIN b_spm_master[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 71.3500 0.5200 71.4500 ;
    END
  END b_spm_master[69]
  PIN b_spm_master[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 70.3500 0.5200 70.4500 ;
    END
  END b_spm_master[68]
  PIN b_spm_master[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 69.3500 0.5200 69.4500 ;
    END
  END b_spm_master[67]
  PIN b_spm_master[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 68.3500 0.5200 68.4500 ;
    END
  END b_spm_master[66]
  PIN b_spm_master[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 67.3500 0.5200 67.4500 ;
    END
  END b_spm_master[65]
  PIN b_spm_master[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 66.3500 0.5200 66.4500 ;
    END
  END b_spm_master[64]
  PIN b_spm_master[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 65.3500 0.5200 65.4500 ;
    END
  END b_spm_master[63]
  PIN b_spm_master[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 64.3500 0.5200 64.4500 ;
    END
  END b_spm_master[62]
  PIN b_spm_master[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 63.3500 0.5200 63.4500 ;
    END
  END b_spm_master[61]
  PIN b_spm_master[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 62.3500 0.5200 62.4500 ;
    END
  END b_spm_master[60]
  PIN b_spm_master[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 61.3500 0.5200 61.4500 ;
    END
  END b_spm_master[59]
  PIN b_spm_master[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 60.3500 0.5200 60.4500 ;
    END
  END b_spm_master[58]
  PIN b_spm_master[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 59.3500 0.5200 59.4500 ;
    END
  END b_spm_master[57]
  PIN b_spm_master[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 58.3500 0.5200 58.4500 ;
    END
  END b_spm_master[56]
  PIN b_spm_master[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 57.3500 0.5200 57.4500 ;
    END
  END b_spm_master[55]
  PIN b_spm_master[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 56.3500 0.5200 56.4500 ;
    END
  END b_spm_master[54]
  PIN b_spm_master[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 55.3500 0.5200 55.4500 ;
    END
  END b_spm_master[53]
  PIN b_spm_master[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 54.3500 0.5200 54.4500 ;
    END
  END b_spm_master[52]
  PIN b_spm_master[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 53.3500 0.5200 53.4500 ;
    END
  END b_spm_master[51]
  PIN b_spm_master[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 52.3500 0.5200 52.4500 ;
    END
  END b_spm_master[50]
  PIN b_spm_master[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 51.3500 0.5200 51.4500 ;
    END
  END b_spm_master[49]
  PIN b_spm_master[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 50.3500 0.5200 50.4500 ;
    END
  END b_spm_master[48]
  PIN b_spm_master[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 49.3500 0.5200 49.4500 ;
    END
  END b_spm_master[47]
  PIN b_spm_master[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 48.3500 0.5200 48.4500 ;
    END
  END b_spm_master[46]
  PIN b_spm_master[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 47.3500 0.5200 47.4500 ;
    END
  END b_spm_master[45]
  PIN b_spm_master[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 46.3500 0.5200 46.4500 ;
    END
  END b_spm_master[44]
  PIN b_spm_master[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 45.3500 0.5200 45.4500 ;
    END
  END b_spm_master[43]
  PIN b_spm_master[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 44.3500 0.5200 44.4500 ;
    END
  END b_spm_master[42]
  PIN b_spm_master[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 43.3500 0.5200 43.4500 ;
    END
  END b_spm_master[41]
  PIN b_spm_master[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 42.3500 0.5200 42.4500 ;
    END
  END b_spm_master[40]
  PIN b_spm_master[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 41.3500 0.5200 41.4500 ;
    END
  END b_spm_master[39]
  PIN b_spm_master[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 40.3500 0.5200 40.4500 ;
    END
  END b_spm_master[38]
  PIN b_spm_master[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 39.3500 0.5200 39.4500 ;
    END
  END b_spm_master[37]
  PIN b_spm_master[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 38.3500 0.5200 38.4500 ;
    END
  END b_spm_master[36]
  PIN b_spm_master[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 37.3500 0.5200 37.4500 ;
    END
  END b_spm_master[35]
  PIN b_spm_master[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 36.3500 0.5200 36.4500 ;
    END
  END b_spm_master[34]
  PIN b_spm_master[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 35.3500 0.5200 35.4500 ;
    END
  END b_spm_master[33]
  PIN b_spm_master[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 34.3500 0.5200 34.4500 ;
    END
  END b_spm_master[32]
  PIN b_spm_master[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 33.3500 0.5200 33.4500 ;
    END
  END b_spm_master[31]
  PIN b_spm_master[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 32.3500 0.5200 32.4500 ;
    END
  END b_spm_master[30]
  PIN b_spm_master[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 31.3500 0.5200 31.4500 ;
    END
  END b_spm_master[29]
  PIN b_spm_master[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 30.3500 0.5200 30.4500 ;
    END
  END b_spm_master[28]
  PIN b_spm_master[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 29.3500 0.5200 29.4500 ;
    END
  END b_spm_master[27]
  PIN b_spm_master[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 28.3500 0.5200 28.4500 ;
    END
  END b_spm_master[26]
  PIN b_spm_master[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 27.3500 0.5200 27.4500 ;
    END
  END b_spm_master[25]
  PIN b_spm_master[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 26.3500 0.5200 26.4500 ;
    END
  END b_spm_master[24]
  PIN b_spm_master[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 25.3500 0.5200 25.4500 ;
    END
  END b_spm_master[23]
  PIN b_spm_master[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 24.3500 0.5200 24.4500 ;
    END
  END b_spm_master[22]
  PIN b_spm_master[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 23.3500 0.5200 23.4500 ;
    END
  END b_spm_master[21]
  PIN b_spm_master[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 22.3500 0.5200 22.4500 ;
    END
  END b_spm_master[20]
  PIN b_spm_master[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 21.3500 0.5200 21.4500 ;
    END
  END b_spm_master[19]
  PIN b_spm_master[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 20.3500 0.5200 20.4500 ;
    END
  END b_spm_master[18]
  PIN b_spm_master[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 19.3500 0.5200 19.4500 ;
    END
  END b_spm_master[17]
  PIN b_spm_master[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 18.3500 0.5200 18.4500 ;
    END
  END b_spm_master[16]
  PIN b_spm_master[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 17.3500 0.5200 17.4500 ;
    END
  END b_spm_master[15]
  PIN b_spm_master[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 16.3500 0.5200 16.4500 ;
    END
  END b_spm_master[14]
  PIN b_spm_master[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 15.3500 0.5200 15.4500 ;
    END
  END b_spm_master[13]
  PIN b_spm_master[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 14.3500 0.5200 14.4500 ;
    END
  END b_spm_master[12]
  PIN b_spm_master[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 13.3500 0.5200 13.4500 ;
    END
  END b_spm_master[11]
  PIN b_spm_master[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 12.3500 0.5200 12.4500 ;
    END
  END b_spm_master[10]
  PIN b_spm_master[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 11.3500 0.5200 11.4500 ;
    END
  END b_spm_master[9]
  PIN b_spm_master[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 10.3500 0.5200 10.4500 ;
    END
  END b_spm_master[8]
  PIN b_spm_master[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 9.3500 0.5200 9.4500 ;
    END
  END b_spm_master[7]
  PIN b_spm_master[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 8.3500 0.5200 8.4500 ;
    END
  END b_spm_master[6]
  PIN b_spm_master[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 7.3500 0.5200 7.4500 ;
    END
  END b_spm_master[5]
  PIN b_spm_master[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 6.3500 0.5200 6.4500 ;
    END
  END b_spm_master[4]
  PIN b_spm_master[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 5.3500 0.5200 5.4500 ;
    END
  END b_spm_master[3]
  PIN b_spm_master[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 4.3500 0.5200 4.4500 ;
    END
  END b_spm_master[2]
  PIN b_spm_master[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 3.3500 0.5200 3.4500 ;
    END
  END b_spm_master[1]
  PIN b_spm_master[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 2.3500 0.5200 2.4500 ;
    END
  END b_spm_master[0]
  PIN a_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 0.3500 0.5200 0.4500 ;
    END
  END a_clk
  PIN b_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 1.3500 0.5200 1.4500 ;
    END
  END b_clk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0000 139.3500 0.5200 139.4500 ;
    END
  END reset
  OBS
    LAYER OVERLAP ;
    LAYER AP ;
      RECT 0.0000 0.0000 500.0000 208.0000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 500.0000 208.0000 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 500.0000 208.0000 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 500.0000 208.0000 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 500.0000 208.0000 ;
    LAYER M3 ;
      RECT 0.0000 0.0000 500.0000 208.0000 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 500.0000 208.0000 ;
    LAYER M1 ;
      RECT 0.0000 0.0000 500.0000 208.0000 ;
  END
END spm

END LIBRARY
