##
## LEF for PtnCells ;
## created by Encounter v13.13-s017_1 on Thu Mar 20 12:06:46 2014
##

VERSION 5.6 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO processor
  CLASS BLOCK ;
  FOREIGN processor 0 0 ;
  ORIGIN 0.0000 0.0000 ;
  SIZE 1383.2000 BY 1175.2000 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1500 0.0000 0.2500 0.4200 ;
    END
  END clk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 116.1500 0.0000 116.2500 0.4200 ;
    END
  END reset
  PIN p_spm_master[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 394.3500 0.0000 394.4500 0.4200 ;
    END
  END p_spm_master[72]
  PIN p_spm_master[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 393.3500 0.0000 393.4500 0.4200 ;
    END
  END p_spm_master[71]
  PIN p_spm_master[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 392.3500 0.0000 392.4500 0.4200 ;
    END
  END p_spm_master[70]
  PIN p_spm_master[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 391.3500 0.0000 391.4500 0.4200 ;
    END
  END p_spm_master[69]
  PIN p_spm_master[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 390.3500 0.0000 390.4500 0.4200 ;
    END
  END p_spm_master[68]
  PIN p_spm_master[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 389.3500 0.0000 389.4500 0.4200 ;
    END
  END p_spm_master[67]
  PIN p_spm_master[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 388.3500 0.0000 388.4500 0.4200 ;
    END
  END p_spm_master[66]
  PIN p_spm_master[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 387.3500 0.0000 387.4500 0.4200 ;
    END
  END p_spm_master[65]
  PIN p_spm_master[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 386.3500 0.0000 386.4500 0.4200 ;
    END
  END p_spm_master[64]
  PIN p_spm_master[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 385.3500 0.0000 385.4500 0.4200 ;
    END
  END p_spm_master[63]
  PIN p_spm_master[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 384.3500 0.0000 384.4500 0.4200 ;
    END
  END p_spm_master[62]
  PIN p_spm_master[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 383.3500 0.0000 383.4500 0.4200 ;
    END
  END p_spm_master[61]
  PIN p_spm_master[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 382.3500 0.0000 382.4500 0.4200 ;
    END
  END p_spm_master[60]
  PIN p_spm_master[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 381.3500 0.0000 381.4500 0.4200 ;
    END
  END p_spm_master[59]
  PIN p_spm_master[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 380.3500 0.0000 380.4500 0.4200 ;
    END
  END p_spm_master[58]
  PIN p_spm_master[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 379.3500 0.0000 379.4500 0.4200 ;
    END
  END p_spm_master[57]
  PIN p_spm_master[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 378.3500 0.0000 378.4500 0.4200 ;
    END
  END p_spm_master[56]
  PIN p_spm_master[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 377.3500 0.0000 377.4500 0.4200 ;
    END
  END p_spm_master[55]
  PIN p_spm_master[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 376.3500 0.0000 376.4500 0.4200 ;
    END
  END p_spm_master[54]
  PIN p_spm_master[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 375.3500 0.0000 375.4500 0.4200 ;
    END
  END p_spm_master[53]
  PIN p_spm_master[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 374.3500 0.0000 374.4500 0.4200 ;
    END
  END p_spm_master[52]
  PIN p_spm_master[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 373.3500 0.0000 373.4500 0.4200 ;
    END
  END p_spm_master[51]
  PIN p_spm_master[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 372.3500 0.0000 372.4500 0.4200 ;
    END
  END p_spm_master[50]
  PIN p_spm_master[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 371.3500 0.0000 371.4500 0.4200 ;
    END
  END p_spm_master[49]
  PIN p_spm_master[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 370.3500 0.0000 370.4500 0.4200 ;
    END
  END p_spm_master[48]
  PIN p_spm_master[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 369.3500 0.0000 369.4500 0.4200 ;
    END
  END p_spm_master[47]
  PIN p_spm_master[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 368.3500 0.0000 368.4500 0.4200 ;
    END
  END p_spm_master[46]
  PIN p_spm_master[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 367.3500 0.0000 367.4500 0.4200 ;
    END
  END p_spm_master[45]
  PIN p_spm_master[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 366.3500 0.0000 366.4500 0.4200 ;
    END
  END p_spm_master[44]
  PIN p_spm_master[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 365.3500 0.0000 365.4500 0.4200 ;
    END
  END p_spm_master[43]
  PIN p_spm_master[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 364.3500 0.0000 364.4500 0.4200 ;
    END
  END p_spm_master[42]
  PIN p_spm_master[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 363.3500 0.0000 363.4500 0.4200 ;
    END
  END p_spm_master[41]
  PIN p_spm_master[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 362.3500 0.0000 362.4500 0.4200 ;
    END
  END p_spm_master[40]
  PIN p_spm_master[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 361.3500 0.0000 361.4500 0.4200 ;
    END
  END p_spm_master[39]
  PIN p_spm_master[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 360.3500 0.0000 360.4500 0.4200 ;
    END
  END p_spm_master[38]
  PIN p_spm_master[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 359.3500 0.0000 359.4500 0.4200 ;
    END
  END p_spm_master[37]
  PIN p_spm_master[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 358.3500 0.0000 358.4500 0.4200 ;
    END
  END p_spm_master[36]
  PIN p_spm_master[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 357.3500 0.0000 357.4500 0.4200 ;
    END
  END p_spm_master[35]
  PIN p_spm_master[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 356.3500 0.0000 356.4500 0.4200 ;
    END
  END p_spm_master[34]
  PIN p_spm_master[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 355.3500 0.0000 355.4500 0.4200 ;
    END
  END p_spm_master[33]
  PIN p_spm_master[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 354.3500 0.0000 354.4500 0.4200 ;
    END
  END p_spm_master[32]
  PIN p_spm_master[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 353.3500 0.0000 353.4500 0.4200 ;
    END
  END p_spm_master[31]
  PIN p_spm_master[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 352.3500 0.0000 352.4500 0.4200 ;
    END
  END p_spm_master[30]
  PIN p_spm_master[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 351.3500 0.0000 351.4500 0.4200 ;
    END
  END p_spm_master[29]
  PIN p_spm_master[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 350.3500 0.0000 350.4500 0.4200 ;
    END
  END p_spm_master[28]
  PIN p_spm_master[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 349.3500 0.0000 349.4500 0.4200 ;
    END
  END p_spm_master[27]
  PIN p_spm_master[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 348.3500 0.0000 348.4500 0.4200 ;
    END
  END p_spm_master[26]
  PIN p_spm_master[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 347.3500 0.0000 347.4500 0.4200 ;
    END
  END p_spm_master[25]
  PIN p_spm_master[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 346.3500 0.0000 346.4500 0.4200 ;
    END
  END p_spm_master[24]
  PIN p_spm_master[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 345.3500 0.0000 345.4500 0.4200 ;
    END
  END p_spm_master[23]
  PIN p_spm_master[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 344.3500 0.0000 344.4500 0.4200 ;
    END
  END p_spm_master[22]
  PIN p_spm_master[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 343.3500 0.0000 343.4500 0.4200 ;
    END
  END p_spm_master[21]
  PIN p_spm_master[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 342.3500 0.0000 342.4500 0.4200 ;
    END
  END p_spm_master[20]
  PIN p_spm_master[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 341.3500 0.0000 341.4500 0.4200 ;
    END
  END p_spm_master[19]
  PIN p_spm_master[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 340.3500 0.0000 340.4500 0.4200 ;
    END
  END p_spm_master[18]
  PIN p_spm_master[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 339.3500 0.0000 339.4500 0.4200 ;
    END
  END p_spm_master[17]
  PIN p_spm_master[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 338.3500 0.0000 338.4500 0.4200 ;
    END
  END p_spm_master[16]
  PIN p_spm_master[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 337.3500 0.0000 337.4500 0.4200 ;
    END
  END p_spm_master[15]
  PIN p_spm_master[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 336.3500 0.0000 336.4500 0.4200 ;
    END
  END p_spm_master[14]
  PIN p_spm_master[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 335.3500 0.0000 335.4500 0.4200 ;
    END
  END p_spm_master[13]
  PIN p_spm_master[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 334.3500 0.0000 334.4500 0.4200 ;
    END
  END p_spm_master[12]
  PIN p_spm_master[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 333.3500 0.0000 333.4500 0.4200 ;
    END
  END p_spm_master[11]
  PIN p_spm_master[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 332.3500 0.0000 332.4500 0.4200 ;
    END
  END p_spm_master[10]
  PIN p_spm_master[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 331.3500 0.0000 331.4500 0.4200 ;
    END
  END p_spm_master[9]
  PIN p_spm_master[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 330.3500 0.0000 330.4500 0.4200 ;
    END
  END p_spm_master[8]
  PIN p_spm_master[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 329.3500 0.0000 329.4500 0.4200 ;
    END
  END p_spm_master[7]
  PIN p_spm_master[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 328.3500 0.0000 328.4500 0.4200 ;
    END
  END p_spm_master[6]
  PIN p_spm_master[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 327.3500 0.0000 327.4500 0.4200 ;
    END
  END p_spm_master[5]
  PIN p_spm_master[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 326.3500 0.0000 326.4500 0.4200 ;
    END
  END p_spm_master[4]
  PIN p_spm_master[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 325.3500 0.0000 325.4500 0.4200 ;
    END
  END p_spm_master[3]
  PIN p_spm_master[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 324.3500 0.0000 324.4500 0.4200 ;
    END
  END p_spm_master[2]
  PIN p_spm_master[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 323.3500 0.0000 323.4500 0.4200 ;
    END
  END p_spm_master[1]
  PIN p_spm_master[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 322.3500 0.0000 322.4500 0.4200 ;
    END
  END p_spm_master[0]
  PIN p_spm_slave[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 458.3500 0.0000 458.4500 0.4200 ;
    END
  END p_spm_slave[63]
  PIN p_spm_slave[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 457.3500 0.0000 457.4500 0.4200 ;
    END
  END p_spm_slave[62]
  PIN p_spm_slave[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 456.3500 0.0000 456.4500 0.4200 ;
    END
  END p_spm_slave[61]
  PIN p_spm_slave[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 455.3500 0.0000 455.4500 0.4200 ;
    END
  END p_spm_slave[60]
  PIN p_spm_slave[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 454.3500 0.0000 454.4500 0.4200 ;
    END
  END p_spm_slave[59]
  PIN p_spm_slave[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 453.3500 0.0000 453.4500 0.4200 ;
    END
  END p_spm_slave[58]
  PIN p_spm_slave[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 452.3500 0.0000 452.4500 0.4200 ;
    END
  END p_spm_slave[57]
  PIN p_spm_slave[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 451.3500 0.0000 451.4500 0.4200 ;
    END
  END p_spm_slave[56]
  PIN p_spm_slave[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 450.3500 0.0000 450.4500 0.4200 ;
    END
  END p_spm_slave[55]
  PIN p_spm_slave[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 449.3500 0.0000 449.4500 0.4200 ;
    END
  END p_spm_slave[54]
  PIN p_spm_slave[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 448.3500 0.0000 448.4500 0.4200 ;
    END
  END p_spm_slave[53]
  PIN p_spm_slave[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 447.3500 0.0000 447.4500 0.4200 ;
    END
  END p_spm_slave[52]
  PIN p_spm_slave[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 446.3500 0.0000 446.4500 0.4200 ;
    END
  END p_spm_slave[51]
  PIN p_spm_slave[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 445.3500 0.0000 445.4500 0.4200 ;
    END
  END p_spm_slave[50]
  PIN p_spm_slave[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 444.3500 0.0000 444.4500 0.4200 ;
    END
  END p_spm_slave[49]
  PIN p_spm_slave[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 443.3500 0.0000 443.4500 0.4200 ;
    END
  END p_spm_slave[48]
  PIN p_spm_slave[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 442.3500 0.0000 442.4500 0.4200 ;
    END
  END p_spm_slave[47]
  PIN p_spm_slave[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 441.3500 0.0000 441.4500 0.4200 ;
    END
  END p_spm_slave[46]
  PIN p_spm_slave[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 440.3500 0.0000 440.4500 0.4200 ;
    END
  END p_spm_slave[45]
  PIN p_spm_slave[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 439.3500 0.0000 439.4500 0.4200 ;
    END
  END p_spm_slave[44]
  PIN p_spm_slave[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 438.3500 0.0000 438.4500 0.4200 ;
    END
  END p_spm_slave[43]
  PIN p_spm_slave[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 437.3500 0.0000 437.4500 0.4200 ;
    END
  END p_spm_slave[42]
  PIN p_spm_slave[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 436.3500 0.0000 436.4500 0.4200 ;
    END
  END p_spm_slave[41]
  PIN p_spm_slave[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 435.3500 0.0000 435.4500 0.4200 ;
    END
  END p_spm_slave[40]
  PIN p_spm_slave[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 434.3500 0.0000 434.4500 0.4200 ;
    END
  END p_spm_slave[39]
  PIN p_spm_slave[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 433.3500 0.0000 433.4500 0.4200 ;
    END
  END p_spm_slave[38]
  PIN p_spm_slave[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 432.3500 0.0000 432.4500 0.4200 ;
    END
  END p_spm_slave[37]
  PIN p_spm_slave[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 431.3500 0.0000 431.4500 0.4200 ;
    END
  END p_spm_slave[36]
  PIN p_spm_slave[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 430.3500 0.0000 430.4500 0.4200 ;
    END
  END p_spm_slave[35]
  PIN p_spm_slave[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 429.3500 0.0000 429.4500 0.4200 ;
    END
  END p_spm_slave[34]
  PIN p_spm_slave[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 428.3500 0.0000 428.4500 0.4200 ;
    END
  END p_spm_slave[33]
  PIN p_spm_slave[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 427.3500 0.0000 427.4500 0.4200 ;
    END
  END p_spm_slave[32]
  PIN p_spm_slave[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 426.3500 0.0000 426.4500 0.4200 ;
    END
  END p_spm_slave[31]
  PIN p_spm_slave[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 425.3500 0.0000 425.4500 0.4200 ;
    END
  END p_spm_slave[30]
  PIN p_spm_slave[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 424.3500 0.0000 424.4500 0.4200 ;
    END
  END p_spm_slave[29]
  PIN p_spm_slave[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 423.3500 0.0000 423.4500 0.4200 ;
    END
  END p_spm_slave[28]
  PIN p_spm_slave[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 422.3500 0.0000 422.4500 0.4200 ;
    END
  END p_spm_slave[27]
  PIN p_spm_slave[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 421.3500 0.0000 421.4500 0.4200 ;
    END
  END p_spm_slave[26]
  PIN p_spm_slave[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 420.3500 0.0000 420.4500 0.4200 ;
    END
  END p_spm_slave[25]
  PIN p_spm_slave[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 419.3500 0.0000 419.4500 0.4200 ;
    END
  END p_spm_slave[24]
  PIN p_spm_slave[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 418.3500 0.0000 418.4500 0.4200 ;
    END
  END p_spm_slave[23]
  PIN p_spm_slave[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 417.3500 0.0000 417.4500 0.4200 ;
    END
  END p_spm_slave[22]
  PIN p_spm_slave[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 416.3500 0.0000 416.4500 0.4200 ;
    END
  END p_spm_slave[21]
  PIN p_spm_slave[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 415.3500 0.0000 415.4500 0.4200 ;
    END
  END p_spm_slave[20]
  PIN p_spm_slave[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 414.3500 0.0000 414.4500 0.4200 ;
    END
  END p_spm_slave[19]
  PIN p_spm_slave[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 413.3500 0.0000 413.4500 0.4200 ;
    END
  END p_spm_slave[18]
  PIN p_spm_slave[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 412.3500 0.0000 412.4500 0.4200 ;
    END
  END p_spm_slave[17]
  PIN p_spm_slave[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 411.3500 0.0000 411.4500 0.4200 ;
    END
  END p_spm_slave[16]
  PIN p_spm_slave[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 410.3500 0.0000 410.4500 0.4200 ;
    END
  END p_spm_slave[15]
  PIN p_spm_slave[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 409.3500 0.0000 409.4500 0.4200 ;
    END
  END p_spm_slave[14]
  PIN p_spm_slave[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 408.3500 0.0000 408.4500 0.4200 ;
    END
  END p_spm_slave[13]
  PIN p_spm_slave[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 407.3500 0.0000 407.4500 0.4200 ;
    END
  END p_spm_slave[12]
  PIN p_spm_slave[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 406.3500 0.0000 406.4500 0.4200 ;
    END
  END p_spm_slave[11]
  PIN p_spm_slave[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 405.3500 0.0000 405.4500 0.4200 ;
    END
  END p_spm_slave[10]
  PIN p_spm_slave[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 404.3500 0.0000 404.4500 0.4200 ;
    END
  END p_spm_slave[9]
  PIN p_spm_slave[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 403.3500 0.0000 403.4500 0.4200 ;
    END
  END p_spm_slave[8]
  PIN p_spm_slave[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 402.3500 0.0000 402.4500 0.4200 ;
    END
  END p_spm_slave[7]
  PIN p_spm_slave[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 401.3500 0.0000 401.4500 0.4200 ;
    END
  END p_spm_slave[6]
  PIN p_spm_slave[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 400.3500 0.0000 400.4500 0.4200 ;
    END
  END p_spm_slave[5]
  PIN p_spm_slave[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 399.3500 0.0000 399.4500 0.4200 ;
    END
  END p_spm_slave[4]
  PIN p_spm_slave[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 398.3500 0.0000 398.4500 0.4200 ;
    END
  END p_spm_slave[3]
  PIN p_spm_slave[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 397.3500 0.0000 397.4500 0.4200 ;
    END
  END p_spm_slave[2]
  PIN p_spm_slave[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 396.3500 0.0000 396.4500 0.4200 ;
    END
  END p_spm_slave[1]
  PIN p_spm_slave[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 395.3500 0.0000 395.4500 0.4200 ;
    END
  END p_spm_slave[0]
  PIN p_ocp_master[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.1500 0.0000 72.2500 0.4200 ;
    END
  END p_ocp_master[71]
  PIN p_ocp_master[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.1500 0.0000 71.2500 0.4200 ;
    END
  END p_ocp_master[70]
  PIN p_ocp_master[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.1500 0.0000 70.2500 0.4200 ;
    END
  END p_ocp_master[69]
  PIN p_ocp_master[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.1500 0.0000 69.2500 0.4200 ;
    END
  END p_ocp_master[68]
  PIN p_ocp_master[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.1500 0.0000 68.2500 0.4200 ;
    END
  END p_ocp_master[67]
  PIN p_ocp_master[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.1500 0.0000 67.2500 0.4200 ;
    END
  END p_ocp_master[66]
  PIN p_ocp_master[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.1500 0.0000 66.2500 0.4200 ;
    END
  END p_ocp_master[65]
  PIN p_ocp_master[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.1500 0.0000 65.2500 0.4200 ;
    END
  END p_ocp_master[64]
  PIN p_ocp_master[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.1500 0.0000 64.2500 0.4200 ;
    END
  END p_ocp_master[63]
  PIN p_ocp_master[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.1500 0.0000 63.2500 0.4200 ;
    END
  END p_ocp_master[62]
  PIN p_ocp_master[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.1500 0.0000 62.2500 0.4200 ;
    END
  END p_ocp_master[61]
  PIN p_ocp_master[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.1500 0.0000 61.2500 0.4200 ;
    END
  END p_ocp_master[60]
  PIN p_ocp_master[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.1500 0.0000 60.2500 0.4200 ;
    END
  END p_ocp_master[59]
  PIN p_ocp_master[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.1500 0.0000 59.2500 0.4200 ;
    END
  END p_ocp_master[58]
  PIN p_ocp_master[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.1500 0.0000 58.2500 0.4200 ;
    END
  END p_ocp_master[57]
  PIN p_ocp_master[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.1500 0.0000 57.2500 0.4200 ;
    END
  END p_ocp_master[56]
  PIN p_ocp_master[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.1500 0.0000 56.2500 0.4200 ;
    END
  END p_ocp_master[55]
  PIN p_ocp_master[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.1500 0.0000 55.2500 0.4200 ;
    END
  END p_ocp_master[54]
  PIN p_ocp_master[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.1500 0.0000 54.2500 0.4200 ;
    END
  END p_ocp_master[53]
  PIN p_ocp_master[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.1500 0.0000 53.2500 0.4200 ;
    END
  END p_ocp_master[52]
  PIN p_ocp_master[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.1500 0.0000 52.2500 0.4200 ;
    END
  END p_ocp_master[51]
  PIN p_ocp_master[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.1500 0.0000 51.2500 0.4200 ;
    END
  END p_ocp_master[50]
  PIN p_ocp_master[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.1500 0.0000 50.2500 0.4200 ;
    END
  END p_ocp_master[49]
  PIN p_ocp_master[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.1500 0.0000 49.2500 0.4200 ;
    END
  END p_ocp_master[48]
  PIN p_ocp_master[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.1500 0.0000 48.2500 0.4200 ;
    END
  END p_ocp_master[47]
  PIN p_ocp_master[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.1500 0.0000 47.2500 0.4200 ;
    END
  END p_ocp_master[46]
  PIN p_ocp_master[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.1500 0.0000 46.2500 0.4200 ;
    END
  END p_ocp_master[45]
  PIN p_ocp_master[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.1500 0.0000 45.2500 0.4200 ;
    END
  END p_ocp_master[44]
  PIN p_ocp_master[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.1500 0.0000 44.2500 0.4200 ;
    END
  END p_ocp_master[43]
  PIN p_ocp_master[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.1500 0.0000 43.2500 0.4200 ;
    END
  END p_ocp_master[42]
  PIN p_ocp_master[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.1500 0.0000 42.2500 0.4200 ;
    END
  END p_ocp_master[41]
  PIN p_ocp_master[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.1500 0.0000 41.2500 0.4200 ;
    END
  END p_ocp_master[40]
  PIN p_ocp_master[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.1500 0.0000 40.2500 0.4200 ;
    END
  END p_ocp_master[39]
  PIN p_ocp_master[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.1500 0.0000 39.2500 0.4200 ;
    END
  END p_ocp_master[38]
  PIN p_ocp_master[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.1500 0.0000 38.2500 0.4200 ;
    END
  END p_ocp_master[37]
  PIN p_ocp_master[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.1500 0.0000 37.2500 0.4200 ;
    END
  END p_ocp_master[36]
  PIN p_ocp_master[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.1500 0.0000 36.2500 0.4200 ;
    END
  END p_ocp_master[35]
  PIN p_ocp_master[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.1500 0.0000 35.2500 0.4200 ;
    END
  END p_ocp_master[34]
  PIN p_ocp_master[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.1500 0.0000 34.2500 0.4200 ;
    END
  END p_ocp_master[33]
  PIN p_ocp_master[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.1500 0.0000 33.2500 0.4200 ;
    END
  END p_ocp_master[32]
  PIN p_ocp_master[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.1500 0.0000 32.2500 0.4200 ;
    END
  END p_ocp_master[31]
  PIN p_ocp_master[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.1500 0.0000 31.2500 0.4200 ;
    END
  END p_ocp_master[30]
  PIN p_ocp_master[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.1500 0.0000 30.2500 0.4200 ;
    END
  END p_ocp_master[29]
  PIN p_ocp_master[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.1500 0.0000 29.2500 0.4200 ;
    END
  END p_ocp_master[28]
  PIN p_ocp_master[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.1500 0.0000 28.2500 0.4200 ;
    END
  END p_ocp_master[27]
  PIN p_ocp_master[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.1500 0.0000 27.2500 0.4200 ;
    END
  END p_ocp_master[26]
  PIN p_ocp_master[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.1500 0.0000 26.2500 0.4200 ;
    END
  END p_ocp_master[25]
  PIN p_ocp_master[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.1500 0.0000 25.2500 0.4200 ;
    END
  END p_ocp_master[24]
  PIN p_ocp_master[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.1500 0.0000 24.2500 0.4200 ;
    END
  END p_ocp_master[23]
  PIN p_ocp_master[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.1500 0.0000 23.2500 0.4200 ;
    END
  END p_ocp_master[22]
  PIN p_ocp_master[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.1500 0.0000 22.2500 0.4200 ;
    END
  END p_ocp_master[21]
  PIN p_ocp_master[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.1500 0.0000 21.2500 0.4200 ;
    END
  END p_ocp_master[20]
  PIN p_ocp_master[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.1500 0.0000 20.2500 0.4200 ;
    END
  END p_ocp_master[19]
  PIN p_ocp_master[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.1500 0.0000 19.2500 0.4200 ;
    END
  END p_ocp_master[18]
  PIN p_ocp_master[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.1500 0.0000 18.2500 0.4200 ;
    END
  END p_ocp_master[17]
  PIN p_ocp_master[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.1500 0.0000 17.2500 0.4200 ;
    END
  END p_ocp_master[16]
  PIN p_ocp_master[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.1500 0.0000 16.2500 0.4200 ;
    END
  END p_ocp_master[15]
  PIN p_ocp_master[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.1500 0.0000 15.2500 0.4200 ;
    END
  END p_ocp_master[14]
  PIN p_ocp_master[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.1500 0.0000 14.2500 0.4200 ;
    END
  END p_ocp_master[13]
  PIN p_ocp_master[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.1500 0.0000 13.2500 0.4200 ;
    END
  END p_ocp_master[12]
  PIN p_ocp_master[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.1500 0.0000 12.2500 0.4200 ;
    END
  END p_ocp_master[11]
  PIN p_ocp_master[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.1500 0.0000 11.2500 0.4200 ;
    END
  END p_ocp_master[10]
  PIN p_ocp_master[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.1500 0.0000 10.2500 0.4200 ;
    END
  END p_ocp_master[9]
  PIN p_ocp_master[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.1500 0.0000 9.2500 0.4200 ;
    END
  END p_ocp_master[8]
  PIN p_ocp_master[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.1500 0.0000 8.2500 0.4200 ;
    END
  END p_ocp_master[7]
  PIN p_ocp_master[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7.1500 0.0000 7.2500 0.4200 ;
    END
  END p_ocp_master[6]
  PIN p_ocp_master[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6.1500 0.0000 6.2500 0.4200 ;
    END
  END p_ocp_master[5]
  PIN p_ocp_master[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5.1500 0.0000 5.2500 0.4200 ;
    END
  END p_ocp_master[4]
  PIN p_ocp_master[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4.1500 0.0000 4.2500 0.4200 ;
    END
  END p_ocp_master[3]
  PIN p_ocp_master[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3.1500 0.0000 3.2500 0.4200 ;
    END
  END p_ocp_master[2]
  PIN p_ocp_master[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2.1500 0.0000 2.2500 0.4200 ;
    END
  END p_ocp_master[1]
  PIN p_ocp_master[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.1500 0.0000 1.2500 0.4200 ;
    END
  END p_ocp_master[0]
  PIN p_ocp_slave[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.1500 0.0000 107.2500 0.4200 ;
    END
  END p_ocp_slave[34]
  PIN p_ocp_slave[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.1500 0.0000 106.2500 0.4200 ;
    END
  END p_ocp_slave[33]
  PIN p_ocp_slave[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.1500 0.0000 105.2500 0.4200 ;
    END
  END p_ocp_slave[32]
  PIN p_ocp_slave[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.1500 0.0000 104.2500 0.4200 ;
    END
  END p_ocp_slave[31]
  PIN p_ocp_slave[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.1500 0.0000 103.2500 0.4200 ;
    END
  END p_ocp_slave[30]
  PIN p_ocp_slave[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.1500 0.0000 102.2500 0.4200 ;
    END
  END p_ocp_slave[29]
  PIN p_ocp_slave[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.1500 0.0000 101.2500 0.4200 ;
    END
  END p_ocp_slave[28]
  PIN p_ocp_slave[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.1500 0.0000 100.2500 0.4200 ;
    END
  END p_ocp_slave[27]
  PIN p_ocp_slave[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.1500 0.0000 99.2500 0.4200 ;
    END
  END p_ocp_slave[26]
  PIN p_ocp_slave[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.1500 0.0000 98.2500 0.4200 ;
    END
  END p_ocp_slave[25]
  PIN p_ocp_slave[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.1500 0.0000 97.2500 0.4200 ;
    END
  END p_ocp_slave[24]
  PIN p_ocp_slave[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.1500 0.0000 96.2500 0.4200 ;
    END
  END p_ocp_slave[23]
  PIN p_ocp_slave[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.1500 0.0000 95.2500 0.4200 ;
    END
  END p_ocp_slave[22]
  PIN p_ocp_slave[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.1500 0.0000 94.2500 0.4200 ;
    END
  END p_ocp_slave[21]
  PIN p_ocp_slave[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.1500 0.0000 93.2500 0.4200 ;
    END
  END p_ocp_slave[20]
  PIN p_ocp_slave[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92.1500 0.0000 92.2500 0.4200 ;
    END
  END p_ocp_slave[19]
  PIN p_ocp_slave[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 91.1500 0.0000 91.2500 0.4200 ;
    END
  END p_ocp_slave[18]
  PIN p_ocp_slave[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.1500 0.0000 90.2500 0.4200 ;
    END
  END p_ocp_slave[17]
  PIN p_ocp_slave[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.1500 0.0000 89.2500 0.4200 ;
    END
  END p_ocp_slave[16]
  PIN p_ocp_slave[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.1500 0.0000 88.2500 0.4200 ;
    END
  END p_ocp_slave[15]
  PIN p_ocp_slave[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.1500 0.0000 87.2500 0.4200 ;
    END
  END p_ocp_slave[14]
  PIN p_ocp_slave[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.1500 0.0000 86.2500 0.4200 ;
    END
  END p_ocp_slave[13]
  PIN p_ocp_slave[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.1500 0.0000 85.2500 0.4200 ;
    END
  END p_ocp_slave[12]
  PIN p_ocp_slave[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 84.1500 0.0000 84.2500 0.4200 ;
    END
  END p_ocp_slave[11]
  PIN p_ocp_slave[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.1500 0.0000 83.2500 0.4200 ;
    END
  END p_ocp_slave[10]
  PIN p_ocp_slave[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.1500 0.0000 82.2500 0.4200 ;
    END
  END p_ocp_slave[9]
  PIN p_ocp_slave[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.1500 0.0000 81.2500 0.4200 ;
    END
  END p_ocp_slave[8]
  PIN p_ocp_slave[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.1500 0.0000 80.2500 0.4200 ;
    END
  END p_ocp_slave[7]
  PIN p_ocp_slave[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.1500 0.0000 79.2500 0.4200 ;
    END
  END p_ocp_slave[6]
  PIN p_ocp_slave[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.1500 0.0000 78.2500 0.4200 ;
    END
  END p_ocp_slave[5]
  PIN p_ocp_slave[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.1500 0.0000 77.2500 0.4200 ;
    END
  END p_ocp_slave[4]
  PIN p_ocp_slave[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.1500 0.0000 76.2500 0.4200 ;
    END
  END p_ocp_slave[3]
  PIN p_ocp_slave[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.1500 0.0000 75.2500 0.4200 ;
    END
  END p_ocp_slave[2]
  PIN p_ocp_slave[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.1500 0.0000 74.2500 0.4200 ;
    END
  END p_ocp_slave[1]
  PIN p_ocp_slave[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.1500 0.0000 73.2500 0.4200 ;
    END
  END p_ocp_slave[0]
  PIN p_settings[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.1500 0.0000 115.2500 0.4200 ;
    END
  END p_settings[7]
  PIN p_settings[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.1500 0.0000 114.2500 0.4200 ;
    END
  END p_settings[6]
  PIN p_settings[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 113.1500 0.0000 113.2500 0.4200 ;
    END
  END p_settings[5]
  PIN p_settings[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.1500 0.0000 112.2500 0.4200 ;
    END
  END p_settings[4]
  PIN p_settings[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.1500 0.0000 111.2500 0.4200 ;
    END
  END p_settings[3]
  PIN p_settings[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.1500 0.0000 110.2500 0.4200 ;
    END
  END p_settings[2]
  PIN p_settings[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.1500 0.0000 109.2500 0.4200 ;
    END
  END p_settings[1]
  PIN p_settings[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.1500 0.0000 108.2500 0.4200 ;
    END
  END p_settings[0]
  OBS
    LAYER OVERLAP ;
    LAYER AP ;
      RECT 0.0000 0.0000 1383.2000 1175.2000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 1383.2000 1175.2000 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 1383.2000 1175.2000 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 1383.2000 1175.2000 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 1383.2000 1175.2000 ;
    LAYER M3 ;
      RECT 0.0000 0.0000 1383.2000 1175.2000 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 1383.2000 1175.2000 ;
    LAYER M1 ;
      RECT 0.0000 0.0000 1383.2000 1175.2000 ;
  END
END processor

END LIBRARY
