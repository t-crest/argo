module tdp_ram_14_5
  (input  a_clk,
   input  a_wr,
   input  [4:0] a_addr,
   input  [13:0] a_din,
   input  b_clk,
   input  b_wr,
   input  [4:0] b_addr,
   input  [13:0] b_din,
   output [13:0] a_dout,
   output [13:0] b_dout);
  reg [13:0] n3000_data; // mem_rd
  reg [13:0] n3003_data; // mem_rd
  assign a_dout = n3003_data;
  assign b_dout = n3000_data;
  /* mem/tdp_ram.vhd:57:5  */
  reg [13:0] mem[31:0] ; // memory
  initial begin
    mem[31] = 14'b00000000000000;
    mem[30] = 14'b00000000000000;
    mem[29] = 14'b00000000000000;
    mem[28] = 14'b00000000000000;
    mem[27] = 14'b00000000000000;
    mem[26] = 14'b00000000000000;
    mem[25] = 14'b00000000000000;
    mem[24] = 14'b00000000000000;
    mem[23] = 14'b00000000000000;
    mem[22] = 14'b00000000000000;
    mem[21] = 14'b00000000000000;
    mem[20] = 14'b00000000000000;
    mem[19] = 14'b00000000000000;
    mem[18] = 14'b00000000000000;
    mem[17] = 14'b00000000000000;
    mem[16] = 14'b00000000000000;
    mem[15] = 14'b00000000000000;
    mem[14] = 14'b00000000000000;
    mem[13] = 14'b00000000000000;
    mem[12] = 14'b00000000000000;
    mem[11] = 14'b00000000000000;
    mem[10] = 14'b00000000000000;
    mem[9] = 14'b00000000000000;
    mem[8] = 14'b00000000000000;
    mem[7] = 14'b00000000000000;
    mem[6] = 14'b00000000000000;
    mem[5] = 14'b00000000000000;
    mem[4] = 14'b00000000000000;
    mem[3] = 14'b00000000000000;
    mem[2] = 14'b00000000000000;
    mem[1] = 14'b00000000000000;
    mem[0] = 14'b00000000000000;
    end
  always @(posedge b_clk)
    if (b_wr)
      mem[b_addr] <= b_din;
  always @(posedge b_clk)
    if (1'b1)
      n3000_data <= mem[b_addr];
  always @(posedge a_clk)
    if (a_wr)
      mem[a_addr] <= a_din;
  always @(posedge a_clk)
    if (1'b1)
      n3003_data <= mem[a_addr];
  /* mem/tdp_ram.vhd:104:17  */
  /* mem/tdp_ram.vhd:88:17  */
  /* mem/tdp_ram.vhd:103:9  */
endmodule

module tdp_ram_16_6
  (input  a_clk,
   input  a_wr,
   input  [5:0] a_addr,
   input  [15:0] a_din,
   input  b_clk,
   input  b_wr,
   input  [5:0] b_addr,
   input  [15:0] b_din,
   output [15:0] a_dout,
   output [15:0] b_dout);
  reg [15:0] n2961_data; // mem_rd
  reg [15:0] n2964_data; // mem_rd
  assign a_dout = n2964_data;
  assign b_dout = n2961_data;
  /* mem/tdp_ram.vhd:57:5  */
  reg [15:0] mem[63:0] ; // memory
  initial begin
    mem[63] = 16'b0000000000000000;
    mem[62] = 16'b0000000000000000;
    mem[61] = 16'b0000000000000000;
    mem[60] = 16'b0000000000000000;
    mem[59] = 16'b0000000000000000;
    mem[58] = 16'b0000000000000000;
    mem[57] = 16'b0000000000000000;
    mem[56] = 16'b0000000000000000;
    mem[55] = 16'b0000000000000000;
    mem[54] = 16'b0000000000000000;
    mem[53] = 16'b0000000000000000;
    mem[52] = 16'b0000000000000000;
    mem[51] = 16'b0000000000000000;
    mem[50] = 16'b0000000000000000;
    mem[49] = 16'b0000000000000000;
    mem[48] = 16'b0000000000000000;
    mem[47] = 16'b0000000000000000;
    mem[46] = 16'b0000000000000000;
    mem[45] = 16'b0000000000000000;
    mem[44] = 16'b0000000000000000;
    mem[43] = 16'b0000000000000000;
    mem[42] = 16'b0000000000000000;
    mem[41] = 16'b0000000000000000;
    mem[40] = 16'b0000000000000000;
    mem[39] = 16'b0000000000000000;
    mem[38] = 16'b0000000000000000;
    mem[37] = 16'b0000000000000000;
    mem[36] = 16'b0000000000000000;
    mem[35] = 16'b0000000000000000;
    mem[34] = 16'b0000000000000000;
    mem[33] = 16'b0000000000000000;
    mem[32] = 16'b0000000000000000;
    mem[31] = 16'b0000000000000000;
    mem[30] = 16'b0000000000000000;
    mem[29] = 16'b0000000000000000;
    mem[28] = 16'b0000000000000000;
    mem[27] = 16'b0000000000000000;
    mem[26] = 16'b0000000000000000;
    mem[25] = 16'b0000000000000000;
    mem[24] = 16'b0000000000000000;
    mem[23] = 16'b0000000000000000;
    mem[22] = 16'b0000000000000000;
    mem[21] = 16'b0000000000000000;
    mem[20] = 16'b0000000000000000;
    mem[19] = 16'b0000000000000000;
    mem[18] = 16'b0000000000000000;
    mem[17] = 16'b0000000000000000;
    mem[16] = 16'b0000000000000000;
    mem[15] = 16'b0000000000000000;
    mem[14] = 16'b0000000000000000;
    mem[13] = 16'b0000000000000000;
    mem[12] = 16'b0000000000000000;
    mem[11] = 16'b0000000000000000;
    mem[10] = 16'b0000000000000000;
    mem[9] = 16'b0000000000000000;
    mem[8] = 16'b0000000000000000;
    mem[7] = 16'b0000000000000000;
    mem[6] = 16'b0000000000000000;
    mem[5] = 16'b0000000000000000;
    mem[4] = 16'b0000000000000000;
    mem[3] = 16'b0000000000000000;
    mem[2] = 16'b0000000000000000;
    mem[1] = 16'b0000000000000000;
    mem[0] = 16'b0000000000000000;
    end
  always @(posedge b_clk)
    if (b_wr)
      mem[b_addr] <= b_din;
  always @(posedge b_clk)
    if (1'b1)
      n2961_data <= mem[b_addr];
  always @(posedge a_clk)
    if (a_wr)
      mem[a_addr] <= a_din;
  always @(posedge a_clk)
    if (1'b1)
      n2964_data <= mem[a_addr];
  /* mem/tdp_ram.vhd:104:17  */
  /* mem/tdp_ram.vhd:88:17  */
  /* mem/tdp_ram.vhd:103:9  */
endmodule

module tdp_ram_29_6
  (input  a_clk,
   input  a_wr,
   input  [5:0] a_addr,
   input  [28:0] a_din,
   input  b_clk,
   input  b_wr,
   input  [5:0] b_addr,
   input  [28:0] b_din,
   output [28:0] a_dout,
   output [28:0] b_dout);
  reg [28:0] n2922_data; // mem_rd
  reg [28:0] n2925_data; // mem_rd
  assign a_dout = n2925_data;
  assign b_dout = n2922_data;
  /* mem/tdp_ram.vhd:57:5  */
  reg [28:0] mem[63:0] ; // memory
  initial begin
    mem[63] = 29'b00000000000000000000000000000;
    mem[62] = 29'b00000000000000000000000000000;
    mem[61] = 29'b00000000000000000000000000000;
    mem[60] = 29'b00000000000000000000000000000;
    mem[59] = 29'b00000000000000000000000000000;
    mem[58] = 29'b00000000000000000000000000000;
    mem[57] = 29'b00000000000000000000000000000;
    mem[56] = 29'b00000000000000000000000000000;
    mem[55] = 29'b00000000000000000000000000000;
    mem[54] = 29'b00000000000000000000000000000;
    mem[53] = 29'b00000000000000000000000000000;
    mem[52] = 29'b00000000000000000000000000000;
    mem[51] = 29'b00000000000000000000000000000;
    mem[50] = 29'b00000000000000000000000000000;
    mem[49] = 29'b00000000000000000000000000000;
    mem[48] = 29'b00000000000000000000000000000;
    mem[47] = 29'b00000000000000000000000000000;
    mem[46] = 29'b00000000000000000000000000000;
    mem[45] = 29'b00000000000000000000000000000;
    mem[44] = 29'b00000000000000000000000000000;
    mem[43] = 29'b00000000000000000000000000000;
    mem[42] = 29'b00000000000000000000000000000;
    mem[41] = 29'b00000000000000000000000000000;
    mem[40] = 29'b00000000000000000000000000000;
    mem[39] = 29'b00000000000000000000000000000;
    mem[38] = 29'b00000000000000000000000000000;
    mem[37] = 29'b00000000000000000000000000000;
    mem[36] = 29'b00000000000000000000000000000;
    mem[35] = 29'b00000000000000000000000000000;
    mem[34] = 29'b00000000000000000000000000000;
    mem[33] = 29'b00000000000000000000000000000;
    mem[32] = 29'b00000000000000000000000000000;
    mem[31] = 29'b00000000000000000000000000000;
    mem[30] = 29'b00000000000000000000000000000;
    mem[29] = 29'b00000000000000000000000000000;
    mem[28] = 29'b00000000000000000000000000000;
    mem[27] = 29'b00000000000000000000000000000;
    mem[26] = 29'b00000000000000000000000000000;
    mem[25] = 29'b00000000000000000000000000000;
    mem[24] = 29'b00000000000000000000000000000;
    mem[23] = 29'b00000000000000000000000000000;
    mem[22] = 29'b00000000000000000000000000000;
    mem[21] = 29'b00000000000000000000000000000;
    mem[20] = 29'b00000000000000000000000000000;
    mem[19] = 29'b00000000000000000000000000000;
    mem[18] = 29'b00000000000000000000000000000;
    mem[17] = 29'b00000000000000000000000000000;
    mem[16] = 29'b00000000000000000000000000000;
    mem[15] = 29'b00000000000000000000000000000;
    mem[14] = 29'b00000000000000000000000000000;
    mem[13] = 29'b00000000000000000000000000000;
    mem[12] = 29'b00000000000000000000000000000;
    mem[11] = 29'b00000000000000000000000000000;
    mem[10] = 29'b00000000000000000000000000000;
    mem[9] = 29'b00000000000000000000000000000;
    mem[8] = 29'b00000000000000000000000000000;
    mem[7] = 29'b00000000000000000000000000000;
    mem[6] = 29'b00000000000000000000000000000;
    mem[5] = 29'b00000000000000000000000000000;
    mem[4] = 29'b00000000000000000000000000000;
    mem[3] = 29'b00000000000000000000000000000;
    mem[2] = 29'b00000000000000000000000000000;
    mem[1] = 29'b00000000000000000000000000000;
    mem[0] = 29'b00000000000000000000000000000;
    end
  always @(posedge b_clk)
    if (b_wr)
      mem[b_addr] <= b_din;
  always @(posedge b_clk)
    if (1'b1)
      n2922_data <= mem[b_addr];
  always @(posedge a_clk)
    if (a_wr)
      mem[a_addr] <= a_din;
  always @(posedge a_clk)
    if (1'b1)
      n2925_data <= mem[a_addr];
  /* mem/tdp_ram.vhd:104:17  */
  /* mem/tdp_ram.vhd:88:17  */
  /* mem/tdp_ram.vhd:103:9  */
endmodule

module tdp_ram_30_8
  (input  a_clk,
   input  a_wr,
   input  [7:0] a_addr,
   input  [29:0] a_din,
   input  b_clk,
   input  b_wr,
   input  [7:0] b_addr,
   input  [29:0] b_din,
   output [29:0] a_dout,
   output [29:0] b_dout);
  reg [29:0] n2883_data; // mem_rd
  reg [29:0] n2886_data; // mem_rd
  assign a_dout = n2886_data;
  assign b_dout = n2883_data;
  /* mem/tdp_ram.vhd:57:5  */
  reg [29:0] mem[255:0] ; // memory
  initial begin
    mem[255] = 30'b000000000000000000000000000000;
    mem[254] = 30'b000000000000000000000000000000;
    mem[253] = 30'b000000000000000000000000000000;
    mem[252] = 30'b000000000000000000000000000000;
    mem[251] = 30'b000000000000000000000000000000;
    mem[250] = 30'b000000000000000000000000000000;
    mem[249] = 30'b000000000000000000000000000000;
    mem[248] = 30'b000000000000000000000000000000;
    mem[247] = 30'b000000000000000000000000000000;
    mem[246] = 30'b000000000000000000000000000000;
    mem[245] = 30'b000000000000000000000000000000;
    mem[244] = 30'b000000000000000000000000000000;
    mem[243] = 30'b000000000000000000000000000000;
    mem[242] = 30'b000000000000000000000000000000;
    mem[241] = 30'b000000000000000000000000000000;
    mem[240] = 30'b000000000000000000000000000000;
    mem[239] = 30'b000000000000000000000000000000;
    mem[238] = 30'b000000000000000000000000000000;
    mem[237] = 30'b000000000000000000000000000000;
    mem[236] = 30'b000000000000000000000000000000;
    mem[235] = 30'b000000000000000000000000000000;
    mem[234] = 30'b000000000000000000000000000000;
    mem[233] = 30'b000000000000000000000000000000;
    mem[232] = 30'b000000000000000000000000000000;
    mem[231] = 30'b000000000000000000000000000000;
    mem[230] = 30'b000000000000000000000000000000;
    mem[229] = 30'b000000000000000000000000000000;
    mem[228] = 30'b000000000000000000000000000000;
    mem[227] = 30'b000000000000000000000000000000;
    mem[226] = 30'b000000000000000000000000000000;
    mem[225] = 30'b000000000000000000000000000000;
    mem[224] = 30'b000000000000000000000000000000;
    mem[223] = 30'b000000000000000000000000000000;
    mem[222] = 30'b000000000000000000000000000000;
    mem[221] = 30'b000000000000000000000000000000;
    mem[220] = 30'b000000000000000000000000000000;
    mem[219] = 30'b000000000000000000000000000000;
    mem[218] = 30'b000000000000000000000000000000;
    mem[217] = 30'b000000000000000000000000000000;
    mem[216] = 30'b000000000000000000000000000000;
    mem[215] = 30'b000000000000000000000000000000;
    mem[214] = 30'b000000000000000000000000000000;
    mem[213] = 30'b000000000000000000000000000000;
    mem[212] = 30'b000000000000000000000000000000;
    mem[211] = 30'b000000000000000000000000000000;
    mem[210] = 30'b000000000000000000000000000000;
    mem[209] = 30'b000000000000000000000000000000;
    mem[208] = 30'b000000000000000000000000000000;
    mem[207] = 30'b000000000000000000000000000000;
    mem[206] = 30'b000000000000000000000000000000;
    mem[205] = 30'b000000000000000000000000000000;
    mem[204] = 30'b000000000000000000000000000000;
    mem[203] = 30'b000000000000000000000000000000;
    mem[202] = 30'b000000000000000000000000000000;
    mem[201] = 30'b000000000000000000000000000000;
    mem[200] = 30'b000000000000000000000000000000;
    mem[199] = 30'b000000000000000000000000000000;
    mem[198] = 30'b000000000000000000000000000000;
    mem[197] = 30'b000000000000000000000000000000;
    mem[196] = 30'b000000000000000000000000000000;
    mem[195] = 30'b000000000000000000000000000000;
    mem[194] = 30'b000000000000000000000000000000;
    mem[193] = 30'b000000000000000000000000000000;
    mem[192] = 30'b000000000000000000000000000000;
    mem[191] = 30'b000000000000000000000000000000;
    mem[190] = 30'b000000000000000000000000000000;
    mem[189] = 30'b000000000000000000000000000000;
    mem[188] = 30'b000000000000000000000000000000;
    mem[187] = 30'b000000000000000000000000000000;
    mem[186] = 30'b000000000000000000000000000000;
    mem[185] = 30'b000000000000000000000000000000;
    mem[184] = 30'b000000000000000000000000000000;
    mem[183] = 30'b000000000000000000000000000000;
    mem[182] = 30'b000000000000000000000000000000;
    mem[181] = 30'b000000000000000000000000000000;
    mem[180] = 30'b000000000000000000000000000000;
    mem[179] = 30'b000000000000000000000000000000;
    mem[178] = 30'b000000000000000000000000000000;
    mem[177] = 30'b000000000000000000000000000000;
    mem[176] = 30'b000000000000000000000000000000;
    mem[175] = 30'b000000000000000000000000000000;
    mem[174] = 30'b000000000000000000000000000000;
    mem[173] = 30'b000000000000000000000000000000;
    mem[172] = 30'b000000000000000000000000000000;
    mem[171] = 30'b000000000000000000000000000000;
    mem[170] = 30'b000000000000000000000000000000;
    mem[169] = 30'b000000000000000000000000000000;
    mem[168] = 30'b000000000000000000000000000000;
    mem[167] = 30'b000000000000000000000000000000;
    mem[166] = 30'b000000000000000000000000000000;
    mem[165] = 30'b000000000000000000000000000000;
    mem[164] = 30'b000000000000000000000000000000;
    mem[163] = 30'b000000000000000000000000000000;
    mem[162] = 30'b000000000000000000000000000000;
    mem[161] = 30'b000000000000000000000000000000;
    mem[160] = 30'b000000000000000000000000000000;
    mem[159] = 30'b000000000000000000000000000000;
    mem[158] = 30'b000000000000000000000000000000;
    mem[157] = 30'b000000000000000000000000000000;
    mem[156] = 30'b000000000000000000000000000000;
    mem[155] = 30'b000000000000000000000000000000;
    mem[154] = 30'b000000000000000000000000000000;
    mem[153] = 30'b000000000000000000000000000000;
    mem[152] = 30'b000000000000000000000000000000;
    mem[151] = 30'b000000000000000000000000000000;
    mem[150] = 30'b000000000000000000000000000000;
    mem[149] = 30'b000000000000000000000000000000;
    mem[148] = 30'b000000000000000000000000000000;
    mem[147] = 30'b000000000000000000000000000000;
    mem[146] = 30'b000000000000000000000000000000;
    mem[145] = 30'b000000000000000000000000000000;
    mem[144] = 30'b000000000000000000000000000000;
    mem[143] = 30'b000000000000000000000000000000;
    mem[142] = 30'b000000000000000000000000000000;
    mem[141] = 30'b000000000000000000000000000000;
    mem[140] = 30'b000000000000000000000000000000;
    mem[139] = 30'b000000000000000000000000000000;
    mem[138] = 30'b000000000000000000000000000000;
    mem[137] = 30'b000000000000000000000000000000;
    mem[136] = 30'b000000000000000000000000000000;
    mem[135] = 30'b000000000000000000000000000000;
    mem[134] = 30'b000000000000000000000000000000;
    mem[133] = 30'b000000000000000000000000000000;
    mem[132] = 30'b000000000000000000000000000000;
    mem[131] = 30'b000000000000000000000000000000;
    mem[130] = 30'b000000000000000000000000000000;
    mem[129] = 30'b000000000000000000000000000000;
    mem[128] = 30'b000000000000000000000000000000;
    mem[127] = 30'b000000000000000000000000000000;
    mem[126] = 30'b000000000000000000000000000000;
    mem[125] = 30'b000000000000000000000000000000;
    mem[124] = 30'b000000000000000000000000000000;
    mem[123] = 30'b000000000000000000000000000000;
    mem[122] = 30'b000000000000000000000000000000;
    mem[121] = 30'b000000000000000000000000000000;
    mem[120] = 30'b000000000000000000000000000000;
    mem[119] = 30'b000000000000000000000000000000;
    mem[118] = 30'b000000000000000000000000000000;
    mem[117] = 30'b000000000000000000000000000000;
    mem[116] = 30'b000000000000000000000000000000;
    mem[115] = 30'b000000000000000000000000000000;
    mem[114] = 30'b000000000000000000000000000000;
    mem[113] = 30'b000000000000000000000000000000;
    mem[112] = 30'b000000000000000000000000000000;
    mem[111] = 30'b000000000000000000000000000000;
    mem[110] = 30'b000000000000000000000000000000;
    mem[109] = 30'b000000000000000000000000000000;
    mem[108] = 30'b000000000000000000000000000000;
    mem[107] = 30'b000000000000000000000000000000;
    mem[106] = 30'b000000000000000000000000000000;
    mem[105] = 30'b000000000000000000000000000000;
    mem[104] = 30'b000000000000000000000000000000;
    mem[103] = 30'b000000000000000000000000000000;
    mem[102] = 30'b000000000000000000000000000000;
    mem[101] = 30'b000000000000000000000000000000;
    mem[100] = 30'b000000000000000000000000000000;
    mem[99] = 30'b000000000000000000000000000000;
    mem[98] = 30'b000000000000000000000000000000;
    mem[97] = 30'b000000000000000000000000000000;
    mem[96] = 30'b000000000000000000000000000000;
    mem[95] = 30'b000000000000000000000000000000;
    mem[94] = 30'b000000000000000000000000000000;
    mem[93] = 30'b000000000000000000000000000000;
    mem[92] = 30'b000000000000000000000000000000;
    mem[91] = 30'b000000000000000000000000000000;
    mem[90] = 30'b000000000000000000000000000000;
    mem[89] = 30'b000000000000000000000000000000;
    mem[88] = 30'b000000000000000000000000000000;
    mem[87] = 30'b000000000000000000000000000000;
    mem[86] = 30'b000000000000000000000000000000;
    mem[85] = 30'b000000000000000000000000000000;
    mem[84] = 30'b000000000000000000000000000000;
    mem[83] = 30'b000000000000000000000000000000;
    mem[82] = 30'b000000000000000000000000000000;
    mem[81] = 30'b000000000000000000000000000000;
    mem[80] = 30'b000000000000000000000000000000;
    mem[79] = 30'b000000000000000000000000000000;
    mem[78] = 30'b000000000000000000000000000000;
    mem[77] = 30'b000000000000000000000000000000;
    mem[76] = 30'b000000000000000000000000000000;
    mem[75] = 30'b000000000000000000000000000000;
    mem[74] = 30'b000000000000000000000000000000;
    mem[73] = 30'b000000000000000000000000000000;
    mem[72] = 30'b000000000000000000000000000000;
    mem[71] = 30'b000000000000000000000000000000;
    mem[70] = 30'b000000000000000000000000000000;
    mem[69] = 30'b000000000000000000000000000000;
    mem[68] = 30'b000000000000000000000000000000;
    mem[67] = 30'b000000000000000000000000000000;
    mem[66] = 30'b000000000000000000000000000000;
    mem[65] = 30'b000000000000000000000000000000;
    mem[64] = 30'b000000000000000000000000000000;
    mem[63] = 30'b000000000000000000000000000000;
    mem[62] = 30'b000000000000000000000000000000;
    mem[61] = 30'b000000000000000000000000000000;
    mem[60] = 30'b000000000000000000000000000000;
    mem[59] = 30'b000000000000000000000000000000;
    mem[58] = 30'b000000000000000000000000000000;
    mem[57] = 30'b000000000000000000000000000000;
    mem[56] = 30'b000000000000000000000000000000;
    mem[55] = 30'b000000000000000000000000000000;
    mem[54] = 30'b000000000000000000000000000000;
    mem[53] = 30'b000000000000000000000000000000;
    mem[52] = 30'b000000000000000000000000000000;
    mem[51] = 30'b000000000000000000000000000000;
    mem[50] = 30'b000000000000000000000000000000;
    mem[49] = 30'b000000000000000000000000000000;
    mem[48] = 30'b000000000000000000000000000000;
    mem[47] = 30'b000000000000000000000000000000;
    mem[46] = 30'b000000000000000000000000000000;
    mem[45] = 30'b000000000000000000000000000000;
    mem[44] = 30'b000000000000000000000000000000;
    mem[43] = 30'b000000000000000000000000000000;
    mem[42] = 30'b000000000000000000000000000000;
    mem[41] = 30'b000000000000000000000000000000;
    mem[40] = 30'b000000000000000000000000000000;
    mem[39] = 30'b000000000000000000000000000000;
    mem[38] = 30'b000000000000000000000000000000;
    mem[37] = 30'b000000000000000000000000000000;
    mem[36] = 30'b000000000000000000000000000000;
    mem[35] = 30'b000000000000000000000000000000;
    mem[34] = 30'b000000000000000000000000000000;
    mem[33] = 30'b000000000000000000000000000000;
    mem[32] = 30'b000000000000000000000000000000;
    mem[31] = 30'b000000000000000000000000000000;
    mem[30] = 30'b000000000000000000000000000000;
    mem[29] = 30'b000000000000000000000000000000;
    mem[28] = 30'b000000000000000000000000000000;
    mem[27] = 30'b000000000000000000000000000000;
    mem[26] = 30'b000000000000000000000000000000;
    mem[25] = 30'b000000000000000000000000000000;
    mem[24] = 30'b000000000000000000000000000000;
    mem[23] = 30'b000000000000000000000000000000;
    mem[22] = 30'b000000000000000000000000000000;
    mem[21] = 30'b000000000000000000000000000000;
    mem[20] = 30'b000000000000000000000000000000;
    mem[19] = 30'b000000000000000000000000000000;
    mem[18] = 30'b000000000000000000000000000000;
    mem[17] = 30'b000000000000000000000000000000;
    mem[16] = 30'b000000000000000000000000000000;
    mem[15] = 30'b000000000000000000000000000000;
    mem[14] = 30'b000000000000000000000000000000;
    mem[13] = 30'b000000000000000000000000000000;
    mem[12] = 30'b000000000000000000000000000000;
    mem[11] = 30'b000000000000000000000000000000;
    mem[10] = 30'b000000000000000000000000000000;
    mem[9] = 30'b000000000000000000000000000000;
    mem[8] = 30'b000000000000000000000000000000;
    mem[7] = 30'b000000000000000000000000000000;
    mem[6] = 30'b000000000000000000000000000000;
    mem[5] = 30'b000000000000000000000000000000;
    mem[4] = 30'b000000000000000000000000000000;
    mem[3] = 30'b000000000000000000000000000000;
    mem[2] = 30'b000000000000000000000000000000;
    mem[1] = 30'b000000000000000000000000000000;
    mem[0] = 30'b000000000000000000000000000000;
    end
  always @(posedge b_clk)
    if (b_wr)
      mem[b_addr] <= b_din;
  always @(posedge b_clk)
    if (1'b1)
      n2883_data <= mem[b_addr];
  always @(posedge a_clk)
    if (a_wr)
      mem[a_addr] <= a_din;
  always @(posedge a_clk)
    if (1'b1)
      n2886_data <= mem[a_addr];
  /* mem/tdp_ram.vhd:104:17  */
  /* mem/tdp_ram.vhd:88:17  */
  /* mem/tdp_ram.vhd:103:9  */
endmodule

module xbar
  (input  [19:0] func,
   input  [179:0] inport,
   output [179:0] outport);
  wire [3:0] sel0;
  wire [3:0] sel1;
  wire [3:0] sel2;
  wire [3:0] sel3;
  wire [3:0] sel4;
  wire [3:0] n1822_o;
  wire [3:0] n1823_o;
  wire [3:0] n1824_o;
  wire [3:0] n1825_o;
  wire [3:0] n1826_o;
  wire [35:0] n1827_o;
  wire [34:0] n1828_o;
  wire n1829_o;
  wire n1830_o;
  wire n1831_o;
  wire n1832_o;
  wire n1833_o;
  wire n1834_o;
  wire n1835_o;
  wire n1836_o;
  wire n1837_o;
  wire n1838_o;
  wire n1839_o;
  wire n1840_o;
  wire n1841_o;
  wire n1842_o;
  wire n1843_o;
  wire n1844_o;
  wire n1845_o;
  wire n1846_o;
  wire n1847_o;
  wire n1848_o;
  wire n1849_o;
  wire n1850_o;
  wire n1851_o;
  wire n1852_o;
  wire n1853_o;
  wire n1854_o;
  wire n1855_o;
  wire n1856_o;
  wire n1857_o;
  wire n1858_o;
  wire n1859_o;
  wire n1860_o;
  wire n1861_o;
  wire n1862_o;
  wire n1863_o;
  wire [3:0] n1864_o;
  wire [3:0] n1865_o;
  wire [3:0] n1866_o;
  wire [3:0] n1867_o;
  wire [3:0] n1868_o;
  wire [3:0] n1869_o;
  wire [3:0] n1870_o;
  wire [3:0] n1871_o;
  wire [2:0] n1872_o;
  wire [15:0] n1873_o;
  wire [15:0] n1874_o;
  wire [34:0] n1875_o;
  wire [34:0] n1876_o;
  wire [35:0] n1877_o;
  wire [34:0] n1878_o;
  wire n1879_o;
  wire n1880_o;
  wire n1881_o;
  wire n1882_o;
  wire n1883_o;
  wire n1884_o;
  wire n1885_o;
  wire n1886_o;
  wire n1887_o;
  wire n1888_o;
  wire n1889_o;
  wire n1890_o;
  wire n1891_o;
  wire n1892_o;
  wire n1893_o;
  wire n1894_o;
  wire n1895_o;
  wire n1896_o;
  wire n1897_o;
  wire n1898_o;
  wire n1899_o;
  wire n1900_o;
  wire n1901_o;
  wire n1902_o;
  wire n1903_o;
  wire n1904_o;
  wire n1905_o;
  wire n1906_o;
  wire n1907_o;
  wire n1908_o;
  wire n1909_o;
  wire n1910_o;
  wire n1911_o;
  wire n1912_o;
  wire n1913_o;
  wire [3:0] n1914_o;
  wire [3:0] n1915_o;
  wire [3:0] n1916_o;
  wire [3:0] n1917_o;
  wire [3:0] n1918_o;
  wire [3:0] n1919_o;
  wire [3:0] n1920_o;
  wire [3:0] n1921_o;
  wire [2:0] n1922_o;
  wire [15:0] n1923_o;
  wire [15:0] n1924_o;
  wire [34:0] n1925_o;
  wire [34:0] n1926_o;
  wire [34:0] n1927_o;
  wire [35:0] n1928_o;
  wire [34:0] n1929_o;
  wire n1930_o;
  wire n1931_o;
  wire n1932_o;
  wire n1933_o;
  wire n1934_o;
  wire n1935_o;
  wire n1936_o;
  wire n1937_o;
  wire n1938_o;
  wire n1939_o;
  wire n1940_o;
  wire n1941_o;
  wire n1942_o;
  wire n1943_o;
  wire n1944_o;
  wire n1945_o;
  wire n1946_o;
  wire n1947_o;
  wire n1948_o;
  wire n1949_o;
  wire n1950_o;
  wire n1951_o;
  wire n1952_o;
  wire n1953_o;
  wire n1954_o;
  wire n1955_o;
  wire n1956_o;
  wire n1957_o;
  wire n1958_o;
  wire n1959_o;
  wire n1960_o;
  wire n1961_o;
  wire n1962_o;
  wire n1963_o;
  wire n1964_o;
  wire [3:0] n1965_o;
  wire [3:0] n1966_o;
  wire [3:0] n1967_o;
  wire [3:0] n1968_o;
  wire [3:0] n1969_o;
  wire [3:0] n1970_o;
  wire [3:0] n1971_o;
  wire [3:0] n1972_o;
  wire [2:0] n1973_o;
  wire [15:0] n1974_o;
  wire [15:0] n1975_o;
  wire [34:0] n1976_o;
  wire [34:0] n1977_o;
  wire [34:0] n1978_o;
  wire [35:0] n1979_o;
  wire [34:0] n1980_o;
  wire n1981_o;
  wire n1982_o;
  wire n1983_o;
  wire n1984_o;
  wire n1985_o;
  wire n1986_o;
  wire n1987_o;
  wire n1988_o;
  wire n1989_o;
  wire n1990_o;
  wire n1991_o;
  wire n1992_o;
  wire n1993_o;
  wire n1994_o;
  wire n1995_o;
  wire n1996_o;
  wire n1997_o;
  wire n1998_o;
  wire n1999_o;
  wire n2000_o;
  wire n2001_o;
  wire n2002_o;
  wire n2003_o;
  wire n2004_o;
  wire n2005_o;
  wire n2006_o;
  wire n2007_o;
  wire n2008_o;
  wire n2009_o;
  wire n2010_o;
  wire n2011_o;
  wire n2012_o;
  wire n2013_o;
  wire n2014_o;
  wire n2015_o;
  wire [3:0] n2016_o;
  wire [3:0] n2017_o;
  wire [3:0] n2018_o;
  wire [3:0] n2019_o;
  wire [3:0] n2020_o;
  wire [3:0] n2021_o;
  wire [3:0] n2022_o;
  wire [3:0] n2023_o;
  wire [2:0] n2024_o;
  wire [15:0] n2025_o;
  wire [15:0] n2026_o;
  wire [34:0] n2027_o;
  wire [34:0] n2028_o;
  wire [34:0] n2029_o;
  wire [35:0] n2030_o;
  wire [34:0] n2031_o;
  wire n2032_o;
  wire n2033_o;
  wire n2034_o;
  wire n2035_o;
  wire n2036_o;
  wire n2037_o;
  wire n2038_o;
  wire n2039_o;
  wire n2040_o;
  wire n2041_o;
  wire n2042_o;
  wire n2043_o;
  wire n2044_o;
  wire n2045_o;
  wire n2046_o;
  wire n2047_o;
  wire n2048_o;
  wire n2049_o;
  wire n2050_o;
  wire n2051_o;
  wire n2052_o;
  wire n2053_o;
  wire n2054_o;
  wire n2055_o;
  wire n2056_o;
  wire n2057_o;
  wire n2058_o;
  wire n2059_o;
  wire n2060_o;
  wire n2061_o;
  wire n2062_o;
  wire n2063_o;
  wire n2064_o;
  wire n2065_o;
  wire n2066_o;
  wire [3:0] n2067_o;
  wire [3:0] n2068_o;
  wire [3:0] n2069_o;
  wire [3:0] n2070_o;
  wire [3:0] n2071_o;
  wire [3:0] n2072_o;
  wire [3:0] n2073_o;
  wire [3:0] n2074_o;
  wire [2:0] n2075_o;
  wire [15:0] n2076_o;
  wire [15:0] n2077_o;
  wire [34:0] n2078_o;
  wire [34:0] n2079_o;
  wire [35:0] n2080_o;
  wire [34:0] n2081_o;
  wire n2082_o;
  wire n2083_o;
  wire n2084_o;
  wire n2085_o;
  wire n2086_o;
  wire n2087_o;
  wire n2088_o;
  wire n2089_o;
  wire n2090_o;
  wire n2091_o;
  wire n2092_o;
  wire n2093_o;
  wire n2094_o;
  wire n2095_o;
  wire n2096_o;
  wire n2097_o;
  wire n2098_o;
  wire n2099_o;
  wire n2100_o;
  wire n2101_o;
  wire n2102_o;
  wire n2103_o;
  wire n2104_o;
  wire n2105_o;
  wire n2106_o;
  wire n2107_o;
  wire n2108_o;
  wire n2109_o;
  wire n2110_o;
  wire n2111_o;
  wire n2112_o;
  wire n2113_o;
  wire n2114_o;
  wire n2115_o;
  wire n2116_o;
  wire [3:0] n2117_o;
  wire [3:0] n2118_o;
  wire [3:0] n2119_o;
  wire [3:0] n2120_o;
  wire [3:0] n2121_o;
  wire [3:0] n2122_o;
  wire [3:0] n2123_o;
  wire [3:0] n2124_o;
  wire [2:0] n2125_o;
  wire [15:0] n2126_o;
  wire [15:0] n2127_o;
  wire [34:0] n2128_o;
  wire [34:0] n2129_o;
  wire [34:0] n2130_o;
  wire [35:0] n2131_o;
  wire [34:0] n2132_o;
  wire n2133_o;
  wire n2134_o;
  wire n2135_o;
  wire n2136_o;
  wire n2137_o;
  wire n2138_o;
  wire n2139_o;
  wire n2140_o;
  wire n2141_o;
  wire n2142_o;
  wire n2143_o;
  wire n2144_o;
  wire n2145_o;
  wire n2146_o;
  wire n2147_o;
  wire n2148_o;
  wire n2149_o;
  wire n2150_o;
  wire n2151_o;
  wire n2152_o;
  wire n2153_o;
  wire n2154_o;
  wire n2155_o;
  wire n2156_o;
  wire n2157_o;
  wire n2158_o;
  wire n2159_o;
  wire n2160_o;
  wire n2161_o;
  wire n2162_o;
  wire n2163_o;
  wire n2164_o;
  wire n2165_o;
  wire n2166_o;
  wire n2167_o;
  wire [3:0] n2168_o;
  wire [3:0] n2169_o;
  wire [3:0] n2170_o;
  wire [3:0] n2171_o;
  wire [3:0] n2172_o;
  wire [3:0] n2173_o;
  wire [3:0] n2174_o;
  wire [3:0] n2175_o;
  wire [2:0] n2176_o;
  wire [15:0] n2177_o;
  wire [15:0] n2178_o;
  wire [34:0] n2179_o;
  wire [34:0] n2180_o;
  wire [34:0] n2181_o;
  wire [35:0] n2182_o;
  wire [34:0] n2183_o;
  wire n2184_o;
  wire n2185_o;
  wire n2186_o;
  wire n2187_o;
  wire n2188_o;
  wire n2189_o;
  wire n2190_o;
  wire n2191_o;
  wire n2192_o;
  wire n2193_o;
  wire n2194_o;
  wire n2195_o;
  wire n2196_o;
  wire n2197_o;
  wire n2198_o;
  wire n2199_o;
  wire n2200_o;
  wire n2201_o;
  wire n2202_o;
  wire n2203_o;
  wire n2204_o;
  wire n2205_o;
  wire n2206_o;
  wire n2207_o;
  wire n2208_o;
  wire n2209_o;
  wire n2210_o;
  wire n2211_o;
  wire n2212_o;
  wire n2213_o;
  wire n2214_o;
  wire n2215_o;
  wire n2216_o;
  wire n2217_o;
  wire n2218_o;
  wire [3:0] n2219_o;
  wire [3:0] n2220_o;
  wire [3:0] n2221_o;
  wire [3:0] n2222_o;
  wire [3:0] n2223_o;
  wire [3:0] n2224_o;
  wire [3:0] n2225_o;
  wire [3:0] n2226_o;
  wire [2:0] n2227_o;
  wire [15:0] n2228_o;
  wire [15:0] n2229_o;
  wire [34:0] n2230_o;
  wire [34:0] n2231_o;
  wire [34:0] n2232_o;
  wire [35:0] n2233_o;
  wire [34:0] n2234_o;
  wire n2235_o;
  wire n2236_o;
  wire n2237_o;
  wire n2238_o;
  wire n2239_o;
  wire n2240_o;
  wire n2241_o;
  wire n2242_o;
  wire n2243_o;
  wire n2244_o;
  wire n2245_o;
  wire n2246_o;
  wire n2247_o;
  wire n2248_o;
  wire n2249_o;
  wire n2250_o;
  wire n2251_o;
  wire n2252_o;
  wire n2253_o;
  wire n2254_o;
  wire n2255_o;
  wire n2256_o;
  wire n2257_o;
  wire n2258_o;
  wire n2259_o;
  wire n2260_o;
  wire n2261_o;
  wire n2262_o;
  wire n2263_o;
  wire n2264_o;
  wire n2265_o;
  wire n2266_o;
  wire n2267_o;
  wire n2268_o;
  wire n2269_o;
  wire [3:0] n2270_o;
  wire [3:0] n2271_o;
  wire [3:0] n2272_o;
  wire [3:0] n2273_o;
  wire [3:0] n2274_o;
  wire [3:0] n2275_o;
  wire [3:0] n2276_o;
  wire [3:0] n2277_o;
  wire [2:0] n2278_o;
  wire [15:0] n2279_o;
  wire [15:0] n2280_o;
  wire [34:0] n2281_o;
  wire [34:0] n2282_o;
  wire [35:0] n2283_o;
  wire [34:0] n2284_o;
  wire n2285_o;
  wire n2286_o;
  wire n2287_o;
  wire n2288_o;
  wire n2289_o;
  wire n2290_o;
  wire n2291_o;
  wire n2292_o;
  wire n2293_o;
  wire n2294_o;
  wire n2295_o;
  wire n2296_o;
  wire n2297_o;
  wire n2298_o;
  wire n2299_o;
  wire n2300_o;
  wire n2301_o;
  wire n2302_o;
  wire n2303_o;
  wire n2304_o;
  wire n2305_o;
  wire n2306_o;
  wire n2307_o;
  wire n2308_o;
  wire n2309_o;
  wire n2310_o;
  wire n2311_o;
  wire n2312_o;
  wire n2313_o;
  wire n2314_o;
  wire n2315_o;
  wire n2316_o;
  wire n2317_o;
  wire n2318_o;
  wire n2319_o;
  wire [3:0] n2320_o;
  wire [3:0] n2321_o;
  wire [3:0] n2322_o;
  wire [3:0] n2323_o;
  wire [3:0] n2324_o;
  wire [3:0] n2325_o;
  wire [3:0] n2326_o;
  wire [3:0] n2327_o;
  wire [2:0] n2328_o;
  wire [15:0] n2329_o;
  wire [15:0] n2330_o;
  wire [34:0] n2331_o;
  wire [34:0] n2332_o;
  wire [34:0] n2333_o;
  wire [35:0] n2334_o;
  wire [34:0] n2335_o;
  wire n2336_o;
  wire n2337_o;
  wire n2338_o;
  wire n2339_o;
  wire n2340_o;
  wire n2341_o;
  wire n2342_o;
  wire n2343_o;
  wire n2344_o;
  wire n2345_o;
  wire n2346_o;
  wire n2347_o;
  wire n2348_o;
  wire n2349_o;
  wire n2350_o;
  wire n2351_o;
  wire n2352_o;
  wire n2353_o;
  wire n2354_o;
  wire n2355_o;
  wire n2356_o;
  wire n2357_o;
  wire n2358_o;
  wire n2359_o;
  wire n2360_o;
  wire n2361_o;
  wire n2362_o;
  wire n2363_o;
  wire n2364_o;
  wire n2365_o;
  wire n2366_o;
  wire n2367_o;
  wire n2368_o;
  wire n2369_o;
  wire n2370_o;
  wire [3:0] n2371_o;
  wire [3:0] n2372_o;
  wire [3:0] n2373_o;
  wire [3:0] n2374_o;
  wire [3:0] n2375_o;
  wire [3:0] n2376_o;
  wire [3:0] n2377_o;
  wire [3:0] n2378_o;
  wire [2:0] n2379_o;
  wire [15:0] n2380_o;
  wire [15:0] n2381_o;
  wire [34:0] n2382_o;
  wire [34:0] n2383_o;
  wire [34:0] n2384_o;
  wire [35:0] n2385_o;
  wire [34:0] n2386_o;
  wire n2387_o;
  wire n2388_o;
  wire n2389_o;
  wire n2390_o;
  wire n2391_o;
  wire n2392_o;
  wire n2393_o;
  wire n2394_o;
  wire n2395_o;
  wire n2396_o;
  wire n2397_o;
  wire n2398_o;
  wire n2399_o;
  wire n2400_o;
  wire n2401_o;
  wire n2402_o;
  wire n2403_o;
  wire n2404_o;
  wire n2405_o;
  wire n2406_o;
  wire n2407_o;
  wire n2408_o;
  wire n2409_o;
  wire n2410_o;
  wire n2411_o;
  wire n2412_o;
  wire n2413_o;
  wire n2414_o;
  wire n2415_o;
  wire n2416_o;
  wire n2417_o;
  wire n2418_o;
  wire n2419_o;
  wire n2420_o;
  wire n2421_o;
  wire [3:0] n2422_o;
  wire [3:0] n2423_o;
  wire [3:0] n2424_o;
  wire [3:0] n2425_o;
  wire [3:0] n2426_o;
  wire [3:0] n2427_o;
  wire [3:0] n2428_o;
  wire [3:0] n2429_o;
  wire [2:0] n2430_o;
  wire [15:0] n2431_o;
  wire [15:0] n2432_o;
  wire [34:0] n2433_o;
  wire [34:0] n2434_o;
  wire [34:0] n2435_o;
  wire [35:0] n2436_o;
  wire [34:0] n2437_o;
  wire n2438_o;
  wire n2439_o;
  wire n2440_o;
  wire n2441_o;
  wire n2442_o;
  wire n2443_o;
  wire n2444_o;
  wire n2445_o;
  wire n2446_o;
  wire n2447_o;
  wire n2448_o;
  wire n2449_o;
  wire n2450_o;
  wire n2451_o;
  wire n2452_o;
  wire n2453_o;
  wire n2454_o;
  wire n2455_o;
  wire n2456_o;
  wire n2457_o;
  wire n2458_o;
  wire n2459_o;
  wire n2460_o;
  wire n2461_o;
  wire n2462_o;
  wire n2463_o;
  wire n2464_o;
  wire n2465_o;
  wire n2466_o;
  wire n2467_o;
  wire n2468_o;
  wire n2469_o;
  wire n2470_o;
  wire n2471_o;
  wire n2472_o;
  wire [3:0] n2473_o;
  wire [3:0] n2474_o;
  wire [3:0] n2475_o;
  wire [3:0] n2476_o;
  wire [3:0] n2477_o;
  wire [3:0] n2478_o;
  wire [3:0] n2479_o;
  wire [3:0] n2480_o;
  wire [2:0] n2481_o;
  wire [15:0] n2482_o;
  wire [15:0] n2483_o;
  wire [34:0] n2484_o;
  wire [34:0] n2485_o;
  wire [35:0] n2486_o;
  wire [34:0] n2487_o;
  wire n2488_o;
  wire n2489_o;
  wire n2490_o;
  wire n2491_o;
  wire n2492_o;
  wire n2493_o;
  wire n2494_o;
  wire n2495_o;
  wire n2496_o;
  wire n2497_o;
  wire n2498_o;
  wire n2499_o;
  wire n2500_o;
  wire n2501_o;
  wire n2502_o;
  wire n2503_o;
  wire n2504_o;
  wire n2505_o;
  wire n2506_o;
  wire n2507_o;
  wire n2508_o;
  wire n2509_o;
  wire n2510_o;
  wire n2511_o;
  wire n2512_o;
  wire n2513_o;
  wire n2514_o;
  wire n2515_o;
  wire n2516_o;
  wire n2517_o;
  wire n2518_o;
  wire n2519_o;
  wire n2520_o;
  wire n2521_o;
  wire n2522_o;
  wire [3:0] n2523_o;
  wire [3:0] n2524_o;
  wire [3:0] n2525_o;
  wire [3:0] n2526_o;
  wire [3:0] n2527_o;
  wire [3:0] n2528_o;
  wire [3:0] n2529_o;
  wire [3:0] n2530_o;
  wire [2:0] n2531_o;
  wire [15:0] n2532_o;
  wire [15:0] n2533_o;
  wire [34:0] n2534_o;
  wire [34:0] n2535_o;
  wire [34:0] n2536_o;
  wire [35:0] n2537_o;
  wire [34:0] n2538_o;
  wire n2539_o;
  wire n2540_o;
  wire n2541_o;
  wire n2542_o;
  wire n2543_o;
  wire n2544_o;
  wire n2545_o;
  wire n2546_o;
  wire n2547_o;
  wire n2548_o;
  wire n2549_o;
  wire n2550_o;
  wire n2551_o;
  wire n2552_o;
  wire n2553_o;
  wire n2554_o;
  wire n2555_o;
  wire n2556_o;
  wire n2557_o;
  wire n2558_o;
  wire n2559_o;
  wire n2560_o;
  wire n2561_o;
  wire n2562_o;
  wire n2563_o;
  wire n2564_o;
  wire n2565_o;
  wire n2566_o;
  wire n2567_o;
  wire n2568_o;
  wire n2569_o;
  wire n2570_o;
  wire n2571_o;
  wire n2572_o;
  wire n2573_o;
  wire [3:0] n2574_o;
  wire [3:0] n2575_o;
  wire [3:0] n2576_o;
  wire [3:0] n2577_o;
  wire [3:0] n2578_o;
  wire [3:0] n2579_o;
  wire [3:0] n2580_o;
  wire [3:0] n2581_o;
  wire [2:0] n2582_o;
  wire [15:0] n2583_o;
  wire [15:0] n2584_o;
  wire [34:0] n2585_o;
  wire [34:0] n2586_o;
  wire [34:0] n2587_o;
  wire [35:0] n2588_o;
  wire [34:0] n2589_o;
  wire n2590_o;
  wire n2591_o;
  wire n2592_o;
  wire n2593_o;
  wire n2594_o;
  wire n2595_o;
  wire n2596_o;
  wire n2597_o;
  wire n2598_o;
  wire n2599_o;
  wire n2600_o;
  wire n2601_o;
  wire n2602_o;
  wire n2603_o;
  wire n2604_o;
  wire n2605_o;
  wire n2606_o;
  wire n2607_o;
  wire n2608_o;
  wire n2609_o;
  wire n2610_o;
  wire n2611_o;
  wire n2612_o;
  wire n2613_o;
  wire n2614_o;
  wire n2615_o;
  wire n2616_o;
  wire n2617_o;
  wire n2618_o;
  wire n2619_o;
  wire n2620_o;
  wire n2621_o;
  wire n2622_o;
  wire n2623_o;
  wire n2624_o;
  wire [3:0] n2625_o;
  wire [3:0] n2626_o;
  wire [3:0] n2627_o;
  wire [3:0] n2628_o;
  wire [3:0] n2629_o;
  wire [3:0] n2630_o;
  wire [3:0] n2631_o;
  wire [3:0] n2632_o;
  wire [2:0] n2633_o;
  wire [15:0] n2634_o;
  wire [15:0] n2635_o;
  wire [34:0] n2636_o;
  wire [34:0] n2637_o;
  wire [34:0] n2638_o;
  wire [35:0] n2639_o;
  wire [34:0] n2640_o;
  wire n2641_o;
  wire n2642_o;
  wire n2643_o;
  wire n2644_o;
  wire n2645_o;
  wire n2646_o;
  wire n2647_o;
  wire n2648_o;
  wire n2649_o;
  wire n2650_o;
  wire n2651_o;
  wire n2652_o;
  wire n2653_o;
  wire n2654_o;
  wire n2655_o;
  wire n2656_o;
  wire n2657_o;
  wire n2658_o;
  wire n2659_o;
  wire n2660_o;
  wire n2661_o;
  wire n2662_o;
  wire n2663_o;
  wire n2664_o;
  wire n2665_o;
  wire n2666_o;
  wire n2667_o;
  wire n2668_o;
  wire n2669_o;
  wire n2670_o;
  wire n2671_o;
  wire n2672_o;
  wire n2673_o;
  wire n2674_o;
  wire n2675_o;
  wire [3:0] n2676_o;
  wire [3:0] n2677_o;
  wire [3:0] n2678_o;
  wire [3:0] n2679_o;
  wire [3:0] n2680_o;
  wire [3:0] n2681_o;
  wire [3:0] n2682_o;
  wire [3:0] n2683_o;
  wire [2:0] n2684_o;
  wire [15:0] n2685_o;
  wire [15:0] n2686_o;
  wire [34:0] n2687_o;
  wire [34:0] n2688_o;
  wire [35:0] n2689_o;
  wire [34:0] n2690_o;
  wire n2691_o;
  wire n2692_o;
  wire n2693_o;
  wire n2694_o;
  wire n2695_o;
  wire n2696_o;
  wire n2697_o;
  wire n2698_o;
  wire n2699_o;
  wire n2700_o;
  wire n2701_o;
  wire n2702_o;
  wire n2703_o;
  wire n2704_o;
  wire n2705_o;
  wire n2706_o;
  wire n2707_o;
  wire n2708_o;
  wire n2709_o;
  wire n2710_o;
  wire n2711_o;
  wire n2712_o;
  wire n2713_o;
  wire n2714_o;
  wire n2715_o;
  wire n2716_o;
  wire n2717_o;
  wire n2718_o;
  wire n2719_o;
  wire n2720_o;
  wire n2721_o;
  wire n2722_o;
  wire n2723_o;
  wire n2724_o;
  wire n2725_o;
  wire [3:0] n2726_o;
  wire [3:0] n2727_o;
  wire [3:0] n2728_o;
  wire [3:0] n2729_o;
  wire [3:0] n2730_o;
  wire [3:0] n2731_o;
  wire [3:0] n2732_o;
  wire [3:0] n2733_o;
  wire [2:0] n2734_o;
  wire [15:0] n2735_o;
  wire [15:0] n2736_o;
  wire [34:0] n2737_o;
  wire [34:0] n2738_o;
  wire [34:0] n2739_o;
  wire [35:0] n2740_o;
  wire [34:0] n2741_o;
  wire n2742_o;
  wire n2743_o;
  wire n2744_o;
  wire n2745_o;
  wire n2746_o;
  wire n2747_o;
  wire n2748_o;
  wire n2749_o;
  wire n2750_o;
  wire n2751_o;
  wire n2752_o;
  wire n2753_o;
  wire n2754_o;
  wire n2755_o;
  wire n2756_o;
  wire n2757_o;
  wire n2758_o;
  wire n2759_o;
  wire n2760_o;
  wire n2761_o;
  wire n2762_o;
  wire n2763_o;
  wire n2764_o;
  wire n2765_o;
  wire n2766_o;
  wire n2767_o;
  wire n2768_o;
  wire n2769_o;
  wire n2770_o;
  wire n2771_o;
  wire n2772_o;
  wire n2773_o;
  wire n2774_o;
  wire n2775_o;
  wire n2776_o;
  wire [3:0] n2777_o;
  wire [3:0] n2778_o;
  wire [3:0] n2779_o;
  wire [3:0] n2780_o;
  wire [3:0] n2781_o;
  wire [3:0] n2782_o;
  wire [3:0] n2783_o;
  wire [3:0] n2784_o;
  wire [2:0] n2785_o;
  wire [15:0] n2786_o;
  wire [15:0] n2787_o;
  wire [34:0] n2788_o;
  wire [34:0] n2789_o;
  wire [34:0] n2790_o;
  wire [35:0] n2791_o;
  wire [34:0] n2792_o;
  wire n2793_o;
  wire n2794_o;
  wire n2795_o;
  wire n2796_o;
  wire n2797_o;
  wire n2798_o;
  wire n2799_o;
  wire n2800_o;
  wire n2801_o;
  wire n2802_o;
  wire n2803_o;
  wire n2804_o;
  wire n2805_o;
  wire n2806_o;
  wire n2807_o;
  wire n2808_o;
  wire n2809_o;
  wire n2810_o;
  wire n2811_o;
  wire n2812_o;
  wire n2813_o;
  wire n2814_o;
  wire n2815_o;
  wire n2816_o;
  wire n2817_o;
  wire n2818_o;
  wire n2819_o;
  wire n2820_o;
  wire n2821_o;
  wire n2822_o;
  wire n2823_o;
  wire n2824_o;
  wire n2825_o;
  wire n2826_o;
  wire n2827_o;
  wire [3:0] n2828_o;
  wire [3:0] n2829_o;
  wire [3:0] n2830_o;
  wire [3:0] n2831_o;
  wire [3:0] n2832_o;
  wire [3:0] n2833_o;
  wire [3:0] n2834_o;
  wire [3:0] n2835_o;
  wire [2:0] n2836_o;
  wire [15:0] n2837_o;
  wire [15:0] n2838_o;
  wire [34:0] n2839_o;
  wire [34:0] n2840_o;
  wire [34:0] n2841_o;
  wire [179:0] n2847_o;
  assign outport = n2847_o;
  /* routers/synchronous/xbar.vhd:59:16  */
  assign sel0 = n1822_o; // (signal)
  /* routers/synchronous/xbar.vhd:59:22  */
  assign sel1 = n1823_o; // (signal)
  /* routers/synchronous/xbar.vhd:59:28  */
  assign sel2 = n1824_o; // (signal)
  /* routers/synchronous/xbar.vhd:59:34  */
  assign sel3 = n1825_o; // (signal)
  /* routers/synchronous/xbar.vhd:59:40  */
  assign sel4 = n1826_o; // (signal)
  /* routers/synchronous/xbar.vhd:61:21  */
  assign n1822_o = func[3:0];
  /* routers/synchronous/xbar.vhd:62:21  */
  assign n1823_o = func[7:4];
  /* routers/synchronous/xbar.vhd:63:21  */
  assign n1824_o = func[11:8];
  /* routers/synchronous/xbar.vhd:64:21  */
  assign n1825_o = func[15:12];
  /* routers/synchronous/xbar.vhd:65:21  */
  assign n1826_o = func[19:16];
  /* routers/synchronous/xbar.vhd:67:35  */
  assign n1827_o = inport[71:36];
  /* routers/synchronous/xbar.vhd:67:39  */
  assign n1828_o = n1827_o[35:1];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1829_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1830_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1831_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1832_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1833_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1834_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1835_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1836_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1837_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1838_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1839_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1840_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1841_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1842_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1843_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1844_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1845_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1846_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1847_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1848_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1849_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1850_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1851_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1852_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1853_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1854_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1855_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1856_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1857_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1858_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1859_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1860_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1861_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1862_o = sel1[0];
  /* routers/synchronous/xbar.vhd:67:67  */
  assign n1863_o = sel1[0];
  assign n1864_o = {n1863_o, n1862_o, n1861_o, n1860_o};
  assign n1865_o = {n1859_o, n1858_o, n1857_o, n1856_o};
  assign n1866_o = {n1855_o, n1854_o, n1853_o, n1852_o};
  assign n1867_o = {n1851_o, n1850_o, n1849_o, n1848_o};
  assign n1868_o = {n1847_o, n1846_o, n1845_o, n1844_o};
  assign n1869_o = {n1843_o, n1842_o, n1841_o, n1840_o};
  assign n1870_o = {n1839_o, n1838_o, n1837_o, n1836_o};
  assign n1871_o = {n1835_o, n1834_o, n1833_o, n1832_o};
  assign n1872_o = {n1831_o, n1830_o, n1829_o};
  assign n1873_o = {n1864_o, n1865_o, n1866_o, n1867_o};
  assign n1874_o = {n1868_o, n1869_o, n1870_o, n1871_o};
  assign n1875_o = {n1873_o, n1874_o, n1872_o};
  /* routers/synchronous/xbar.vhd:67:44  */
  assign n1876_o = n1828_o & n1875_o;
  /* routers/synchronous/xbar.vhd:68:42  */
  assign n1877_o = inport[107:72];
  /* routers/synchronous/xbar.vhd:68:46  */
  assign n1878_o = n1877_o[35:1];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1879_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1880_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1881_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1882_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1883_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1884_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1885_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1886_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1887_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1888_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1889_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1890_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1891_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1892_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1893_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1894_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1895_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1896_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1897_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1898_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1899_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1900_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1901_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1902_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1903_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1904_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1905_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1906_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1907_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1908_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1909_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1910_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1911_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1912_o = sel2[0];
  /* routers/synchronous/xbar.vhd:68:74  */
  assign n1913_o = sel2[0];
  assign n1914_o = {n1913_o, n1912_o, n1911_o, n1910_o};
  assign n1915_o = {n1909_o, n1908_o, n1907_o, n1906_o};
  assign n1916_o = {n1905_o, n1904_o, n1903_o, n1902_o};
  assign n1917_o = {n1901_o, n1900_o, n1899_o, n1898_o};
  assign n1918_o = {n1897_o, n1896_o, n1895_o, n1894_o};
  assign n1919_o = {n1893_o, n1892_o, n1891_o, n1890_o};
  assign n1920_o = {n1889_o, n1888_o, n1887_o, n1886_o};
  assign n1921_o = {n1885_o, n1884_o, n1883_o, n1882_o};
  assign n1922_o = {n1881_o, n1880_o, n1879_o};
  assign n1923_o = {n1914_o, n1915_o, n1916_o, n1917_o};
  assign n1924_o = {n1918_o, n1919_o, n1920_o, n1921_o};
  assign n1925_o = {n1923_o, n1924_o, n1922_o};
  /* routers/synchronous/xbar.vhd:68:51  */
  assign n1926_o = n1878_o & n1925_o;
  /* routers/synchronous/xbar.vhd:67:73  */
  assign n1927_o = n1876_o | n1926_o;
  /* routers/synchronous/xbar.vhd:69:42  */
  assign n1928_o = inport[143:108];
  /* routers/synchronous/xbar.vhd:69:46  */
  assign n1929_o = n1928_o[35:1];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1930_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1931_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1932_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1933_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1934_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1935_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1936_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1937_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1938_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1939_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1940_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1941_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1942_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1943_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1944_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1945_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1946_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1947_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1948_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1949_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1950_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1951_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1952_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1953_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1954_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1955_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1956_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1957_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1958_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1959_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1960_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1961_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1962_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1963_o = sel3[0];
  /* routers/synchronous/xbar.vhd:69:74  */
  assign n1964_o = sel3[0];
  assign n1965_o = {n1964_o, n1963_o, n1962_o, n1961_o};
  assign n1966_o = {n1960_o, n1959_o, n1958_o, n1957_o};
  assign n1967_o = {n1956_o, n1955_o, n1954_o, n1953_o};
  assign n1968_o = {n1952_o, n1951_o, n1950_o, n1949_o};
  assign n1969_o = {n1948_o, n1947_o, n1946_o, n1945_o};
  assign n1970_o = {n1944_o, n1943_o, n1942_o, n1941_o};
  assign n1971_o = {n1940_o, n1939_o, n1938_o, n1937_o};
  assign n1972_o = {n1936_o, n1935_o, n1934_o, n1933_o};
  assign n1973_o = {n1932_o, n1931_o, n1930_o};
  assign n1974_o = {n1965_o, n1966_o, n1967_o, n1968_o};
  assign n1975_o = {n1969_o, n1970_o, n1971_o, n1972_o};
  assign n1976_o = {n1974_o, n1975_o, n1973_o};
  /* routers/synchronous/xbar.vhd:69:51  */
  assign n1977_o = n1929_o & n1976_o;
  /* routers/synchronous/xbar.vhd:68:80  */
  assign n1978_o = n1927_o | n1977_o;
  /* routers/synchronous/xbar.vhd:70:42  */
  assign n1979_o = inport[179:144];
  /* routers/synchronous/xbar.vhd:70:46  */
  assign n1980_o = n1979_o[35:1];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n1981_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n1982_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n1983_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n1984_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n1985_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n1986_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n1987_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n1988_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n1989_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n1990_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n1991_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n1992_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n1993_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n1994_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n1995_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n1996_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n1997_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n1998_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n1999_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n2000_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n2001_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n2002_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n2003_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n2004_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n2005_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n2006_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n2007_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n2008_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n2009_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n2010_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n2011_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n2012_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n2013_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n2014_o = sel4[0];
  /* routers/synchronous/xbar.vhd:70:74  */
  assign n2015_o = sel4[0];
  assign n2016_o = {n2015_o, n2014_o, n2013_o, n2012_o};
  assign n2017_o = {n2011_o, n2010_o, n2009_o, n2008_o};
  assign n2018_o = {n2007_o, n2006_o, n2005_o, n2004_o};
  assign n2019_o = {n2003_o, n2002_o, n2001_o, n2000_o};
  assign n2020_o = {n1999_o, n1998_o, n1997_o, n1996_o};
  assign n2021_o = {n1995_o, n1994_o, n1993_o, n1992_o};
  assign n2022_o = {n1991_o, n1990_o, n1989_o, n1988_o};
  assign n2023_o = {n1987_o, n1986_o, n1985_o, n1984_o};
  assign n2024_o = {n1983_o, n1982_o, n1981_o};
  assign n2025_o = {n2016_o, n2017_o, n2018_o, n2019_o};
  assign n2026_o = {n2020_o, n2021_o, n2022_o, n2023_o};
  assign n2027_o = {n2025_o, n2026_o, n2024_o};
  /* routers/synchronous/xbar.vhd:70:51  */
  assign n2028_o = n1980_o & n2027_o;
  /* routers/synchronous/xbar.vhd:69:80  */
  assign n2029_o = n1978_o | n2028_o;
  /* routers/synchronous/xbar.vhd:71:35  */
  assign n2030_o = inport[35:0];
  /* routers/synchronous/xbar.vhd:71:39  */
  assign n2031_o = n2030_o[35:1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2032_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2033_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2034_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2035_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2036_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2037_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2038_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2039_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2040_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2041_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2042_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2043_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2044_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2045_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2046_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2047_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2048_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2049_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2050_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2051_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2052_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2053_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2054_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2055_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2056_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2057_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2058_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2059_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2060_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2061_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2062_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2063_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2064_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2065_o = sel0[1];
  /* routers/synchronous/xbar.vhd:71:67  */
  assign n2066_o = sel0[1];
  assign n2067_o = {n2066_o, n2065_o, n2064_o, n2063_o};
  assign n2068_o = {n2062_o, n2061_o, n2060_o, n2059_o};
  assign n2069_o = {n2058_o, n2057_o, n2056_o, n2055_o};
  assign n2070_o = {n2054_o, n2053_o, n2052_o, n2051_o};
  assign n2071_o = {n2050_o, n2049_o, n2048_o, n2047_o};
  assign n2072_o = {n2046_o, n2045_o, n2044_o, n2043_o};
  assign n2073_o = {n2042_o, n2041_o, n2040_o, n2039_o};
  assign n2074_o = {n2038_o, n2037_o, n2036_o, n2035_o};
  assign n2075_o = {n2034_o, n2033_o, n2032_o};
  assign n2076_o = {n2067_o, n2068_o, n2069_o, n2070_o};
  assign n2077_o = {n2071_o, n2072_o, n2073_o, n2074_o};
  assign n2078_o = {n2076_o, n2077_o, n2075_o};
  /* routers/synchronous/xbar.vhd:71:44  */
  assign n2079_o = n2031_o & n2078_o;
  /* routers/synchronous/xbar.vhd:72:42  */
  assign n2080_o = inport[107:72];
  /* routers/synchronous/xbar.vhd:72:46  */
  assign n2081_o = n2080_o[35:1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2082_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2083_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2084_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2085_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2086_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2087_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2088_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2089_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2090_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2091_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2092_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2093_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2094_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2095_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2096_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2097_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2098_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2099_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2100_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2101_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2102_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2103_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2104_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2105_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2106_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2107_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2108_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2109_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2110_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2111_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2112_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2113_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2114_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2115_o = sel2[1];
  /* routers/synchronous/xbar.vhd:72:74  */
  assign n2116_o = sel2[1];
  assign n2117_o = {n2116_o, n2115_o, n2114_o, n2113_o};
  assign n2118_o = {n2112_o, n2111_o, n2110_o, n2109_o};
  assign n2119_o = {n2108_o, n2107_o, n2106_o, n2105_o};
  assign n2120_o = {n2104_o, n2103_o, n2102_o, n2101_o};
  assign n2121_o = {n2100_o, n2099_o, n2098_o, n2097_o};
  assign n2122_o = {n2096_o, n2095_o, n2094_o, n2093_o};
  assign n2123_o = {n2092_o, n2091_o, n2090_o, n2089_o};
  assign n2124_o = {n2088_o, n2087_o, n2086_o, n2085_o};
  assign n2125_o = {n2084_o, n2083_o, n2082_o};
  assign n2126_o = {n2117_o, n2118_o, n2119_o, n2120_o};
  assign n2127_o = {n2121_o, n2122_o, n2123_o, n2124_o};
  assign n2128_o = {n2126_o, n2127_o, n2125_o};
  /* routers/synchronous/xbar.vhd:72:51  */
  assign n2129_o = n2081_o & n2128_o;
  /* routers/synchronous/xbar.vhd:71:73  */
  assign n2130_o = n2079_o | n2129_o;
  /* routers/synchronous/xbar.vhd:73:42  */
  assign n2131_o = inport[143:108];
  /* routers/synchronous/xbar.vhd:73:46  */
  assign n2132_o = n2131_o[35:1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2133_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2134_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2135_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2136_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2137_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2138_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2139_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2140_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2141_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2142_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2143_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2144_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2145_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2146_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2147_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2148_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2149_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2150_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2151_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2152_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2153_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2154_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2155_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2156_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2157_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2158_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2159_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2160_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2161_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2162_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2163_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2164_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2165_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2166_o = sel3[1];
  /* routers/synchronous/xbar.vhd:73:74  */
  assign n2167_o = sel3[1];
  assign n2168_o = {n2167_o, n2166_o, n2165_o, n2164_o};
  assign n2169_o = {n2163_o, n2162_o, n2161_o, n2160_o};
  assign n2170_o = {n2159_o, n2158_o, n2157_o, n2156_o};
  assign n2171_o = {n2155_o, n2154_o, n2153_o, n2152_o};
  assign n2172_o = {n2151_o, n2150_o, n2149_o, n2148_o};
  assign n2173_o = {n2147_o, n2146_o, n2145_o, n2144_o};
  assign n2174_o = {n2143_o, n2142_o, n2141_o, n2140_o};
  assign n2175_o = {n2139_o, n2138_o, n2137_o, n2136_o};
  assign n2176_o = {n2135_o, n2134_o, n2133_o};
  assign n2177_o = {n2168_o, n2169_o, n2170_o, n2171_o};
  assign n2178_o = {n2172_o, n2173_o, n2174_o, n2175_o};
  assign n2179_o = {n2177_o, n2178_o, n2176_o};
  /* routers/synchronous/xbar.vhd:73:51  */
  assign n2180_o = n2132_o & n2179_o;
  /* routers/synchronous/xbar.vhd:72:80  */
  assign n2181_o = n2130_o | n2180_o;
  /* routers/synchronous/xbar.vhd:74:42  */
  assign n2182_o = inport[179:144];
  /* routers/synchronous/xbar.vhd:74:46  */
  assign n2183_o = n2182_o[35:1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2184_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2185_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2186_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2187_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2188_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2189_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2190_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2191_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2192_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2193_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2194_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2195_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2196_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2197_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2198_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2199_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2200_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2201_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2202_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2203_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2204_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2205_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2206_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2207_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2208_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2209_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2210_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2211_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2212_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2213_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2214_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2215_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2216_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2217_o = sel4[1];
  /* routers/synchronous/xbar.vhd:74:74  */
  assign n2218_o = sel4[1];
  assign n2219_o = {n2218_o, n2217_o, n2216_o, n2215_o};
  assign n2220_o = {n2214_o, n2213_o, n2212_o, n2211_o};
  assign n2221_o = {n2210_o, n2209_o, n2208_o, n2207_o};
  assign n2222_o = {n2206_o, n2205_o, n2204_o, n2203_o};
  assign n2223_o = {n2202_o, n2201_o, n2200_o, n2199_o};
  assign n2224_o = {n2198_o, n2197_o, n2196_o, n2195_o};
  assign n2225_o = {n2194_o, n2193_o, n2192_o, n2191_o};
  assign n2226_o = {n2190_o, n2189_o, n2188_o, n2187_o};
  assign n2227_o = {n2186_o, n2185_o, n2184_o};
  assign n2228_o = {n2219_o, n2220_o, n2221_o, n2222_o};
  assign n2229_o = {n2223_o, n2224_o, n2225_o, n2226_o};
  assign n2230_o = {n2228_o, n2229_o, n2227_o};
  /* routers/synchronous/xbar.vhd:74:51  */
  assign n2231_o = n2183_o & n2230_o;
  /* routers/synchronous/xbar.vhd:73:80  */
  assign n2232_o = n2181_o | n2231_o;
  /* routers/synchronous/xbar.vhd:75:35  */
  assign n2233_o = inport[35:0];
  /* routers/synchronous/xbar.vhd:75:39  */
  assign n2234_o = n2233_o[35:1];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2235_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2236_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2237_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2238_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2239_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2240_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2241_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2242_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2243_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2244_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2245_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2246_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2247_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2248_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2249_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2250_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2251_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2252_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2253_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2254_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2255_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2256_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2257_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2258_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2259_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2260_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2261_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2262_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2263_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2264_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2265_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2266_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2267_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2268_o = sel0[2];
  /* routers/synchronous/xbar.vhd:75:67  */
  assign n2269_o = sel0[2];
  assign n2270_o = {n2269_o, n2268_o, n2267_o, n2266_o};
  assign n2271_o = {n2265_o, n2264_o, n2263_o, n2262_o};
  assign n2272_o = {n2261_o, n2260_o, n2259_o, n2258_o};
  assign n2273_o = {n2257_o, n2256_o, n2255_o, n2254_o};
  assign n2274_o = {n2253_o, n2252_o, n2251_o, n2250_o};
  assign n2275_o = {n2249_o, n2248_o, n2247_o, n2246_o};
  assign n2276_o = {n2245_o, n2244_o, n2243_o, n2242_o};
  assign n2277_o = {n2241_o, n2240_o, n2239_o, n2238_o};
  assign n2278_o = {n2237_o, n2236_o, n2235_o};
  assign n2279_o = {n2270_o, n2271_o, n2272_o, n2273_o};
  assign n2280_o = {n2274_o, n2275_o, n2276_o, n2277_o};
  assign n2281_o = {n2279_o, n2280_o, n2278_o};
  /* routers/synchronous/xbar.vhd:75:44  */
  assign n2282_o = n2234_o & n2281_o;
  /* routers/synchronous/xbar.vhd:76:42  */
  assign n2283_o = inport[71:36];
  /* routers/synchronous/xbar.vhd:76:46  */
  assign n2284_o = n2283_o[35:1];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2285_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2286_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2287_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2288_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2289_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2290_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2291_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2292_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2293_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2294_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2295_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2296_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2297_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2298_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2299_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2300_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2301_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2302_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2303_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2304_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2305_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2306_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2307_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2308_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2309_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2310_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2311_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2312_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2313_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2314_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2315_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2316_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2317_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2318_o = sel1[2];
  /* routers/synchronous/xbar.vhd:76:74  */
  assign n2319_o = sel1[2];
  assign n2320_o = {n2319_o, n2318_o, n2317_o, n2316_o};
  assign n2321_o = {n2315_o, n2314_o, n2313_o, n2312_o};
  assign n2322_o = {n2311_o, n2310_o, n2309_o, n2308_o};
  assign n2323_o = {n2307_o, n2306_o, n2305_o, n2304_o};
  assign n2324_o = {n2303_o, n2302_o, n2301_o, n2300_o};
  assign n2325_o = {n2299_o, n2298_o, n2297_o, n2296_o};
  assign n2326_o = {n2295_o, n2294_o, n2293_o, n2292_o};
  assign n2327_o = {n2291_o, n2290_o, n2289_o, n2288_o};
  assign n2328_o = {n2287_o, n2286_o, n2285_o};
  assign n2329_o = {n2320_o, n2321_o, n2322_o, n2323_o};
  assign n2330_o = {n2324_o, n2325_o, n2326_o, n2327_o};
  assign n2331_o = {n2329_o, n2330_o, n2328_o};
  /* routers/synchronous/xbar.vhd:76:51  */
  assign n2332_o = n2284_o & n2331_o;
  /* routers/synchronous/xbar.vhd:75:73  */
  assign n2333_o = n2282_o | n2332_o;
  /* routers/synchronous/xbar.vhd:77:42  */
  assign n2334_o = inport[143:108];
  /* routers/synchronous/xbar.vhd:77:46  */
  assign n2335_o = n2334_o[35:1];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2336_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2337_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2338_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2339_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2340_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2341_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2342_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2343_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2344_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2345_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2346_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2347_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2348_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2349_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2350_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2351_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2352_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2353_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2354_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2355_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2356_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2357_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2358_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2359_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2360_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2361_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2362_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2363_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2364_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2365_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2366_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2367_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2368_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2369_o = sel3[2];
  /* routers/synchronous/xbar.vhd:77:74  */
  assign n2370_o = sel3[2];
  assign n2371_o = {n2370_o, n2369_o, n2368_o, n2367_o};
  assign n2372_o = {n2366_o, n2365_o, n2364_o, n2363_o};
  assign n2373_o = {n2362_o, n2361_o, n2360_o, n2359_o};
  assign n2374_o = {n2358_o, n2357_o, n2356_o, n2355_o};
  assign n2375_o = {n2354_o, n2353_o, n2352_o, n2351_o};
  assign n2376_o = {n2350_o, n2349_o, n2348_o, n2347_o};
  assign n2377_o = {n2346_o, n2345_o, n2344_o, n2343_o};
  assign n2378_o = {n2342_o, n2341_o, n2340_o, n2339_o};
  assign n2379_o = {n2338_o, n2337_o, n2336_o};
  assign n2380_o = {n2371_o, n2372_o, n2373_o, n2374_o};
  assign n2381_o = {n2375_o, n2376_o, n2377_o, n2378_o};
  assign n2382_o = {n2380_o, n2381_o, n2379_o};
  /* routers/synchronous/xbar.vhd:77:51  */
  assign n2383_o = n2335_o & n2382_o;
  /* routers/synchronous/xbar.vhd:76:80  */
  assign n2384_o = n2333_o | n2383_o;
  /* routers/synchronous/xbar.vhd:78:42  */
  assign n2385_o = inport[179:144];
  /* routers/synchronous/xbar.vhd:78:46  */
  assign n2386_o = n2385_o[35:1];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2387_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2388_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2389_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2390_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2391_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2392_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2393_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2394_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2395_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2396_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2397_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2398_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2399_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2400_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2401_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2402_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2403_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2404_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2405_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2406_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2407_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2408_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2409_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2410_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2411_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2412_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2413_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2414_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2415_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2416_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2417_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2418_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2419_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2420_o = sel4[2];
  /* routers/synchronous/xbar.vhd:78:74  */
  assign n2421_o = sel4[2];
  assign n2422_o = {n2421_o, n2420_o, n2419_o, n2418_o};
  assign n2423_o = {n2417_o, n2416_o, n2415_o, n2414_o};
  assign n2424_o = {n2413_o, n2412_o, n2411_o, n2410_o};
  assign n2425_o = {n2409_o, n2408_o, n2407_o, n2406_o};
  assign n2426_o = {n2405_o, n2404_o, n2403_o, n2402_o};
  assign n2427_o = {n2401_o, n2400_o, n2399_o, n2398_o};
  assign n2428_o = {n2397_o, n2396_o, n2395_o, n2394_o};
  assign n2429_o = {n2393_o, n2392_o, n2391_o, n2390_o};
  assign n2430_o = {n2389_o, n2388_o, n2387_o};
  assign n2431_o = {n2422_o, n2423_o, n2424_o, n2425_o};
  assign n2432_o = {n2426_o, n2427_o, n2428_o, n2429_o};
  assign n2433_o = {n2431_o, n2432_o, n2430_o};
  /* routers/synchronous/xbar.vhd:78:51  */
  assign n2434_o = n2386_o & n2433_o;
  /* routers/synchronous/xbar.vhd:77:80  */
  assign n2435_o = n2384_o | n2434_o;
  /* routers/synchronous/xbar.vhd:79:35  */
  assign n2436_o = inport[35:0];
  /* routers/synchronous/xbar.vhd:79:39  */
  assign n2437_o = n2436_o[35:1];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2438_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2439_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2440_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2441_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2442_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2443_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2444_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2445_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2446_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2447_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2448_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2449_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2450_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2451_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2452_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2453_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2454_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2455_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2456_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2457_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2458_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2459_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2460_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2461_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2462_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2463_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2464_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2465_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2466_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2467_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2468_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2469_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2470_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2471_o = sel0[3];
  /* routers/synchronous/xbar.vhd:79:67  */
  assign n2472_o = sel0[3];
  assign n2473_o = {n2472_o, n2471_o, n2470_o, n2469_o};
  assign n2474_o = {n2468_o, n2467_o, n2466_o, n2465_o};
  assign n2475_o = {n2464_o, n2463_o, n2462_o, n2461_o};
  assign n2476_o = {n2460_o, n2459_o, n2458_o, n2457_o};
  assign n2477_o = {n2456_o, n2455_o, n2454_o, n2453_o};
  assign n2478_o = {n2452_o, n2451_o, n2450_o, n2449_o};
  assign n2479_o = {n2448_o, n2447_o, n2446_o, n2445_o};
  assign n2480_o = {n2444_o, n2443_o, n2442_o, n2441_o};
  assign n2481_o = {n2440_o, n2439_o, n2438_o};
  assign n2482_o = {n2473_o, n2474_o, n2475_o, n2476_o};
  assign n2483_o = {n2477_o, n2478_o, n2479_o, n2480_o};
  assign n2484_o = {n2482_o, n2483_o, n2481_o};
  /* routers/synchronous/xbar.vhd:79:44  */
  assign n2485_o = n2437_o & n2484_o;
  /* routers/synchronous/xbar.vhd:80:42  */
  assign n2486_o = inport[71:36];
  /* routers/synchronous/xbar.vhd:80:46  */
  assign n2487_o = n2486_o[35:1];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2488_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2489_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2490_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2491_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2492_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2493_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2494_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2495_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2496_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2497_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2498_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2499_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2500_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2501_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2502_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2503_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2504_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2505_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2506_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2507_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2508_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2509_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2510_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2511_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2512_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2513_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2514_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2515_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2516_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2517_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2518_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2519_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2520_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2521_o = sel1[3];
  /* routers/synchronous/xbar.vhd:80:74  */
  assign n2522_o = sel1[3];
  assign n2523_o = {n2522_o, n2521_o, n2520_o, n2519_o};
  assign n2524_o = {n2518_o, n2517_o, n2516_o, n2515_o};
  assign n2525_o = {n2514_o, n2513_o, n2512_o, n2511_o};
  assign n2526_o = {n2510_o, n2509_o, n2508_o, n2507_o};
  assign n2527_o = {n2506_o, n2505_o, n2504_o, n2503_o};
  assign n2528_o = {n2502_o, n2501_o, n2500_o, n2499_o};
  assign n2529_o = {n2498_o, n2497_o, n2496_o, n2495_o};
  assign n2530_o = {n2494_o, n2493_o, n2492_o, n2491_o};
  assign n2531_o = {n2490_o, n2489_o, n2488_o};
  assign n2532_o = {n2523_o, n2524_o, n2525_o, n2526_o};
  assign n2533_o = {n2527_o, n2528_o, n2529_o, n2530_o};
  assign n2534_o = {n2532_o, n2533_o, n2531_o};
  /* routers/synchronous/xbar.vhd:80:51  */
  assign n2535_o = n2487_o & n2534_o;
  /* routers/synchronous/xbar.vhd:79:73  */
  assign n2536_o = n2485_o | n2535_o;
  /* routers/synchronous/xbar.vhd:81:42  */
  assign n2537_o = inport[107:72];
  /* routers/synchronous/xbar.vhd:81:46  */
  assign n2538_o = n2537_o[35:1];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2539_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2540_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2541_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2542_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2543_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2544_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2545_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2546_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2547_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2548_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2549_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2550_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2551_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2552_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2553_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2554_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2555_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2556_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2557_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2558_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2559_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2560_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2561_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2562_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2563_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2564_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2565_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2566_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2567_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2568_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2569_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2570_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2571_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2572_o = sel2[3];
  /* routers/synchronous/xbar.vhd:81:74  */
  assign n2573_o = sel2[3];
  assign n2574_o = {n2573_o, n2572_o, n2571_o, n2570_o};
  assign n2575_o = {n2569_o, n2568_o, n2567_o, n2566_o};
  assign n2576_o = {n2565_o, n2564_o, n2563_o, n2562_o};
  assign n2577_o = {n2561_o, n2560_o, n2559_o, n2558_o};
  assign n2578_o = {n2557_o, n2556_o, n2555_o, n2554_o};
  assign n2579_o = {n2553_o, n2552_o, n2551_o, n2550_o};
  assign n2580_o = {n2549_o, n2548_o, n2547_o, n2546_o};
  assign n2581_o = {n2545_o, n2544_o, n2543_o, n2542_o};
  assign n2582_o = {n2541_o, n2540_o, n2539_o};
  assign n2583_o = {n2574_o, n2575_o, n2576_o, n2577_o};
  assign n2584_o = {n2578_o, n2579_o, n2580_o, n2581_o};
  assign n2585_o = {n2583_o, n2584_o, n2582_o};
  /* routers/synchronous/xbar.vhd:81:51  */
  assign n2586_o = n2538_o & n2585_o;
  /* routers/synchronous/xbar.vhd:80:80  */
  assign n2587_o = n2536_o | n2586_o;
  /* routers/synchronous/xbar.vhd:82:42  */
  assign n2588_o = inport[179:144];
  /* routers/synchronous/xbar.vhd:82:46  */
  assign n2589_o = n2588_o[35:1];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2590_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2591_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2592_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2593_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2594_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2595_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2596_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2597_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2598_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2599_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2600_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2601_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2602_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2603_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2604_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2605_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2606_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2607_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2608_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2609_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2610_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2611_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2612_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2613_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2614_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2615_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2616_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2617_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2618_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2619_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2620_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2621_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2622_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2623_o = sel4[3];
  /* routers/synchronous/xbar.vhd:82:74  */
  assign n2624_o = sel4[3];
  assign n2625_o = {n2624_o, n2623_o, n2622_o, n2621_o};
  assign n2626_o = {n2620_o, n2619_o, n2618_o, n2617_o};
  assign n2627_o = {n2616_o, n2615_o, n2614_o, n2613_o};
  assign n2628_o = {n2612_o, n2611_o, n2610_o, n2609_o};
  assign n2629_o = {n2608_o, n2607_o, n2606_o, n2605_o};
  assign n2630_o = {n2604_o, n2603_o, n2602_o, n2601_o};
  assign n2631_o = {n2600_o, n2599_o, n2598_o, n2597_o};
  assign n2632_o = {n2596_o, n2595_o, n2594_o, n2593_o};
  assign n2633_o = {n2592_o, n2591_o, n2590_o};
  assign n2634_o = {n2625_o, n2626_o, n2627_o, n2628_o};
  assign n2635_o = {n2629_o, n2630_o, n2631_o, n2632_o};
  assign n2636_o = {n2634_o, n2635_o, n2633_o};
  /* routers/synchronous/xbar.vhd:82:51  */
  assign n2637_o = n2589_o & n2636_o;
  /* routers/synchronous/xbar.vhd:81:80  */
  assign n2638_o = n2587_o | n2637_o;
  /* routers/synchronous/xbar.vhd:83:35  */
  assign n2639_o = inport[35:0];
  /* routers/synchronous/xbar.vhd:83:39  */
  assign n2640_o = n2639_o[35:1];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2641_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2642_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2643_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2644_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2645_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2646_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2647_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2648_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2649_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2650_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2651_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2652_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2653_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2654_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2655_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2656_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2657_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2658_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2659_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2660_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2661_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2662_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2663_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2664_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2665_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2666_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2667_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2668_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2669_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2670_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2671_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2672_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2673_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2674_o = sel0[0];
  /* routers/synchronous/xbar.vhd:83:67  */
  assign n2675_o = sel0[0];
  assign n2676_o = {n2675_o, n2674_o, n2673_o, n2672_o};
  assign n2677_o = {n2671_o, n2670_o, n2669_o, n2668_o};
  assign n2678_o = {n2667_o, n2666_o, n2665_o, n2664_o};
  assign n2679_o = {n2663_o, n2662_o, n2661_o, n2660_o};
  assign n2680_o = {n2659_o, n2658_o, n2657_o, n2656_o};
  assign n2681_o = {n2655_o, n2654_o, n2653_o, n2652_o};
  assign n2682_o = {n2651_o, n2650_o, n2649_o, n2648_o};
  assign n2683_o = {n2647_o, n2646_o, n2645_o, n2644_o};
  assign n2684_o = {n2643_o, n2642_o, n2641_o};
  assign n2685_o = {n2676_o, n2677_o, n2678_o, n2679_o};
  assign n2686_o = {n2680_o, n2681_o, n2682_o, n2683_o};
  assign n2687_o = {n2685_o, n2686_o, n2684_o};
  /* routers/synchronous/xbar.vhd:83:44  */
  assign n2688_o = n2640_o & n2687_o;
  /* routers/synchronous/xbar.vhd:84:42  */
  assign n2689_o = inport[71:36];
  /* routers/synchronous/xbar.vhd:84:46  */
  assign n2690_o = n2689_o[35:1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2691_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2692_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2693_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2694_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2695_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2696_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2697_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2698_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2699_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2700_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2701_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2702_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2703_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2704_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2705_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2706_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2707_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2708_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2709_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2710_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2711_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2712_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2713_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2714_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2715_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2716_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2717_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2718_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2719_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2720_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2721_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2722_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2723_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2724_o = sel1[1];
  /* routers/synchronous/xbar.vhd:84:74  */
  assign n2725_o = sel1[1];
  assign n2726_o = {n2725_o, n2724_o, n2723_o, n2722_o};
  assign n2727_o = {n2721_o, n2720_o, n2719_o, n2718_o};
  assign n2728_o = {n2717_o, n2716_o, n2715_o, n2714_o};
  assign n2729_o = {n2713_o, n2712_o, n2711_o, n2710_o};
  assign n2730_o = {n2709_o, n2708_o, n2707_o, n2706_o};
  assign n2731_o = {n2705_o, n2704_o, n2703_o, n2702_o};
  assign n2732_o = {n2701_o, n2700_o, n2699_o, n2698_o};
  assign n2733_o = {n2697_o, n2696_o, n2695_o, n2694_o};
  assign n2734_o = {n2693_o, n2692_o, n2691_o};
  assign n2735_o = {n2726_o, n2727_o, n2728_o, n2729_o};
  assign n2736_o = {n2730_o, n2731_o, n2732_o, n2733_o};
  assign n2737_o = {n2735_o, n2736_o, n2734_o};
  /* routers/synchronous/xbar.vhd:84:51  */
  assign n2738_o = n2690_o & n2737_o;
  /* routers/synchronous/xbar.vhd:83:73  */
  assign n2739_o = n2688_o | n2738_o;
  /* routers/synchronous/xbar.vhd:85:42  */
  assign n2740_o = inport[107:72];
  /* routers/synchronous/xbar.vhd:85:46  */
  assign n2741_o = n2740_o[35:1];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2742_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2743_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2744_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2745_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2746_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2747_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2748_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2749_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2750_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2751_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2752_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2753_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2754_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2755_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2756_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2757_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2758_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2759_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2760_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2761_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2762_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2763_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2764_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2765_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2766_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2767_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2768_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2769_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2770_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2771_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2772_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2773_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2774_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2775_o = sel2[2];
  /* routers/synchronous/xbar.vhd:85:74  */
  assign n2776_o = sel2[2];
  assign n2777_o = {n2776_o, n2775_o, n2774_o, n2773_o};
  assign n2778_o = {n2772_o, n2771_o, n2770_o, n2769_o};
  assign n2779_o = {n2768_o, n2767_o, n2766_o, n2765_o};
  assign n2780_o = {n2764_o, n2763_o, n2762_o, n2761_o};
  assign n2781_o = {n2760_o, n2759_o, n2758_o, n2757_o};
  assign n2782_o = {n2756_o, n2755_o, n2754_o, n2753_o};
  assign n2783_o = {n2752_o, n2751_o, n2750_o, n2749_o};
  assign n2784_o = {n2748_o, n2747_o, n2746_o, n2745_o};
  assign n2785_o = {n2744_o, n2743_o, n2742_o};
  assign n2786_o = {n2777_o, n2778_o, n2779_o, n2780_o};
  assign n2787_o = {n2781_o, n2782_o, n2783_o, n2784_o};
  assign n2788_o = {n2786_o, n2787_o, n2785_o};
  /* routers/synchronous/xbar.vhd:85:51  */
  assign n2789_o = n2741_o & n2788_o;
  /* routers/synchronous/xbar.vhd:84:80  */
  assign n2790_o = n2739_o | n2789_o;
  /* routers/synchronous/xbar.vhd:86:42  */
  assign n2791_o = inport[143:108];
  /* routers/synchronous/xbar.vhd:86:46  */
  assign n2792_o = n2791_o[35:1];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2793_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2794_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2795_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2796_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2797_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2798_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2799_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2800_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2801_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2802_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2803_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2804_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2805_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2806_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2807_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2808_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2809_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2810_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2811_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2812_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2813_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2814_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2815_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2816_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2817_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2818_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2819_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2820_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2821_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2822_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2823_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2824_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2825_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2826_o = sel3[3];
  /* routers/synchronous/xbar.vhd:86:74  */
  assign n2827_o = sel3[3];
  assign n2828_o = {n2827_o, n2826_o, n2825_o, n2824_o};
  assign n2829_o = {n2823_o, n2822_o, n2821_o, n2820_o};
  assign n2830_o = {n2819_o, n2818_o, n2817_o, n2816_o};
  assign n2831_o = {n2815_o, n2814_o, n2813_o, n2812_o};
  assign n2832_o = {n2811_o, n2810_o, n2809_o, n2808_o};
  assign n2833_o = {n2807_o, n2806_o, n2805_o, n2804_o};
  assign n2834_o = {n2803_o, n2802_o, n2801_o, n2800_o};
  assign n2835_o = {n2799_o, n2798_o, n2797_o, n2796_o};
  assign n2836_o = {n2795_o, n2794_o, n2793_o};
  assign n2837_o = {n2828_o, n2829_o, n2830_o, n2831_o};
  assign n2838_o = {n2832_o, n2833_o, n2834_o, n2835_o};
  assign n2839_o = {n2837_o, n2838_o, n2836_o};
  /* routers/synchronous/xbar.vhd:86:51  */
  assign n2840_o = n2792_o & n2839_o;
  /* routers/synchronous/xbar.vhd:85:80  */
  assign n2841_o = n2790_o | n2840_o;
  assign n2847_o = {n2841_o, 1'bZ, n2638_o, 1'bZ, n2435_o, 1'bZ, n2232_o, 1'bZ, n2029_o, 1'bZ};
endmodule

module hpu
  (input  clk,
   input  reset,
   input  inline_req,
   input  [34:0] inline_data,
   output outline_req,
   output [34:0] outline_data,
   output [3:0] sel);
  wire [35:0] n1760_o;
  wire n1762_o;
  wire [34:0] n1763_o;
  wire vld;
  wire sop;
  wire eop;
  wire [1:0] dest;
  wire [3:0] selint;
  wire [3:0] selintnext;
  wire [3:0] decodedsel;
  wire [34:0] outint;
  wire n1765_o;
  wire n1766_o;
  wire n1767_o;
  wire [1:0] n1768_o;
  wire n1771_o;
  wire n1772_o;
  wire n1776_o;
  wire n1777_o;
  wire n1781_o;
  wire n1782_o;
  wire n1786_o;
  wire n1787_o;
  wire [3:0] n1789_o;
  wire n1790_o;
  wire n1791_o;
  wire n1792_o;
  wire n1793_o;
  wire [3:0] n1794_o;
  wire [3:0] n1795_o;
  wire n1796_o;
  wire n1797_o;
  wire n1798_o;
  wire [3:0] n1799_o;
  wire [15:0] n1800_o;
  wire [18:0] n1802_o;
  wire [20:0] n1804_o;
  wire [13:0] n1805_o;
  wire [34:0] n1806_o;
  wire [34:0] n1807_o;
  wire [34:0] n1808_o;
  reg [3:0] n1816_q;
  wire [3:0] n1818_o;
  wire [35:0] n1820_o;
  assign outline_req = n1762_o;
  assign outline_data = n1763_o;
  assign sel = n1799_o;
  /* ni/config_bus.vhd:63:5  */
  assign n1760_o = {inline_data, inline_req};
  /* ni/config_bus.vhd:59:5  */
  assign n1762_o = n1820_o[0];
  /* ni/config_bus.vhd:57:5  */
  assign n1763_o = n1820_o[35:1];
  /* routers/synchronous/hpu.vhd:56:16  */
  assign vld = n1765_o; // (signal)
  /* routers/synchronous/hpu.vhd:57:16  */
  assign sop = n1766_o; // (signal)
  /* routers/synchronous/hpu.vhd:59:16  */
  assign eop = n1767_o; // (signal)
  /* routers/synchronous/hpu.vhd:60:16  */
  assign dest = n1768_o; // (signal)
  /* routers/synchronous/hpu.vhd:62:16  */
  assign selint = n1816_q; // (signal)
  /* routers/synchronous/hpu.vhd:62:24  */
  assign selintnext = n1789_o; // (signal)
  /* routers/synchronous/hpu.vhd:63:16  */
  assign decodedsel = n1818_o; // (signal)
  /* routers/synchronous/hpu.vhd:64:16  */
  assign outint = n1807_o; // (signal)
  /* routers/synchronous/hpu.vhd:66:27  */
  assign n1765_o = n1760_o[35];
  /* routers/synchronous/hpu.vhd:67:27  */
  assign n1766_o = n1760_o[34];
  /* routers/synchronous/hpu.vhd:69:27  */
  assign n1767_o = n1760_o[33];
  /* routers/synchronous/hpu.vhd:70:28  */
  assign n1768_o = n1760_o[2:1];
  /* routers/synchronous/hpu.vhd:74:40  */
  assign n1771_o = dest == 2'b00;
  /* routers/synchronous/hpu.vhd:74:30  */
  assign n1772_o = n1771_o ? 1'b1 : 1'b0;
  /* routers/synchronous/hpu.vhd:75:40  */
  assign n1776_o = dest == 2'b01;
  /* routers/synchronous/hpu.vhd:75:30  */
  assign n1777_o = n1776_o ? 1'b1 : 1'b0;
  /* routers/synchronous/hpu.vhd:76:40  */
  assign n1781_o = dest == 2'b10;
  /* routers/synchronous/hpu.vhd:76:30  */
  assign n1782_o = n1781_o ? 1'b1 : 1'b0;
  /* routers/synchronous/hpu.vhd:77:40  */
  assign n1786_o = dest == 2'b11;
  /* routers/synchronous/hpu.vhd:77:30  */
  assign n1787_o = n1786_o ? 1'b1 : 1'b0;
  /* routers/synchronous/hpu.vhd:79:34  */
  assign n1789_o = sop ? decodedsel : n1795_o;
  /* routers/synchronous/hpu.vhd:79:86  */
  assign n1790_o = vld | eop;
  /* routers/synchronous/hpu.vhd:79:86  */
  assign n1791_o = vld | eop;
  /* routers/synchronous/hpu.vhd:79:86  */
  assign n1792_o = vld | eop;
  /* routers/synchronous/hpu.vhd:79:86  */
  assign n1793_o = vld | eop;
  assign n1794_o = {n1793_o, n1792_o, n1791_o, n1790_o};
  /* routers/synchronous/hpu.vhd:79:62  */
  assign n1795_o = selint & n1794_o;
  /* routers/synchronous/hpu.vhd:80:38  */
  assign n1796_o = eop | vld;
  /* routers/synchronous/hpu.vhd:80:57  */
  assign n1797_o = ~sop;
  /* routers/synchronous/hpu.vhd:80:50  */
  assign n1798_o = n1796_o & n1797_o;
  /* routers/synchronous/hpu.vhd:80:23  */
  assign n1799_o = n1798_o ? selint : selintnext;
  /* routers/synchronous/hpu.vhd:81:38  */
  assign n1800_o = n1760_o[32:17];
  /* routers/synchronous/hpu.vhd:81:25  */
  assign n1802_o = {3'b110, n1800_o};
  /* routers/synchronous/hpu.vhd:81:53  */
  assign n1804_o = {n1802_o, 2'b00};
  /* routers/synchronous/hpu.vhd:81:73  */
  assign n1805_o = n1760_o[16:3];
  /* routers/synchronous/hpu.vhd:81:60  */
  assign n1806_o = {n1804_o, n1805_o};
  /* routers/synchronous/hpu.vhd:81:87  */
  assign n1807_o = sop ? n1806_o : n1808_o;
  /* routers/synchronous/hpu.vhd:81:114  */
  assign n1808_o = n1760_o[35:1];
  /* routers/synchronous/hpu.vhd:87:17  */
  always @(posedge clk or posedge reset)
    if (reset)
      n1816_q <= 4'b0000;
    else
      n1816_q <= selintnext;
  assign n1818_o = {n1787_o, n1782_o, n1777_o, n1772_o};
  assign n1820_o = {outint, 1'bZ};
endmodule

module config_bus
  (input  clk,
   input  reset,
   input  [2:0] ocp_config_m_mcmd,
   input  [31:0] ocp_config_m_maddr,
   input  [31:0] ocp_config_m_mdata,
   input  [3:0] ocp_config_m_mbyteen,
   input  ocp_config_m_mrespaccept,
   input  supervisor,
   input  [13:0] config_unit_addr,
   input  config_unit_en,
   input  config_unit_wr,
   input  [31:0] config_unit_wdata,
   input  [31:0] tdm_ctrl_rdata,
   input  tdm_ctrl_error,
   input  [31:0] sched_tbl_rdata,
   input  sched_tbl_error,
   input  [31:0] dma_tbl_rdata,
   input  dma_tbl_error,
   input  [31:0] mc_ctrl_rdata,
   input  mc_ctrl_error,
   input  [31:0] irq_unit_fifo_rdata,
   input  irq_unit_fifo_error,
   output [1:0] ocp_config_s_sresp,
   output [31:0] ocp_config_s_sdata,
   output ocp_config_s_scmdaccept,
   output [13:0] config_addr,
   output config_en,
   output config_wr,
   output [31:0] config_wdata,
   output tdm_ctrl_sel,
   output sched_tbl_sel,
   output dma_tbl_sel,
   output mc_ctrl_sel,
   output irq_unit_fifo_sel);
  wire [71:0] n1624_o;
  wire [1:0] n1626_o;
  wire [31:0] n1627_o;
  wire n1628_o;
  wire [47:0] n1629_o;
  wire [13:0] n1631_o;
  wire n1632_o;
  wire n1633_o;
  wire [31:0] n1634_o;
  wire [32:0] n1635_o;
  wire [32:0] n1637_o;
  wire [32:0] n1639_o;
  wire [32:0] n1641_o;
  wire [32:0] n1643_o;
  wire [1:0] next_ocp_resp;
  wire [1:0] ocp_resp_reg;
  wire [2:0] bank_id;
  wire [2:0] prev_bank_id;
  wire [31:0] n1646_o;
  wire [2:0] n1648_o;
  wire [13:0] n1649_o;
  wire n1650_o;
  wire n1651_o;
  wire [31:0] n1652_o;
  wire n1653_o;
  wire n1654_o;
  wire [2:0] n1655_o;
  wire n1657_o;
  wire n1658_o;
  wire [31:0] n1660_o;
  wire [2:0] n1661_o;
  wire [13:0] n1662_o;
  wire [2:0] n1665_o;
  wire n1667_o;
  wire n1668_o;
  wire [2:0] n1669_o;
  wire n1671_o;
  wire n1673_o;
  wire n1674_o;
  wire n1675_o;
  wire [47:0] n1676_o;
  wire [47:0] n1677_o;
  wire [47:0] n1678_o;
  wire [1:0] n1680_o;
  wire [2:0] n1681_o;
  wire n1683_o;
  wire n1684_o;
  wire n1685_o;
  wire [1:0] n1687_o;
  wire n1696_o;
  wire n1698_o;
  wire n1700_o;
  wire n1702_o;
  wire n1704_o;
  wire n1706_o;
  wire [5:0] n1707_o;
  reg n1710_o;
  reg n1714_o;
  reg n1718_o;
  reg n1722_o;
  reg n1726_o;
  wire [31:0] n1728_o;
  wire n1730_o;
  wire [31:0] n1731_o;
  wire n1733_o;
  wire [31:0] n1734_o;
  wire n1736_o;
  wire [31:0] n1737_o;
  wire n1739_o;
  wire [31:0] n1740_o;
  wire n1742_o;
  wire n1744_o;
  wire [5:0] n1745_o;
  reg [31:0] n1746_o;
  wire [1:0] n1751_o;
  wire [2:0] n1753_o;
  reg [1:0] n1757_q;
  reg [2:0] n1758_q;
  wire [34:0] n1759_o;
  assign ocp_config_s_sresp = n1626_o;
  assign ocp_config_s_sdata = n1627_o;
  assign ocp_config_s_scmdaccept = n1628_o;
  assign config_addr = n1631_o;
  assign config_en = n1632_o;
  assign config_wr = n1633_o;
  assign config_wdata = n1634_o;
  assign tdm_ctrl_sel = n1710_o;
  assign sched_tbl_sel = n1714_o;
  assign dma_tbl_sel = n1718_o;
  assign mc_ctrl_sel = n1722_o;
  assign irq_unit_fifo_sel = n1726_o;
  /* ni/spm_bus.vhd:50:17  */
  assign n1624_o = {ocp_config_m_mrespaccept, ocp_config_m_mbyteen, ocp_config_m_mdata, ocp_config_m_maddr, ocp_config_m_mcmd};
  /* ni/spm_bus.vhd:81:9  */
  assign n1626_o = n1759_o[1:0];
  assign n1627_o = n1759_o[33:2];
  /* ni/spm_bus.vhd:63:9  */
  assign n1628_o = n1759_o[34];
  /* ni/spm_bus.vhd:83:17  */
  assign n1629_o = {config_unit_wdata, config_unit_wr, config_unit_en, config_unit_addr};
  assign n1631_o = n1678_o[13:0];
  assign n1632_o = n1678_o[14];
  assign n1633_o = n1678_o[15];
  assign n1634_o = n1678_o[47:16];
  assign n1635_o = {tdm_ctrl_error, tdm_ctrl_rdata};
  assign n1637_o = {sched_tbl_error, sched_tbl_rdata};
  assign n1639_o = {dma_tbl_error, dma_tbl_rdata};
  assign n1641_o = {mc_ctrl_error, mc_ctrl_rdata};
  assign n1643_o = {irq_unit_fifo_error, irq_unit_fifo_rdata};
  /* ni/config_bus.vhd:88:8  */
  assign next_ocp_resp = n1687_o; // (signal)
  /* ni/config_bus.vhd:88:23  */
  assign ocp_resp_reg = n1757_q; // (signal)
  /* ni/config_bus.vhd:89:8  */
  assign bank_id = n1681_o; // (signal)
  /* ni/config_bus.vhd:89:17  */
  assign prev_bank_id = n1758_q; // (signal)
  /* ni/config_bus.vhd:105:55  */
  assign n1646_o = n1639_o[31:0];
  /* ni/config_bus.vhd:108:30  */
  assign n1648_o = n1629_o[13:11];
  /* ni/config_bus.vhd:110:30  */
  assign n1649_o = n1629_o[13:0];
  /* ni/config_bus.vhd:111:28  */
  assign n1650_o = n1629_o[14];
  /* ni/config_bus.vhd:112:28  */
  assign n1651_o = n1629_o[15];
  /* ni/config_bus.vhd:113:31  */
  assign n1652_o = n1629_o[47:16];
  /* ni/config_bus.vhd:120:18  */
  assign n1653_o = n1629_o[14];
  /* ni/config_bus.vhd:120:21  */
  assign n1654_o = ~n1653_o;
  /* ni/config_bus.vhd:120:44  */
  assign n1655_o = n1624_o[2:0];
  /* ni/config_bus.vhd:120:49  */
  assign n1657_o = n1655_o != 3'b000;
  /* ni/config_bus.vhd:120:27  */
  assign n1658_o = n1654_o & n1657_o;
  /* ni/config_bus.vhd:124:66  */
  assign n1660_o = n1624_o[66:35];
  /* ni/config_bus.vhd:126:43  */
  assign n1661_o = n1624_o[18:16];
  /* ni/config_bus.vhd:129:47  */
  assign n1662_o = n1624_o[18:5];
  /* ni/config_bus.vhd:134:21  */
  assign n1665_o = n1624_o[2:0];
  /* ni/config_bus.vhd:134:26  */
  assign n1667_o = n1665_o != 3'b000;
  /* ni/config_bus.vhd:134:42  */
  assign n1668_o = n1667_o & supervisor;
  /* ni/config_bus.vhd:135:21  */
  assign n1669_o = n1624_o[2:0];
  /* ni/config_bus.vhd:135:26  */
  assign n1671_o = n1669_o == 3'b001;
  /* ni/config_bus.vhd:134:5  */
  assign n1673_o = n1674_o ? 1'b1 : 1'b0;
  /* ni/config_bus.vhd:134:5  */
  assign n1674_o = n1668_o & n1671_o;
  /* ni/config_bus.vhd:120:3  */
  assign n1675_o = n1658_o ? 1'b1 : 1'b0;
  assign n1676_o = {n1660_o, n1673_o, 1'b1, n1662_o};
  assign n1677_o = {n1652_o, n1651_o, n1650_o, n1649_o};
  /* ni/config_bus.vhd:120:3  */
  assign n1678_o = n1658_o ? n1676_o : n1677_o;
  /* ni/config_bus.vhd:120:3  */
  assign n1680_o = n1658_o ? 2'b01 : ocp_resp_reg;
  /* ni/config_bus.vhd:120:3  */
  assign n1681_o = n1658_o ? n1661_o : n1648_o;
  /* ni/config_bus.vhd:161:20  */
  assign n1683_o = ocp_resp_reg != 2'b00;
  /* ni/config_bus.vhd:161:56  */
  assign n1684_o = n1624_o[71];
  /* ni/config_bus.vhd:161:38  */
  assign n1685_o = n1683_o & n1684_o;
  /* ni/config_bus.vhd:161:3  */
  assign n1687_o = n1685_o ? 2'b00 : n1680_o;
  /* ni/config_bus.vhd:177:5  */
  assign n1696_o = bank_id == 3'b000;
  /* ni/config_bus.vhd:179:5  */
  assign n1698_o = bank_id == 3'b001;
  /* ni/config_bus.vhd:181:5  */
  assign n1700_o = bank_id == 3'b010;
  /* ni/config_bus.vhd:183:5  */
  assign n1702_o = bank_id == 3'b011;
  /* ni/config_bus.vhd:185:5  */
  assign n1704_o = bank_id == 3'b100;
  /* ni/config_bus.vhd:187:5  */
  assign n1706_o = bank_id == 3'b111;
  assign n1707_o = {n1706_o, n1704_o, n1702_o, n1700_o, n1698_o, n1696_o};
  /* ni/config_bus.vhd:176:3  */
  always @*
    case (n1707_o)
      6'b100000: n1710_o <= 1'b0;
      6'b010000: n1710_o <= 1'b0;
      6'b001000: n1710_o <= 1'b0;
      6'b000100: n1710_o <= 1'b1;
      6'b000010: n1710_o <= 1'b0;
      6'b000001: n1710_o <= 1'b0;
      default: n1710_o <= 1'b0;
    endcase
  /* ni/config_bus.vhd:176:3  */
  always @*
    case (n1707_o)
      6'b100000: n1714_o <= 1'b0;
      6'b010000: n1714_o <= 1'b0;
      6'b001000: n1714_o <= 1'b0;
      6'b000100: n1714_o <= 1'b0;
      6'b000010: n1714_o <= 1'b1;
      6'b000001: n1714_o <= 1'b0;
      default: n1714_o <= 1'b0;
    endcase
  /* ni/config_bus.vhd:176:3  */
  always @*
    case (n1707_o)
      6'b100000: n1718_o <= 1'b0;
      6'b010000: n1718_o <= 1'b0;
      6'b001000: n1718_o <= 1'b0;
      6'b000100: n1718_o <= 1'b0;
      6'b000010: n1718_o <= 1'b0;
      6'b000001: n1718_o <= 1'b1;
      default: n1718_o <= 1'b0;
    endcase
  /* ni/config_bus.vhd:176:3  */
  always @*
    case (n1707_o)
      6'b100000: n1722_o <= 1'b0;
      6'b010000: n1722_o <= 1'b0;
      6'b001000: n1722_o <= 1'b1;
      6'b000100: n1722_o <= 1'b0;
      6'b000010: n1722_o <= 1'b0;
      6'b000001: n1722_o <= 1'b0;
      default: n1722_o <= 1'b0;
    endcase
  /* ni/config_bus.vhd:176:3  */
  always @*
    case (n1707_o)
      6'b100000: n1726_o <= 1'b0;
      6'b010000: n1726_o <= 1'b1;
      6'b001000: n1726_o <= 1'b0;
      6'b000100: n1726_o <= 1'b0;
      6'b000010: n1726_o <= 1'b0;
      6'b000001: n1726_o <= 1'b0;
      default: n1726_o <= 1'b0;
    endcase
  /* ni/config_bus.vhd:194:59  */
  assign n1728_o = n1639_o[31:0];
  /* ni/config_bus.vhd:193:5  */
  assign n1730_o = prev_bank_id == 3'b000;
  /* ni/config_bus.vhd:196:61  */
  assign n1731_o = n1637_o[31:0];
  /* ni/config_bus.vhd:195:5  */
  assign n1733_o = prev_bank_id == 3'b001;
  /* ni/config_bus.vhd:198:60  */
  assign n1734_o = n1635_o[31:0];
  /* ni/config_bus.vhd:197:5  */
  assign n1736_o = prev_bank_id == 3'b010;
  /* ni/config_bus.vhd:200:59  */
  assign n1737_o = n1641_o[31:0];
  /* ni/config_bus.vhd:199:5  */
  assign n1739_o = prev_bank_id == 3'b011;
  /* ni/config_bus.vhd:202:65  */
  assign n1740_o = n1643_o[31:0];
  /* ni/config_bus.vhd:201:5  */
  assign n1742_o = prev_bank_id == 3'b100;
  /* ni/config_bus.vhd:203:5  */
  assign n1744_o = prev_bank_id == 3'b111;
  assign n1745_o = {n1744_o, n1742_o, n1739_o, n1736_o, n1733_o, n1730_o};
  /* ni/config_bus.vhd:192:3  */
  always @*
    case (n1745_o)
      6'b100000: n1746_o <= n1646_o;
      6'b010000: n1746_o <= n1740_o;
      6'b001000: n1746_o <= n1737_o;
      6'b000100: n1746_o <= n1734_o;
      6'b000010: n1746_o <= n1731_o;
      6'b000001: n1746_o <= n1728_o;
      default: n1746_o <= n1646_o;
    endcase
  /* ni/config_bus.vhd:215:7  */
  assign n1751_o = reset ? 2'b00 : next_ocp_resp;
  /* ni/config_bus.vhd:215:7  */
  assign n1753_o = reset ? 3'b000 : bank_id;
  /* ni/config_bus.vhd:214:5  */
  always @(posedge clk)
    n1757_q <= n1751_o;
  /* ni/config_bus.vhd:214:5  */
  always @(posedge clk)
    n1758_q <= n1753_o;
  /* ni/config_bus.vhd:214:5  */
  assign n1759_o = {n1675_o, n1746_o, ocp_resp_reg};
endmodule

module spm_bus
  (input  clk,
   input  reset,
   input  [63:0] spm_slv_rdata,
   input  spm_slv_error,
   input  [13:0] tx_spm_addr,
   input  [1:0] tx_spm_en,
   input  tx_spm_wr,
   input  [63:0] tx_spm_wdata,
   input  [13:0] rx_spm_addr,
   input  [1:0] rx_spm_en,
   input  rx_spm_wr,
   input  [63:0] rx_spm_wdata,
   output [13:0] spm_addr,
   output [1:0] spm_en,
   output spm_wr,
   output [63:0] spm_wdata,
   output [63:0] tx_spm_slv_rdata,
   output tx_spm_slv_error);
  wire [64:0] n1568_o;
  wire [13:0] n1570_o;
  wire [1:0] n1571_o;
  wire n1572_o;
  wire [63:0] n1573_o;
  wire [63:0] n1575_o;
  wire n1576_o;
  wire [80:0] n1577_o;
  wire [80:0] n1578_o;
  wire [80:0] rx_spm_buff;
  wire n1581_o;
  wire n1582_o;
  wire n1583_o;
  wire n1584_o;
  wire n1585_o;
  wire n1586_o;
  wire n1587_o;
  wire n1588_o;
  wire n1589_o;
  wire [80:0] n1590_o;
  wire [80:0] n1591_o;
  wire [80:0] n1592_o;
  wire n1598_o;
  wire n1599_o;
  wire n1600_o;
  wire n1601_o;
  wire n1602_o;
  wire n1603_o;
  wire n1604_o;
  wire n1605_o;
  wire n1606_o;
  wire n1607_o;
  wire n1608_o;
  wire [13:0] n1609_o;
  wire [63:0] n1610_o;
  wire [80:0] n1611_o;
  wire [13:0] n1612_o;
  wire [13:0] n1613_o;
  wire [13:0] n1614_o;
  wire [1:0] n1615_o;
  wire [1:0] n1616_o;
  wire [64:0] n1617_o;
  wire [64:0] n1618_o;
  wire [64:0] n1619_o;
  wire [80:0] n1620_o;
  reg [80:0] n1623_q;
  assign spm_addr = n1570_o;
  assign spm_en = n1571_o;
  assign spm_wr = n1572_o;
  assign spm_wdata = n1573_o;
  assign tx_spm_slv_rdata = n1575_o;
  assign tx_spm_slv_error = n1576_o;
  /* ni/irq_fifo.vhd:146:9  */
  assign n1568_o = {spm_slv_error, spm_slv_rdata};
  /* ni/irq_fifo.vhd:53:17  */
  assign n1570_o = n1592_o[13:0];
  /* ni/irq_fifo.vhd:51:17  */
  assign n1571_o = n1592_o[15:14];
  assign n1572_o = n1592_o[16];
  assign n1573_o = n1592_o[80:17];
  assign n1575_o = n1568_o[63:0];
  /* ni/irq_fifo.vhd:216:9  */
  assign n1576_o = n1568_o[64];
  assign n1577_o = {tx_spm_wdata, tx_spm_wr, tx_spm_en, tx_spm_addr};
  /* ni/irq_fifo.vhd:200:9  */
  assign n1578_o = {rx_spm_wdata, rx_spm_wr, rx_spm_en, rx_spm_addr};
  /* ni/spm_bus.vhd:58:16  */
  assign rx_spm_buff = n1623_q; // (signal)
  /* ni/spm_bus.vhd:65:31  */
  assign n1581_o = n1577_o[14];
  /* ni/spm_bus.vhd:65:55  */
  assign n1582_o = n1577_o[15];
  /* ni/spm_bus.vhd:65:42  */
  assign n1583_o = n1581_o | n1582_o;
  /* ni/spm_bus.vhd:68:44  */
  assign n1584_o = rx_spm_buff[14];
  /* ni/spm_bus.vhd:68:73  */
  assign n1585_o = rx_spm_buff[15];
  /* ni/spm_bus.vhd:68:55  */
  assign n1586_o = n1584_o | n1585_o;
  /* ni/spm_bus.vhd:71:47  */
  assign n1587_o = n1578_o[14];
  /* ni/spm_bus.vhd:71:71  */
  assign n1588_o = n1578_o[15];
  /* ni/spm_bus.vhd:71:58  */
  assign n1589_o = n1587_o | n1588_o;
  /* ni/spm_bus.vhd:71:33  */
  assign n1590_o = n1589_o ? n1578_o : n1577_o;
  /* ni/spm_bus.vhd:68:25  */
  assign n1591_o = n1586_o ? rx_spm_buff : n1590_o;
  /* ni/spm_bus.vhd:65:17  */
  assign n1592_o = n1583_o ? n1577_o : n1591_o;
  /* ni/spm_bus.vhd:87:63  */
  assign n1598_o = n1578_o[14];
  /* ni/spm_bus.vhd:87:81  */
  assign n1599_o = n1577_o[14];
  /* ni/spm_bus.vhd:87:97  */
  assign n1600_o = n1577_o[15];
  /* ni/spm_bus.vhd:87:85  */
  assign n1601_o = n1599_o | n1600_o;
  /* ni/spm_bus.vhd:87:67  */
  assign n1602_o = n1598_o & n1601_o;
  /* ni/spm_bus.vhd:88:63  */
  assign n1603_o = n1578_o[15];
  /* ni/spm_bus.vhd:88:81  */
  assign n1604_o = n1577_o[14];
  /* ni/spm_bus.vhd:88:97  */
  assign n1605_o = n1577_o[15];
  /* ni/spm_bus.vhd:88:85  */
  assign n1606_o = n1604_o | n1605_o;
  /* ni/spm_bus.vhd:88:67  */
  assign n1607_o = n1603_o & n1606_o;
  /* ni/spm_bus.vhd:89:61  */
  assign n1608_o = n1578_o[16];
  /* ni/spm_bus.vhd:90:61  */
  assign n1609_o = n1578_o[13:0];
  /* ni/spm_bus.vhd:91:61  */
  assign n1610_o = n1578_o[80:17];
  assign n1611_o = {n1610_o, n1608_o, n1607_o, n1602_o, n1609_o};
  assign n1612_o = n1611_o[13:0];
  assign n1613_o = rx_spm_buff[13:0];
  /* ni/spm_bus.vhd:84:25  */
  assign n1614_o = reset ? n1613_o : n1612_o;
  assign n1615_o = n1611_o[15:14];
  /* ni/spm_bus.vhd:84:25  */
  assign n1616_o = reset ? 2'b00 : n1615_o;
  assign n1617_o = n1611_o[80:16];
  assign n1618_o = rx_spm_buff[80:16];
  /* ni/spm_bus.vhd:84:25  */
  assign n1619_o = reset ? n1618_o : n1617_o;
  assign n1620_o = {n1619_o, n1616_o, n1614_o};
  /* ni/spm_bus.vhd:83:17  */
  always @(posedge clk)
    n1623_q <= n1620_o;
endmodule

module irq_fifo
  (input  clk,
   input  reset,
   input  [13:0] config_addr,
   input  config_en,
   input  config_wr,
   input  [31:0] config_wdata,
   input  sel,
   input  irq_data_fifo_data_valid,
   input  irq_irq_fifo_data_valid,
   input  [13:0] irq_data_fifo_data,
   output [31:0] config_slv_rdata,
   output config_slv_error,
   output irq_irq_sig,
   output irq_data_sig);
  wire [47:0] n1403_o;
  wire [31:0] n1405_o;
  wire n1406_o;
  wire irq_not_empty;
  wire data_not_empty;
  wire next_error;
  wire irq_read;
  wire data_read;
  wire irq_not_full;
  wire data_not_full;
  wire [4:0] data_w_ptr;
  wire [4:0] data_r_ptr;
  wire [4:0] irq_w_ptr;
  wire [4:0] irq_r_ptr;
  wire [4:0] w_ptr;
  wire [4:0] r_ptr;
  wire [13:0] w_data;
  wire n1411_o;
  wire n1412_o;
  wire n1415_o;
  wire n1416_o;
  wire [4:0] n1420_o;
  wire n1421_o;
  wire n1423_o;
  wire n1425_o;
  wire n1426_o;
  wire n1427_o;
  wire n1428_o;
  wire [4:0] n1432_o;
  wire n1433_o;
  wire n1435_o;
  wire n1437_o;
  wire n1438_o;
  wire n1439_o;
  wire n1440_o;
  wire n1442_o;
  wire [4:0] n1443_o;
  wire n1446_o;
  wire n1447_o;
  wire n1448_o;
  wire n1449_o;
  wire [10:0] n1450_o;
  wire n1452_o;
  wire n1454_o;
  wire [1:0] n1455_o;
  reg n1458_o;
  reg n1461_o;
  reg n1464_o;
  reg [4:0] n1465_o;
  wire n1467_o;
  wire n1469_o;
  wire n1471_o;
  wire [4:0] n1472_o;
  wire n1474_o;
  wire n1477_o;
  wire n1480_o;
  wire n1482_o;
  wire n1484_o;
  wire n1485_o;
  wire n1486_o;
  localparam n1488_o = 1'b0;
  localparam [13:0] n1489_o = 14'b00000000000000;
  wire [13:0] tdpram_n1490;
  wire [13:0] tdpram_a_dout;
  wire [13:0] tdpram_b_dout;
  wire n1497_o;
  wire n1499_o;
  wire [4:0] n1501_o;
  wire [4:0] n1503_o;
  wire [4:0] n1504_o;
  wire [4:0] n1506_o;
  reg [4:0] n1509_q;
  wire n1513_o;
  wire n1515_o;
  wire [4:0] n1517_o;
  wire [4:0] n1519_o;
  wire [4:0] n1520_o;
  wire [4:0] n1522_o;
  reg [4:0] n1525_q;
  wire n1529_o;
  wire n1531_o;
  wire [4:0] n1533_o;
  wire [4:0] n1535_o;
  wire [4:0] n1536_o;
  wire [4:0] n1538_o;
  reg [4:0] n1541_q;
  wire n1545_o;
  wire n1547_o;
  wire [4:0] n1549_o;
  wire [4:0] n1551_o;
  wire [4:0] n1552_o;
  wire [4:0] n1554_o;
  reg [4:0] n1557_q;
  wire n1562_o;
  reg n1566_q;
  wire [32:0] n1567_o;
  assign config_slv_rdata = n1405_o;
  assign config_slv_error = n1406_o;
  assign irq_irq_sig = irq_not_empty;
  assign irq_data_sig = data_not_empty;
  /* ni/rx_unit.vhd:55:17  */
  assign n1403_o = {config_wdata, config_wr, config_en, config_addr};
  /* ni/rx_unit.vhd:52:17  */
  assign n1405_o = n1567_o[31:0];
  /* ni/rx_unit.vhd:50:17  */
  assign n1406_o = n1567_o[32];
  /* ni/irq_fifo.vhd:94:16  */
  assign irq_not_empty = n1412_o; // (signal)
  /* ni/irq_fifo.vhd:94:31  */
  assign data_not_empty = n1416_o; // (signal)
  /* ni/irq_fifo.vhd:94:47  */
  assign next_error = n1474_o; // (signal)
  /* ni/irq_fifo.vhd:94:59  */
  assign irq_read = n1477_o; // (signal)
  /* ni/irq_fifo.vhd:94:69  */
  assign data_read = n1480_o; // (signal)
  /* ni/irq_fifo.vhd:94:80  */
  assign irq_not_full = n1428_o; // (signal)
  /* ni/irq_fifo.vhd:94:94  */
  assign data_not_full = n1440_o; // (signal)
  /* ni/irq_fifo.vhd:95:16  */
  assign data_w_ptr = n1525_q; // (signal)
  /* ni/irq_fifo.vhd:95:28  */
  assign data_r_ptr = n1557_q; // (signal)
  /* ni/irq_fifo.vhd:95:40  */
  assign irq_w_ptr = n1509_q; // (signal)
  /* ni/irq_fifo.vhd:95:51  */
  assign irq_r_ptr = n1541_q; // (signal)
  /* ni/irq_fifo.vhd:95:62  */
  assign w_ptr = n1443_o; // (signal)
  /* ni/irq_fifo.vhd:95:69  */
  assign r_ptr = n1472_o; // (signal)
  /* ni/irq_fifo.vhd:96:16  */
  assign w_data = irq_data_fifo_data; // (signal)
  /* ni/irq_fifo.vhd:106:46  */
  assign n1411_o = irq_w_ptr == irq_r_ptr;
  /* ni/irq_fifo.vhd:106:31  */
  assign n1412_o = n1411_o ? 1'b0 : 1'b1;
  /* ni/irq_fifo.vhd:107:47  */
  assign n1415_o = data_w_ptr == data_r_ptr;
  /* ni/irq_fifo.vhd:107:31  */
  assign n1416_o = n1415_o ? 1'b0 : 1'b1;
  /* ni/irq_fifo.vhd:109:59  */
  assign n1420_o = irq_r_ptr - 5'b00001;
  /* ni/irq_fifo.vhd:109:47  */
  assign n1421_o = irq_w_ptr == n1420_o;
  /* ni/irq_fifo.vhd:109:78  */
  assign n1423_o = irq_w_ptr == 5'b01111;
  /* ni/irq_fifo.vhd:109:146  */
  assign n1425_o = irq_r_ptr == 5'b00000;
  /* ni/irq_fifo.vhd:109:132  */
  assign n1426_o = n1423_o & n1425_o;
  /* ni/irq_fifo.vhd:109:64  */
  assign n1427_o = n1421_o | n1426_o;
  /* ni/irq_fifo.vhd:109:30  */
  assign n1428_o = n1427_o ? 1'b0 : 1'b1;
  /* ni/irq_fifo.vhd:110:61  */
  assign n1432_o = data_r_ptr + 5'b00001;
  /* ni/irq_fifo.vhd:110:48  */
  assign n1433_o = data_w_ptr == n1432_o;
  /* ni/irq_fifo.vhd:110:81  */
  assign n1435_o = data_w_ptr == 5'b10000;
  /* ni/irq_fifo.vhd:110:151  */
  assign n1437_o = data_r_ptr == 5'b11111;
  /* ni/irq_fifo.vhd:110:136  */
  assign n1438_o = n1435_o & n1437_o;
  /* ni/irq_fifo.vhd:110:66  */
  assign n1439_o = n1433_o | n1438_o;
  /* ni/irq_fifo.vhd:110:30  */
  assign n1440_o = n1439_o ? 1'b0 : 1'b1;
  /* ni/irq_fifo.vhd:113:59  */
  assign n1442_o = ~irq_data_fifo_data_valid;
  /* ni/irq_fifo.vhd:113:29  */
  assign n1443_o = n1442_o ? irq_w_ptr : data_w_ptr;
  /* ni/irq_fifo.vhd:123:42  */
  assign n1446_o = n1403_o[14];
  /* ni/irq_fifo.vhd:123:31  */
  assign n1447_o = sel & n1446_o;
  /* ni/irq_fifo.vhd:125:35  */
  assign n1448_o = n1403_o[15];
  /* ni/irq_fifo.vhd:125:38  */
  assign n1449_o = ~n1448_o;
  /* ni/irq_fifo.vhd:126:50  */
  assign n1450_o = n1403_o[10:0];
  /* ni/irq_fifo.vhd:128:11  */
  assign n1452_o = n1450_o == 11'b00000000000;
  /* ni/irq_fifo.vhd:132:11  */
  assign n1454_o = n1450_o == 11'b00000000001;
  assign n1455_o = {n1454_o, n1452_o};
  /* ni/irq_fifo.vhd:126:33  */
  always @*
    case (n1455_o)
      2'b10: n1458_o <= 1'b0;
      2'b01: n1458_o <= 1'b0;
      default: n1458_o <= 1'b1;
    endcase
  /* ni/irq_fifo.vhd:126:33  */
  always @*
    case (n1455_o)
      2'b10: n1461_o <= 1'b0;
      2'b01: n1461_o <= 1'b1;
      default: n1461_o <= 1'b0;
    endcase
  /* ni/irq_fifo.vhd:126:33  */
  always @*
    case (n1455_o)
      2'b10: n1464_o <= 1'b1;
      2'b01: n1464_o <= 1'b0;
      default: n1464_o <= 1'b0;
    endcase
  /* ni/irq_fifo.vhd:126:33  */
  always @*
    case (n1455_o)
      2'b10: n1465_o <= data_r_ptr;
      2'b01: n1465_o <= irq_r_ptr;
      default: n1465_o <= data_r_ptr;
    endcase
  /* ni/irq_fifo.vhd:125:25  */
  assign n1467_o = n1449_o ? n1458_o : 1'b1;
  /* ni/irq_fifo.vhd:125:25  */
  assign n1469_o = n1449_o ? n1461_o : 1'b0;
  /* ni/irq_fifo.vhd:125:25  */
  assign n1471_o = n1449_o ? n1464_o : 1'b0;
  /* ni/irq_fifo.vhd:123:17  */
  assign n1472_o = n1482_o ? n1465_o : data_r_ptr;
  /* ni/irq_fifo.vhd:123:17  */
  assign n1474_o = n1447_o ? n1467_o : 1'b0;
  /* ni/irq_fifo.vhd:123:17  */
  assign n1477_o = n1447_o ? n1469_o : 1'b0;
  /* ni/irq_fifo.vhd:123:17  */
  assign n1480_o = n1447_o ? n1471_o : 1'b0;
  /* ni/irq_fifo.vhd:123:17  */
  assign n1482_o = n1447_o & n1449_o;
  /* ni/irq_fifo.vhd:154:60  */
  assign n1484_o = irq_irq_fifo_data_valid & irq_not_full;
  /* ni/irq_fifo.vhd:154:108  */
  assign n1485_o = irq_data_fifo_data_valid & data_not_full;
  /* ni/irq_fifo.vhd:154:79  */
  assign n1486_o = n1484_o | n1485_o;
  /* ni/irq_fifo.vhd:164:35  */
  assign tdpram_n1490 = tdpram_b_dout; // (signal)
  /* ni/irq_fifo.vhd:146:9  */
  tdp_ram_14_5 tdpram (
    .a_clk(clk),
    .a_wr(n1486_o),
    .a_addr(w_ptr),
    .a_din(w_data),
    .b_clk(clk),
    .b_wr(n1488_o),
    .b_addr(r_ptr),
    .b_din(n1489_o),
    .a_dout(),
    .b_dout(tdpram_b_dout));
  /* ni/irq_fifo.vhd:173:57  */
  assign n1497_o = irq_irq_fifo_data_valid & irq_not_full;
  /* ni/irq_fifo.vhd:174:47  */
  assign n1499_o = irq_w_ptr == 5'b01111;
  /* ni/irq_fifo.vhd:177:64  */
  assign n1501_o = irq_w_ptr + 5'b00001;
  /* ni/irq_fifo.vhd:174:33  */
  assign n1503_o = n1499_o ? 5'b00000 : n1501_o;
  /* ni/irq_fifo.vhd:173:25  */
  assign n1504_o = n1497_o ? n1503_o : irq_w_ptr;
  /* ni/irq_fifo.vhd:171:25  */
  assign n1506_o = reset ? 5'b00000 : n1504_o;
  /* ni/irq_fifo.vhd:170:17  */
  always @(posedge clk)
    n1509_q <= n1506_o;
  /* ni/irq_fifo.vhd:189:58  */
  assign n1513_o = irq_data_fifo_data_valid & data_not_full;
  /* ni/irq_fifo.vhd:190:48  */
  assign n1515_o = data_w_ptr == 5'b10000;
  /* ni/irq_fifo.vhd:193:66  */
  assign n1517_o = data_w_ptr - 5'b00001;
  /* ni/irq_fifo.vhd:190:33  */
  assign n1519_o = n1515_o ? 5'b11111 : n1517_o;
  /* ni/irq_fifo.vhd:189:25  */
  assign n1520_o = n1513_o ? n1519_o : data_w_ptr;
  /* ni/irq_fifo.vhd:187:25  */
  assign n1522_o = reset ? 5'b11111 : n1520_o;
  /* ni/irq_fifo.vhd:186:17  */
  always @(posedge clk)
    n1525_q <= n1522_o;
  /* ni/irq_fifo.vhd:205:49  */
  assign n1529_o = irq_read & irq_not_empty;
  /* ni/irq_fifo.vhd:206:47  */
  assign n1531_o = irq_r_ptr == 5'b01111;
  /* ni/irq_fifo.vhd:209:64  */
  assign n1533_o = irq_r_ptr + 5'b00001;
  /* ni/irq_fifo.vhd:206:33  */
  assign n1535_o = n1531_o ? 5'b00000 : n1533_o;
  /* ni/irq_fifo.vhd:205:25  */
  assign n1536_o = n1529_o ? n1535_o : irq_r_ptr;
  /* ni/irq_fifo.vhd:203:25  */
  assign n1538_o = reset ? 5'b00000 : n1536_o;
  /* ni/irq_fifo.vhd:202:17  */
  always @(posedge clk)
    n1541_q <= n1538_o;
  /* ni/irq_fifo.vhd:221:50  */
  assign n1545_o = data_read & data_not_empty;
  /* ni/irq_fifo.vhd:222:48  */
  assign n1547_o = data_r_ptr == 5'b10000;
  /* ni/irq_fifo.vhd:225:66  */
  assign n1549_o = data_r_ptr - 5'b00001;
  /* ni/irq_fifo.vhd:222:33  */
  assign n1551_o = n1547_o ? 5'b11111 : n1549_o;
  /* ni/irq_fifo.vhd:221:25  */
  assign n1552_o = n1545_o ? n1551_o : data_r_ptr;
  /* ni/irq_fifo.vhd:219:25  */
  assign n1554_o = reset ? 5'b11111 : n1552_o;
  /* ni/irq_fifo.vhd:218:17  */
  always @(posedge clk)
    n1557_q <= n1554_o;
  /* ni/irq_fifo.vhd:234:25  */
  assign n1562_o = reset ? 1'b0 : next_error;
  /* ni/irq_fifo.vhd:233:17  */
  always @(posedge clk)
    n1566_q <= n1562_o;
  /* ni/irq_fifo.vhd:233:17  */
  assign n1567_o = {n1566_q, 18'b000000000000000000, tdpram_n1490};
endmodule

module rx_unit
  (input  clk,
   input  reset,
   input  [34:0] pkt_in,
   output [13:0] spm_addr,
   output [1:0] spm_en,
   output spm_wr,
   output [63:0] spm_wdata,
   output [13:0] config_addr,
   output config_en,
   output config_wr,
   output [31:0] config_wdata,
   output [13:0] irq_fifo_data,
   output irq_fifo_data_valid,
   output irq_fifo_irq_valid);
  wire [13:0] n1213_o;
  wire [1:0] n1214_o;
  wire n1215_o;
  wire [63:0] n1216_o;
  wire [13:0] n1218_o;
  wire n1219_o;
  wire n1220_o;
  wire [31:0] n1221_o;
  wire new_pkt;
  wire new_data_pkt;
  wire new_config_pkt;
  wire new_irq_pkt;
  wire wdata_high_en;
  wire addr_load;
  wire lst_data_pkt;
  wire [13:0] addr;
  wire [13:0] next_addr;
  wire [13:0] int_addr;
  wire [13:0] next_int_addr;
  wire [31:0] wdata_high;
  wire [2:0] state;
  wire [2:0] next_state;
  wire n1225_o;
  wire n1226_o;
  wire n1227_o;
  wire n1228_o;
  wire n1229_o;
  wire n1230_o;
  wire n1231_o;
  wire n1232_o;
  wire n1233_o;
  wire n1234_o;
  wire n1235_o;
  wire n1236_o;
  wire n1237_o;
  wire n1238_o;
  wire n1239_o;
  wire n1240_o;
  wire n1241_o;
  wire n1242_o;
  wire [31:0] n1243_o;
  wire [31:0] n1244_o;
  wire n1245_o;
  wire n1246_o;
  localparam [1:0] n1249_o = 2'b00;
  wire [13:0] n1254_o;
  wire [13:0] n1255_o;
  wire [2:0] n1257_o;
  wire [2:0] n1259_o;
  wire [2:0] n1261_o;
  wire n1263_o;
  wire [13:0] n1265_o;
  wire n1266_o;
  wire n1267_o;
  wire [31:0] n1270_o;
  wire n1271_o;
  wire n1272_o;
  wire n1273_o;
  wire [31:0] n1274_o;
  wire n1277_o;
  wire [2:0] n1280_o;
  wire n1282_o;
  localparam [1:0] n1283_o = 2'b11;
  wire n1285_o;
  wire n1286_o;
  wire [2:0] n1289_o;
  wire n1291_o;
  wire n1294_o;
  wire n1295_o;
  wire [2:0] n1298_o;
  wire n1300_o;
  wire n1304_o;
  wire [31:0] n1307_o;
  wire n1309_o;
  wire [5:0] n1310_o;
  wire n1311_o;
  wire n1312_o;
  reg n1314_o;
  wire n1315_o;
  wire n1316_o;
  reg n1318_o;
  reg n1320_o;
  reg [31:0] n1322_o;
  reg n1325_o;
  reg n1327_o;
  reg [13:0] n1329_o;
  reg n1333_o;
  reg n1337_o;
  reg n1342_o;
  reg [13:0] n1345_o;
  reg [13:0] n1347_o;
  reg [2:0] n1351_o;
  wire [13:0] n1357_o;
  wire [13:0] n1358_o;
  reg [13:0] n1361_q;
  wire [31:0] n1365_o;
  wire [31:0] n1369_o;
  reg [31:0] n1370_q;
  wire [13:0] n1375_o;
  wire [2:0] n1377_o;
  reg [13:0] n1381_q;
  reg [2:0] n1382_q;
  wire n1386_o;
  wire n1387_o;
  wire n1388_o;
  wire n1389_o;
  wire n1390_o;
  wire n1391_o;
  wire n1392_o;
  wire n1393_o;
  wire n1395_o;
  wire n1397_o;
  reg n1400_q;
  wire [80:0] n1401_o;
  wire [47:0] n1402_o;
  assign spm_addr = n1213_o;
  assign spm_en = n1214_o;
  assign spm_wr = n1215_o;
  assign spm_wdata = n1216_o;
  assign config_addr = n1218_o;
  assign config_en = n1219_o;
  assign config_wr = n1220_o;
  assign config_wdata = n1221_o;
  assign irq_fifo_data = n1329_o;
  assign irq_fifo_data_valid = n1246_o;
  assign irq_fifo_irq_valid = n1333_o;
  /* ni/packet_manager.vhd:323:16  */
  assign n1213_o = n1401_o[13:0];
  /* ni/packet_manager.vhd:318:16  */
  assign n1214_o = n1401_o[15:14];
  /* ni/packet_manager.vhd:60:5  */
  assign n1215_o = n1401_o[16];
  /* ni/packet_manager.vhd:51:5  */
  assign n1216_o = n1401_o[80:17];
  assign n1218_o = n1402_o[13:0];
  /* ni/packet_manager.vhd:399:1  */
  assign n1219_o = n1402_o[14];
  assign n1220_o = n1402_o[15];
  /* ni/packet_manager.vhd:387:1  */
  assign n1221_o = n1402_o[47:16];
  /* ni/rx_unit.vhd:63:16  */
  assign new_pkt = n1230_o; // (signal)
  /* ni/rx_unit.vhd:63:25  */
  assign new_data_pkt = n1233_o; // (signal)
  /* ni/rx_unit.vhd:63:39  */
  assign new_config_pkt = n1238_o; // (signal)
  /* ni/rx_unit.vhd:63:55  */
  assign new_irq_pkt = n1242_o; // (signal)
  /* ni/rx_unit.vhd:64:16  */
  assign wdata_high_en = n1337_o; // (signal)
  /* ni/rx_unit.vhd:64:45  */
  assign addr_load = n1342_o; // (signal)
  /* ni/rx_unit.vhd:64:56  */
  assign lst_data_pkt = n1400_q; // (signal)
  /* ni/rx_unit.vhd:65:16  */
  assign addr = n1361_q; // (signal)
  /* ni/rx_unit.vhd:65:22  */
  assign next_addr = n1345_o; // (signal)
  /* ni/rx_unit.vhd:65:33  */
  assign int_addr = n1381_q; // (signal)
  /* ni/rx_unit.vhd:65:43  */
  assign next_int_addr = n1347_o; // (signal)
  /* ni/rx_unit.vhd:67:8  */
  assign wdata_high = n1370_q; // (signal)
  /* ni/rx_unit.vhd:71:16  */
  assign state = n1382_q; // (signal)
  /* ni/rx_unit.vhd:71:23  */
  assign next_state = n1351_o; // (signal)
  /* ni/rx_unit.vhd:75:26  */
  assign n1225_o = pkt_in[34];
  /* ni/rx_unit.vhd:75:53  */
  assign n1226_o = pkt_in[33];
  /* ni/rx_unit.vhd:75:43  */
  assign n1227_o = n1225_o & n1226_o;
  /* ni/rx_unit.vhd:75:85  */
  assign n1228_o = pkt_in[32];
  /* ni/rx_unit.vhd:75:75  */
  assign n1229_o = ~n1228_o;
  /* ni/rx_unit.vhd:75:70  */
  assign n1230_o = n1227_o & n1229_o;
  /* ni/rx_unit.vhd:78:48  */
  assign n1231_o = pkt_in[30];
  /* ni/rx_unit.vhd:78:38  */
  assign n1232_o = ~n1231_o;
  /* ni/rx_unit.vhd:78:33  */
  assign n1233_o = new_pkt & n1232_o;
  /* ni/rx_unit.vhd:81:49  */
  assign n1234_o = pkt_in[31];
  /* ni/rx_unit.vhd:81:39  */
  assign n1235_o = ~n1234_o;
  /* ni/rx_unit.vhd:81:35  */
  assign n1236_o = new_pkt & n1235_o;
  /* ni/rx_unit.vhd:81:106  */
  assign n1237_o = pkt_in[30];
  /* ni/rx_unit.vhd:81:96  */
  assign n1238_o = n1236_o & n1237_o;
  /* ni/rx_unit.vhd:84:42  */
  assign n1239_o = pkt_in[31];
  /* ni/rx_unit.vhd:84:32  */
  assign n1240_o = new_pkt & n1239_o;
  /* ni/rx_unit.vhd:84:98  */
  assign n1241_o = pkt_in[30];
  /* ni/rx_unit.vhd:84:88  */
  assign n1242_o = n1240_o & n1241_o;
  /* ni/rx_unit.vhd:87:62  */
  assign n1243_o = pkt_in[31:0];
  /* ni/rx_unit.vhd:89:65  */
  assign n1244_o = pkt_in[31:0];
  /* ni/rx_unit.vhd:96:55  */
  assign n1245_o = pkt_in[32];
  /* ni/rx_unit.vhd:96:45  */
  assign n1246_o = lst_data_pkt & n1245_o;
  /* ni/rx_unit.vhd:113:43  */
  assign n1254_o = int_addr + 14'b00000000000001;
  /* ni/rx_unit.vhd:117:65  */
  assign n1255_o = pkt_in[29:16];
  /* ni/rx_unit.vhd:122:33  */
  assign n1257_o = new_irq_pkt ? 3'b101 : state;
  /* ni/rx_unit.vhd:120:33  */
  assign n1259_o = new_config_pkt ? 3'b100 : n1257_o;
  /* ni/rx_unit.vhd:118:33  */
  assign n1261_o = new_data_pkt ? 3'b010 : n1259_o;
  /* ni/rx_unit.vhd:115:25  */
  assign n1263_o = state == 3'b000;
  /* ni/rx_unit.vhd:127:55  */
  assign n1265_o = addr + 14'b00000000000001;
  /* ni/rx_unit.vhd:128:43  */
  assign n1266_o = pkt_in[32];
  /* ni/rx_unit.vhd:128:60  */
  assign n1267_o = ~n1266_o;
  /* ni/rx_unit.vhd:134:107  */
  assign n1270_o = pkt_in[31:0];
  assign n1271_o = n1249_o[0];
  /* ni/rx_unit.vhd:128:33  */
  assign n1272_o = n1267_o ? n1271_o : 1'b1;
  /* ni/rx_unit.vhd:128:33  */
  assign n1273_o = n1267_o ? 1'b0 : 1'b1;
  /* ni/rx_unit.vhd:128:33  */
  assign n1274_o = n1267_o ? wdata_high : n1270_o;
  /* ni/rx_unit.vhd:128:33  */
  assign n1277_o = n1267_o ? 1'b1 : 1'b0;
  /* ni/rx_unit.vhd:128:33  */
  assign n1280_o = n1267_o ? 3'b001 : 3'b000;
  /* ni/rx_unit.vhd:126:25  */
  assign n1282_o = state == 3'b010;
  /* ni/rx_unit.vhd:143:43  */
  assign n1285_o = pkt_in[32];
  /* ni/rx_unit.vhd:143:60  */
  assign n1286_o = ~n1285_o;
  /* ni/rx_unit.vhd:143:33  */
  assign n1289_o = n1286_o ? 3'b010 : 3'b000;
  /* ni/rx_unit.vhd:138:25  */
  assign n1291_o = state == 3'b001;
  /* ni/rx_unit.vhd:153:43  */
  assign n1294_o = pkt_in[32];
  /* ni/rx_unit.vhd:153:60  */
  assign n1295_o = ~n1294_o;
  /* ni/rx_unit.vhd:153:33  */
  assign n1298_o = n1295_o ? 3'b011 : 3'b000;
  /* ni/rx_unit.vhd:150:25  */
  assign n1300_o = state == 3'b100;
  /* ni/rx_unit.vhd:159:25  */
  assign n1304_o = state == 3'b011;
  /* ni/rx_unit.vhd:169:99  */
  assign n1307_o = pkt_in[31:0];
  /* ni/rx_unit.vhd:165:25  */
  assign n1309_o = state == 3'b101;
  assign n1310_o = {n1309_o, n1304_o, n1300_o, n1291_o, n1282_o, n1263_o};
  assign n1311_o = n1283_o[0];
  assign n1312_o = n1249_o[0];
  /* ni/rx_unit.vhd:114:17  */
  always @*
    case (n1310_o)
      6'b100000: n1314_o <= 1'b1;
      6'b010000: n1314_o <= n1312_o;
      6'b001000: n1314_o <= n1312_o;
      6'b000100: n1314_o <= n1311_o;
      6'b000010: n1314_o <= n1272_o;
      6'b000001: n1314_o <= n1312_o;
      default: n1314_o <= 1'bX;
    endcase
  assign n1315_o = n1283_o[1];
  assign n1316_o = n1249_o[1];
  /* ni/rx_unit.vhd:114:17  */
  always @*
    case (n1310_o)
      6'b100000: n1318_o <= n1316_o;
      6'b010000: n1318_o <= n1316_o;
      6'b001000: n1318_o <= n1316_o;
      6'b000100: n1318_o <= n1315_o;
      6'b000010: n1318_o <= n1316_o;
      6'b000001: n1318_o <= n1316_o;
      default: n1318_o <= 1'bX;
    endcase
  /* ni/rx_unit.vhd:114:17  */
  always @*
    case (n1310_o)
      6'b100000: n1320_o <= 1'b1;
      6'b010000: n1320_o <= 1'b0;
      6'b001000: n1320_o <= 1'b0;
      6'b000100: n1320_o <= 1'b1;
      6'b000010: n1320_o <= n1273_o;
      6'b000001: n1320_o <= 1'b0;
      default: n1320_o <= 1'bX;
    endcase
  /* ni/rx_unit.vhd:114:17  */
  always @*
    case (n1310_o)
      6'b100000: n1322_o <= n1307_o;
      6'b010000: n1322_o <= wdata_high;
      6'b001000: n1322_o <= wdata_high;
      6'b000100: n1322_o <= wdata_high;
      6'b000010: n1322_o <= n1274_o;
      6'b000001: n1322_o <= wdata_high;
      default: n1322_o <= 32'bX;
    endcase
  /* ni/rx_unit.vhd:114:17  */
  always @*
    case (n1310_o)
      6'b100000: n1325_o <= 1'b0;
      6'b010000: n1325_o <= 1'b1;
      6'b001000: n1325_o <= 1'b1;
      6'b000100: n1325_o <= 1'b0;
      6'b000010: n1325_o <= 1'b0;
      6'b000001: n1325_o <= 1'b0;
      default: n1325_o <= 1'bX;
    endcase
  /* ni/rx_unit.vhd:114:17  */
  always @*
    case (n1310_o)
      6'b100000: n1327_o <= 1'b0;
      6'b010000: n1327_o <= 1'b1;
      6'b001000: n1327_o <= 1'b1;
      6'b000100: n1327_o <= 1'b0;
      6'b000010: n1327_o <= 1'b0;
      6'b000001: n1327_o <= 1'b0;
      default: n1327_o <= 1'bX;
    endcase
  /* ni/rx_unit.vhd:114:17  */
  always @*
    case (n1310_o)
      6'b100000: n1329_o <= addr;
      6'b010000: n1329_o <= addr;
      6'b001000: n1329_o <= addr;
      6'b000100: n1329_o <= int_addr;
      6'b000010: n1329_o <= addr;
      6'b000001: n1329_o <= addr;
      default: n1329_o <= 14'bX;
    endcase
  /* ni/rx_unit.vhd:114:17  */
  always @*
    case (n1310_o)
      6'b100000: n1333_o <= 1'b1;
      6'b010000: n1333_o <= 1'b0;
      6'b001000: n1333_o <= 1'b0;
      6'b000100: n1333_o <= 1'b0;
      6'b000010: n1333_o <= 1'b0;
      6'b000001: n1333_o <= 1'b0;
      default: n1333_o <= 1'bX;
    endcase
  /* ni/rx_unit.vhd:114:17  */
  always @*
    case (n1310_o)
      6'b100000: n1337_o <= 1'b0;
      6'b010000: n1337_o <= 1'b0;
      6'b001000: n1337_o <= 1'b0;
      6'b000100: n1337_o <= 1'b0;
      6'b000010: n1337_o <= n1277_o;
      6'b000001: n1337_o <= 1'b0;
      default: n1337_o <= 1'bX;
    endcase
  /* ni/rx_unit.vhd:114:17  */
  always @*
    case (n1310_o)
      6'b100000: n1342_o <= 1'b0;
      6'b010000: n1342_o <= 1'b0;
      6'b001000: n1342_o <= 1'b0;
      6'b000100: n1342_o <= 1'b0;
      6'b000010: n1342_o <= 1'b0;
      6'b000001: n1342_o <= 1'b1;
      default: n1342_o <= 1'bX;
    endcase
  /* ni/rx_unit.vhd:114:17  */
  always @*
    case (n1310_o)
      6'b100000: n1345_o <= addr;
      6'b010000: n1345_o <= addr;
      6'b001000: n1345_o <= addr;
      6'b000100: n1345_o <= next_int_addr;
      6'b000010: n1345_o <= addr;
      6'b000001: n1345_o <= addr;
      default: n1345_o <= 14'bX;
    endcase
  /* ni/rx_unit.vhd:114:17  */
  always @*
    case (n1310_o)
      6'b100000: n1347_o <= n1254_o;
      6'b010000: n1347_o <= n1254_o;
      6'b001000: n1347_o <= n1254_o;
      6'b000100: n1347_o <= n1254_o;
      6'b000010: n1347_o <= n1265_o;
      6'b000001: n1347_o <= n1255_o;
      default: n1347_o <= 14'bX;
    endcase
  /* ni/rx_unit.vhd:114:17  */
  always @*
    case (n1310_o)
      6'b100000: n1351_o <= 3'b000;
      6'b010000: n1351_o <= 3'b000;
      6'b001000: n1351_o <= n1298_o;
      6'b000100: n1351_o <= n1289_o;
      6'b000010: n1351_o <= n1280_o;
      6'b000001: n1351_o <= n1261_o;
      default: n1351_o <= 3'bX;
    endcase
  /* ni/rx_unit.vhd:180:56  */
  assign n1357_o = pkt_in[29:16];
  /* ni/rx_unit.vhd:179:25  */
  assign n1358_o = addr_load ? n1357_o : next_addr;
  /* ni/rx_unit.vhd:178:17  */
  always @(posedge clk)
    n1361_q <= n1358_o;
  /* ni/rx_unit.vhd:192:62  */
  assign n1365_o = pkt_in[31:0];
  /* ni/rx_unit.vhd:190:17  */
  assign n1369_o = wdata_high_en ? n1365_o : wdata_high;
  /* ni/rx_unit.vhd:190:17  */
  always @(posedge clk)
    n1370_q <= n1369_o;
  /* ni/rx_unit.vhd:201:25  */
  assign n1375_o = reset ? 14'b00000000000000 : next_int_addr;
  /* ni/rx_unit.vhd:201:25  */
  assign n1377_o = reset ? 3'b000 : next_state;
  /* ni/rx_unit.vhd:200:17  */
  always @(posedge clk)
    n1381_q <= n1375_o;
  /* ni/rx_unit.vhd:200:17  */
  always @(posedge clk)
    n1382_q <= n1377_o;
  /* ni/rx_unit.vhd:217:77  */
  assign n1386_o = pkt_in[31];
  /* ni/rx_unit.vhd:217:67  */
  assign n1387_o = new_data_pkt & n1386_o;
  /* ni/rx_unit.vhd:217:49  */
  assign n1388_o = ~n1387_o;
  /* ni/rx_unit.vhd:217:135  */
  assign n1389_o = pkt_in[32];
  /* ni/rx_unit.vhd:217:125  */
  assign n1390_o = n1388_o & n1389_o;
  /* ni/rx_unit.vhd:217:43  */
  assign n1391_o = reset | n1390_o;
  /* ni/rx_unit.vhd:219:56  */
  assign n1392_o = pkt_in[31];
  /* ni/rx_unit.vhd:219:46  */
  assign n1393_o = new_data_pkt & n1392_o;
  /* ni/rx_unit.vhd:219:25  */
  assign n1395_o = n1393_o ? 1'b1 : lst_data_pkt;
  /* ni/rx_unit.vhd:217:25  */
  assign n1397_o = n1391_o ? 1'b0 : n1395_o;
  /* ni/rx_unit.vhd:216:17  */
  always @(posedge clk)
    n1400_q <= n1397_o;
  /* ni/rx_unit.vhd:216:17  */
  assign n1401_o = {n1322_o, n1243_o, n1320_o, n1318_o, n1314_o, addr};
  assign n1402_o = {n1244_o, n1327_o, n1325_o, int_addr};
endmodule

module packet_manager
  (input  clk,
   input  reset,
   input  [13:0] config_addr,
   input  config_en,
   input  config_wr,
   input  [31:0] config_wdata,
   input  sel,
   input  [63:0] spm_slv_rdata,
   input  spm_slv_error,
   input  [5:0] dma_num,
   input  dma_en,
   input  [15:0] route,
   input  mc,
   input  [1:0] mc_idx,
   input  [1:0] mc_p,
   input  [3:0] pkt_len,
   output [31:0] config_slv_rdata,
   output config_slv_error,
   output [13:0] spm_addr,
   output [1:0] spm_en,
   output spm_wr,
   output [63:0] spm_wdata,
   output [34:0] pkt_out);
  wire [47:0] n855_o;
  wire [31:0] n857_o;
  wire n858_o;
  wire [13:0] n860_o;
  wire [1:0] n861_o;
  wire n862_o;
  wire [63:0] n863_o;
  wire [64:0] n864_o;
  wire [2:0] state;
  wire [2:0] next_state;
  wire [44:0] dmatbl_data;
  wire [13:0] count_reg;
  wire [13:0] count_next;
  wire [1:0] pkt_type;
  wire dma_en_reg;
  wire [13:0] read_ptr_reg;
  wire [13:0] read_ptr_next;
  wire hi_lo_next;
  wire hi_lo_reg;
  wire port_b_wr;
  wire [5:0] port_b_addr;
  wire [44:0] port_b_din;
  wire [44:0] port_b_dout;
  wire [5:0] dma_num_reg;
  wire dma_update_en;
  wire [5:0] dma_update_addr;
  wire [44:0] dma_update_data;
  wire port_a_wr_hi;
  wire port_a_wr_lo;
  wire [5:0] port_a_addr;
  wire [44:0] port_a_din;
  wire [44:0] port_a_dout;
  wire config_slv_error_next;
  wire [3:0] pkt_len_reg;
  wire [3:0] pkt_len_next;
  wire [15:0] route_reg;
  wire [31:0] payload_data;
  wire [31:0] payload_data_next;
  wire [13:0] n872_o;
  wire [3:0] n873_o;
  wire [1:0] n874_o;
  wire n876_o;
  wire [1:0] n878_o;
  wire [4:0] n880_o;
  wire [7:0] n882_o;
  wire [18:0] n884_o;
  wire [34:0] n885_o;
  wire n886_o;
  wire [13:0] n888_o;
  wire [13:0] n889_o;
  wire [13:0] n890_o;
  wire [13:0] n892_o;
  wire [13:0] n893_o;
  wire [13:0] n894_o;
  wire n895_o;
  wire [1:0] n896_o;
  wire n898_o;
  wire [1:0] n900_o;
  wire n902_o;
  wire n903_o;
  wire [13:0] n904_o;
  wire [13:0] n905_o;
  wire [13:0] n906_o;
  wire [13:0] n907_o;
  wire [13:0] n908_o;
  wire [13:0] n909_o;
  wire [13:0] n910_o;
  wire [13:0] n911_o;
  wire [13:0] n912_o;
  wire [1:0] n913_o;
  wire n915_o;
  wire [3:0] n916_o;
  wire [3:0] n917_o;
  wire [3:0] n918_o;
  wire [9:0] n919_o;
  wire [3:0] n921_o;
  wire [4:0] n923_o;
  wire [13:0] n924_o;
  wire [18:0] n925_o;
  wire [34:0] n926_o;
  wire [15:0] n927_o;
  wire [15:0] n928_o;
  wire [15:0] n929_o;
  wire [34:0] n931_o;
  wire [2:0] n933_o;
  wire [13:0] n934_o;
  wire n935_o;
  wire [13:0] n936_o;
  wire n939_o;
  wire [13:0] n940_o;
  wire [28:0] n941_o;
  wire [13:0] n942_o;
  wire [13:0] n943_o;
  wire [27:0] n944_o;
  wire [28:0] n945_o;
  wire [28:0] n946_o;
  wire [3:0] n947_o;
  wire [15:0] n948_o;
  wire [15:0] n949_o;
  wire [34:0] n950_o;
  wire [2:0] n952_o;
  wire [13:0] n953_o;
  wire [1:0] n954_o;
  wire [13:0] n955_o;
  wire n957_o;
  wire [13:0] n958_o;
  wire [13:0] n959_o;
  wire [27:0] n960_o;
  wire [28:0] n961_o;
  wire [28:0] n962_o;
  wire [3:0] n963_o;
  wire [1:0] n965_o;
  wire [1:0] n967_o;
  wire [15:0] n968_o;
  wire [15:0] n969_o;
  wire [34:0] n971_o;
  wire [2:0] n972_o;
  wire [13:0] n973_o;
  wire [1:0] n974_o;
  wire [13:0] n975_o;
  wire n977_o;
  wire [13:0] n978_o;
  wire [13:0] n979_o;
  wire [27:0] n980_o;
  wire [28:0] n981_o;
  wire [28:0] n982_o;
  wire [3:0] n983_o;
  wire [1:0] n985_o;
  wire [1:0] n987_o;
  wire n989_o;
  wire [31:0] n990_o;
  wire [3:0] n992_o;
  wire [13:0] n994_o;
  wire n996_o;
  wire n998_o;
  wire n999_o;
  wire [31:0] n1000_o;
  wire [34:0] n1002_o;
  wire [13:0] n1004_o;
  wire [31:0] n1005_o;
  wire [34:0] n1007_o;
  wire [34:0] n1008_o;
  wire [2:0] n1011_o;
  wire [13:0] n1012_o;
  wire n1014_o;
  wire [3:0] n1016_o;
  wire [13:0] n1018_o;
  wire n1020_o;
  wire n1022_o;
  wire n1023_o;
  wire [34:0] n1025_o;
  wire [13:0] n1028_o;
  wire [34:0] n1030_o;
  wire [15:0] n1031_o;
  wire [15:0] n1032_o;
  wire [15:0] n1033_o;
  wire [34:0] n1034_o;
  wire [2:0] n1037_o;
  wire [13:0] n1038_o;
  wire n1040_o;
  wire [34:0] n1042_o;
  wire n1044_o;
  wire [34:0] n1046_o;
  wire n1048_o;
  wire [4:0] n1049_o;
  wire [15:0] n1050_o;
  reg [15:0] n1052_o;
  reg [34:0] n1054_o;
  reg [2:0] n1059_o;
  reg [13:0] n1061_o;
  reg [1:0] n1063_o;
  reg [13:0] n1065_o;
  reg n1068_o;
  wire [13:0] n1070_o;
  reg [13:0] n1072_o;
  wire [27:0] n1073_o;
  wire [28:0] n1074_o;
  reg [28:0] n1076_o;
  wire [1:0] n1078_o;
  reg [3:0] n1080_o;
  wire [1:0] n1081_o;
  reg [1:0] n1084_o;
  wire [13:0] n1085_o;
  reg [13:0] n1088_o;
  wire [1:0] n1089_o;
  reg [1:0] n1092_o;
  wire [13:0] n1093_o;
  reg [13:0] n1096_o;
  wire [5:0] n1103_o;
  localparam [31:0] n1104_o = 32'b00000000000000000000000000000000;
  wire n1105_o;
  wire [27:0] n1106_o;
  wire [15:0] n1107_o;
  wire n1108_o;
  wire n1109_o;
  wire n1110_o;
  wire n1111_o;
  wire n1112_o;
  wire n1113_o;
  wire n1114_o;
  wire n1116_o;
  wire n1118_o;
  wire n1121_o;
  wire n1123_o;
  wire n1124_o;
  wire [27:0] n1125_o;
  wire [15:0] n1126_o;
  wire [15:0] n1127_o;
  wire [15:0] n1128_o;
  wire [11:0] n1129_o;
  wire [11:0] n1130_o;
  wire [11:0] n1131_o;
  wire n1132_o;
  wire n1133_o;
  wire [2:0] n1136_o;
  wire n1140_o;
  wire [5:0] n1141_o;
  wire [28:0] dmatbl1_a_dout;
  wire [28:0] dmatbl1_b_dout;
  wire [28:0] n1143_o;
  wire [28:0] n1145_o;
  wire [15:0] dmatbl2_a_dout;
  wire [15:0] dmatbl2_b_dout;
  wire [15:0] n1147_o;
  wire [15:0] n1149_o;
  wire [3:0] n1152_o;
  wire n1154_o;
  wire n1155_o;
  wire n1158_o;
  wire n1164_o;
  reg n1167_q;
  wire n1171_o;
  reg n1174_q;
  wire n1178_o;
  reg n1182_q;
  wire [2:0] n1186_o;
  reg [2:0] n1189_q;
  reg [13:0] n1199_q;
  reg [13:0] n1200_q;
  reg [5:0] n1201_q;
  reg [3:0] n1202_q;
  reg [15:0] n1203_q;
  reg [31:0] n1204_q;
  wire [44:0] n1205_o;
  wire [44:0] n1206_o;
  wire [44:0] n1207_o;
  wire [44:0] n1208_o;
  wire [31:0] n1209_o;
  wire [32:0] n1210_o;
  wire [80:0] n1211_o;
  assign config_slv_rdata = n857_o;
  assign config_slv_error = n858_o;
  assign spm_addr = n860_o;
  assign spm_en = n861_o;
  assign spm_wr = n862_o;
  assign spm_wdata = n863_o;
  assign pkt_out = n1054_o;
  /* ni/schedule_table.vhd:103:16  */
  assign n855_o = {config_wdata, config_wr, config_en, config_addr};
  /* ni/schedule_table.vhd:59:5  */
  assign n857_o = n1210_o[31:0];
  /* ni/schedule_table.vhd:58:5  */
  assign n858_o = n1210_o[32];
  /* ni/schedule_table.vhd:56:5  */
  assign n860_o = n1211_o[13:0];
  /* ni/schedule_table.vhd:51:5  */
  assign n861_o = n1211_o[15:14];
  assign n862_o = n1211_o[16];
  assign n863_o = n1211_o[80:17];
  /* ni/schedule_table.vhd:190:1  */
  assign n864_o = {spm_slv_error, spm_slv_rdata};
  /* ni/packet_manager.vhd:78:8  */
  assign state = n1189_q; // (signal)
  /* ni/packet_manager.vhd:78:15  */
  assign next_state = n1059_o; // (signal)
  /* ni/packet_manager.vhd:83:8  */
  assign dmatbl_data = port_b_dout; // (signal)
  /* ni/packet_manager.vhd:94:8  */
  assign count_reg = n1199_q; // (signal)
  /* ni/packet_manager.vhd:94:19  */
  assign count_next = n1061_o; // (signal)
  /* ni/packet_manager.vhd:101:8  */
  assign pkt_type = n1063_o; // (signal)
  /* ni/packet_manager.vhd:103:8  */
  assign dma_en_reg = n1167_q; // (signal)
  /* ni/packet_manager.vhd:105:8  */
  assign read_ptr_reg = n1200_q; // (signal)
  /* ni/packet_manager.vhd:105:22  */
  assign read_ptr_next = n1065_o; // (signal)
  /* ni/packet_manager.vhd:107:8  */
  assign hi_lo_next = n1123_o; // (signal)
  /* ni/packet_manager.vhd:108:8  */
  assign hi_lo_reg = n1174_q; // (signal)
  /* ni/packet_manager.vhd:110:8  */
  assign port_b_wr = n1140_o; // (signal)
  /* ni/packet_manager.vhd:111:8  */
  assign port_b_addr = n1141_o; // (signal)
  /* ni/packet_manager.vhd:112:8  */
  assign port_b_din = dma_update_data; // (signal)
  /* ni/packet_manager.vhd:113:8  */
  assign port_b_dout = n1205_o; // (signal)
  /* ni/packet_manager.vhd:115:8  */
  assign dma_num_reg = n1201_q; // (signal)
  /* ni/packet_manager.vhd:116:8  */
  assign dma_update_en = n1068_o; // (signal)
  /* ni/packet_manager.vhd:117:8  */
  assign dma_update_addr = dma_num_reg; // (signal)
  /* ni/packet_manager.vhd:118:8  */
  assign dma_update_data = n1206_o; // (signal)
  /* ni/packet_manager.vhd:131:8  */
  assign port_a_wr_hi = n1118_o; // (signal)
  /* ni/packet_manager.vhd:132:8  */
  assign port_a_wr_lo = n1121_o; // (signal)
  /* ni/packet_manager.vhd:133:8  */
  assign port_a_addr = n1103_o; // (signal)
  /* ni/packet_manager.vhd:134:8  */
  assign port_a_din = n1207_o; // (signal)
  /* ni/packet_manager.vhd:135:8  */
  assign port_a_dout = n1208_o; // (signal)
  /* ni/packet_manager.vhd:137:8  */
  assign config_slv_error_next = n1158_o; // (signal)
  /* ni/packet_manager.vhd:139:8  */
  assign pkt_len_reg = n1202_q; // (signal)
  /* ni/packet_manager.vhd:139:21  */
  assign pkt_len_next = n1080_o; // (signal)
  /* ni/packet_manager.vhd:141:8  */
  assign route_reg = n1203_q; // (signal)
  /* ni/packet_manager.vhd:147:8  */
  assign payload_data = n1204_q; // (signal)
  /* ni/packet_manager.vhd:147:22  */
  assign payload_data_next = n1209_o; // (signal)
  assign n872_o = dmatbl_data[29:16];
  /* ni/packet_manager.vhd:167:3  */
  assign n873_o = dma_en ? pkt_len : pkt_len_reg;
  assign n874_o = dmatbl_data[15:14];
  /* ni/packet_manager.vhd:179:26  */
  assign n876_o = $unsigned(pkt_len_reg) >= $unsigned(4'b0001);
  /* ni/packet_manager.vhd:179:11  */
  assign n878_o = n876_o ? 2'b01 : n874_o;
  /* ni/packet_manager.vhd:182:49  */
  assign n880_o = {3'b110, pkt_type};
  /* ni/packet_manager.vhd:182:60  */
  assign n882_o = {n880_o, 3'b011};
  /* ni/packet_manager.vhd:182:70  */
  assign n884_o = {n882_o, 11'b00000000000};
  /* ni/packet_manager.vhd:182:103  */
  assign n885_o = {n884_o, route_reg};
  assign n886_o = dmatbl_data[44];
  assign n888_o = dmatbl_data[29:16];
  assign n889_o = dmatbl_data[29:16];
  assign n890_o = dmatbl_data[43:30];
  /* ni/packet_manager.vhd:191:30  */
  assign n892_o = n890_o - 14'b00000000000001;
  assign n893_o = dmatbl_data[43:30];
  /* ni/packet_manager.vhd:192:20  */
  assign n894_o = {10'b0, pkt_len_reg};  //  uext
  /* ni/packet_manager.vhd:192:20  */
  assign n895_o = $unsigned(n893_o) > $unsigned(n894_o);
  assign n896_o = dmatbl_data[15:14];
  /* ni/packet_manager.vhd:193:29  */
  assign n898_o = n896_o == 2'b10;
  /* ni/packet_manager.vhd:185:9  */
  assign n900_o = n935_o ? 2'b00 : n874_o;
  /* ni/packet_manager.vhd:192:11  */
  assign n902_o = n895_o & n898_o;
  /* ni/packet_manager.vhd:192:11  */
  assign n903_o = n895_o ? 1'b1 : 1'b0;
  /* ni/packet_manager.vhd:199:43  */
  assign n904_o = dmatbl_data[13:0];
  /* ni/packet_manager.vhd:199:68  */
  assign n905_o = {10'b0, pkt_len_reg};  //  uext
  /* ni/packet_manager.vhd:199:68  */
  assign n906_o = n904_o + n905_o;
  assign n907_o = dmatbl_data[29:16];
  /* ni/packet_manager.vhd:200:39  */
  assign n908_o = {10'b0, pkt_len_reg};  //  uext
  /* ni/packet_manager.vhd:200:39  */
  assign n909_o = n907_o + n908_o;
  assign n910_o = dmatbl_data[43:30];
  /* ni/packet_manager.vhd:201:33  */
  assign n911_o = {10'b0, pkt_len_reg};  //  uext
  /* ni/packet_manager.vhd:201:33  */
  assign n912_o = n910_o - n911_o;
  assign n913_o = dmatbl_data[15:14];
  /* ni/packet_manager.vhd:202:27  */
  assign n915_o = n913_o == 2'b01;
  /* ni/packet_manager.vhd:205:43  */
  assign n916_o = dmatbl_data[13:10];
  assign n917_o = n906_o[13:10];
  /* ni/packet_manager.vhd:202:11  */
  assign n918_o = n915_o ? n916_o : n917_o;
  assign n919_o = n906_o[9:0];
  /* ni/packet_manager.vhd:207:39  */
  assign n921_o = pkt_len_reg - 4'b0001;
  /* ni/packet_manager.vhd:208:49  */
  assign n923_o = {3'b110, pkt_type};
  /* ni/packet_manager.vhd:208:68  */
  assign n924_o = dmatbl_data[13:0];
  /* ni/packet_manager.vhd:208:60  */
  assign n925_o = {n923_o, n924_o};
  /* ni/packet_manager.vhd:208:93  */
  assign n926_o = {n925_o, route_reg};
  assign n927_o = {2'b11, n888_o};
  assign n928_o = {2'b00, n872_o};
  /* ni/packet_manager.vhd:185:9  */
  assign n929_o = n886_o ? n927_o : n928_o;
  /* ni/packet_manager.vhd:185:9  */
  assign n931_o = n886_o ? n926_o : 35'b00000000000000000000000000000000000;
  /* ni/packet_manager.vhd:185:9  */
  assign n933_o = n886_o ? 3'b001 : state;
  /* ni/packet_manager.vhd:185:9  */
  assign n934_o = n886_o ? n892_o : count_reg;
  /* ni/packet_manager.vhd:185:9  */
  assign n935_o = n886_o & n902_o;
  /* ni/packet_manager.vhd:185:9  */
  assign n936_o = n886_o ? n889_o : read_ptr_reg;
  /* ni/packet_manager.vhd:185:9  */
  assign n939_o = n886_o ? 1'b1 : 1'b0;
  assign n940_o = {n918_o, n919_o};
  assign n941_o = {n903_o, n912_o, n909_o};
  assign n942_o = dmatbl_data[13:0];
  /* ni/packet_manager.vhd:185:9  */
  assign n943_o = n886_o ? n940_o : n942_o;
  assign n944_o = dmatbl_data[43:16];
  assign n945_o = {1'b0, n944_o};
  /* ni/packet_manager.vhd:185:9  */
  assign n946_o = n886_o ? n941_o : n945_o;
  /* ni/packet_manager.vhd:185:9  */
  assign n947_o = n886_o ? n921_o : n873_o;
  assign n948_o = {2'b00, n872_o};
  /* ni/packet_manager.vhd:177:9  */
  assign n949_o = mc ? n948_o : n929_o;
  /* ni/packet_manager.vhd:177:9  */
  assign n950_o = mc ? n885_o : n931_o;
  /* ni/packet_manager.vhd:177:9  */
  assign n952_o = mc ? 3'b011 : n933_o;
  /* ni/packet_manager.vhd:177:9  */
  assign n953_o = mc ? count_reg : n934_o;
  /* ni/packet_manager.vhd:177:9  */
  assign n954_o = mc ? n878_o : n900_o;
  /* ni/packet_manager.vhd:177:9  */
  assign n955_o = mc ? read_ptr_reg : n936_o;
  /* ni/packet_manager.vhd:177:9  */
  assign n957_o = mc ? 1'b0 : n939_o;
  assign n958_o = dmatbl_data[13:0];
  /* ni/packet_manager.vhd:177:9  */
  assign n959_o = mc ? n958_o : n943_o;
  assign n960_o = dmatbl_data[43:16];
  assign n961_o = {1'b0, n960_o};
  /* ni/packet_manager.vhd:177:9  */
  assign n962_o = mc ? n961_o : n946_o;
  /* ni/packet_manager.vhd:177:9  */
  assign n963_o = mc ? n873_o : n947_o;
  /* ni/packet_manager.vhd:177:9  */
  assign n965_o = mc ? mc_idx : 2'b00;
  /* ni/packet_manager.vhd:177:9  */
  assign n967_o = mc ? mc_p : 2'b00;
  assign n968_o = {2'b00, n872_o};
  /* ni/packet_manager.vhd:176:7  */
  assign n969_o = dma_en_reg ? n949_o : n968_o;
  /* ni/packet_manager.vhd:176:7  */
  assign n971_o = dma_en_reg ? n950_o : 35'b00000000000000000000000000000000000;
  /* ni/packet_manager.vhd:176:7  */
  assign n972_o = dma_en_reg ? n952_o : state;
  /* ni/packet_manager.vhd:176:7  */
  assign n973_o = dma_en_reg ? n953_o : count_reg;
  /* ni/packet_manager.vhd:176:7  */
  assign n974_o = dma_en_reg ? n954_o : n874_o;
  /* ni/packet_manager.vhd:176:7  */
  assign n975_o = dma_en_reg ? n955_o : read_ptr_reg;
  /* ni/packet_manager.vhd:176:7  */
  assign n977_o = dma_en_reg ? n957_o : 1'b0;
  assign n978_o = dmatbl_data[13:0];
  /* ni/packet_manager.vhd:176:7  */
  assign n979_o = dma_en_reg ? n959_o : n978_o;
  assign n980_o = dmatbl_data[43:16];
  assign n981_o = {1'b0, n980_o};
  /* ni/packet_manager.vhd:176:7  */
  assign n982_o = dma_en_reg ? n962_o : n981_o;
  /* ni/packet_manager.vhd:176:7  */
  assign n983_o = dma_en_reg ? n963_o : n873_o;
  /* ni/packet_manager.vhd:176:7  */
  assign n985_o = dma_en_reg ? n965_o : 2'b00;
  /* ni/packet_manager.vhd:176:7  */
  assign n987_o = dma_en_reg ? n967_o : 2'b00;
  /* ni/packet_manager.vhd:175:5  */
  assign n989_o = state == 3'b000;
  /* ni/packet_manager.vhd:213:41  */
  assign n990_o = n864_o[31:0];
  /* ni/packet_manager.vhd:214:35  */
  assign n992_o = pkt_len_reg - 4'b0001;
  /* ni/packet_manager.vhd:215:31  */
  assign n994_o = count_reg - 14'b00000000000001;
  /* ni/packet_manager.vhd:216:22  */
  assign n996_o = $unsigned(pkt_len_reg) > $unsigned(4'b0000);
  /* ni/packet_manager.vhd:216:40  */
  assign n998_o = $unsigned(count_reg) > $unsigned(14'b00000000000000);
  /* ni/packet_manager.vhd:216:26  */
  assign n999_o = n996_o & n998_o;
  /* ni/packet_manager.vhd:218:58  */
  assign n1000_o = n864_o[63:32];
  /* ni/packet_manager.vhd:218:43  */
  assign n1002_o = {3'b100, n1000_o};
  /* ni/packet_manager.vhd:219:39  */
  assign n1004_o = read_ptr_reg + 14'b00000000000001;
  /* ni/packet_manager.vhd:222:62  */
  assign n1005_o = n864_o[63:32];
  /* ni/packet_manager.vhd:222:47  */
  assign n1007_o = {3'b101, n1005_o};
  /* ni/packet_manager.vhd:216:7  */
  assign n1008_o = n999_o ? n1002_o : n1007_o;
  /* ni/packet_manager.vhd:216:7  */
  assign n1011_o = n999_o ? 3'b010 : 3'b000;
  /* ni/packet_manager.vhd:216:7  */
  assign n1012_o = n999_o ? n1004_o : read_ptr_reg;
  /* ni/packet_manager.vhd:212:5  */
  assign n1014_o = state == 3'b001;
  /* ni/packet_manager.vhd:226:35  */
  assign n1016_o = pkt_len_reg - 4'b0001;
  /* ni/packet_manager.vhd:227:31  */
  assign n1018_o = count_reg - 14'b00000000000001;
  /* ni/packet_manager.vhd:228:22  */
  assign n1020_o = $unsigned(pkt_len_reg) > $unsigned(4'b0000);
  /* ni/packet_manager.vhd:228:40  */
  assign n1022_o = $unsigned(count_reg) > $unsigned(14'b00000000000000);
  /* ni/packet_manager.vhd:228:26  */
  assign n1023_o = n1020_o & n1022_o;
  /* ni/packet_manager.vhd:230:43  */
  assign n1025_o = {3'b100, payload_data};
  /* ni/packet_manager.vhd:232:39  */
  assign n1028_o = read_ptr_reg + 14'b00000000000001;
  /* ni/packet_manager.vhd:238:47  */
  assign n1030_o = {3'b101, payload_data};
  assign n1031_o = {2'b11, read_ptr_next};
  assign n1032_o = {2'b00, n872_o};
  /* ni/packet_manager.vhd:228:7  */
  assign n1033_o = n1023_o ? n1031_o : n1032_o;
  /* ni/packet_manager.vhd:228:7  */
  assign n1034_o = n1023_o ? n1025_o : n1030_o;
  /* ni/packet_manager.vhd:228:7  */
  assign n1037_o = n1023_o ? 3'b001 : 3'b000;
  /* ni/packet_manager.vhd:228:7  */
  assign n1038_o = n1023_o ? n1028_o : read_ptr_reg;
  /* ni/packet_manager.vhd:225:5  */
  assign n1040_o = state == 3'b010;
  /* ni/packet_manager.vhd:243:41  */
  assign n1042_o = {3'b100, payload_data};
  /* ni/packet_manager.vhd:241:5  */
  assign n1044_o = state == 3'b011;
  /* ni/packet_manager.vhd:247:45  */
  assign n1046_o = {3'b101, payload_data};
  /* ni/packet_manager.vhd:245:5  */
  assign n1048_o = state == 3'b100;
  assign n1049_o = {n1048_o, n1044_o, n1040_o, n1014_o, n989_o};
  assign n1050_o = {2'b00, n872_o};
  /* ni/packet_manager.vhd:174:3  */
  always @*
    case (n1049_o)
      5'b10000: n1052_o <= n1050_o;
      5'b01000: n1052_o <= n1050_o;
      5'b00100: n1052_o <= n1033_o;
      5'b00010: n1052_o <= n1050_o;
      5'b00001: n1052_o <= n969_o;
      default: n1052_o <= 16'bX;
    endcase
  /* ni/packet_manager.vhd:174:3  */
  always @*
    case (n1049_o)
      5'b10000: n1054_o <= n1046_o;
      5'b01000: n1054_o <= n1042_o;
      5'b00100: n1054_o <= n1034_o;
      5'b00010: n1054_o <= n1008_o;
      5'b00001: n1054_o <= n971_o;
      default: n1054_o <= 35'bX;
    endcase
  /* ni/packet_manager.vhd:174:3  */
  always @*
    case (n1049_o)
      5'b10000: n1059_o <= 3'b000;
      5'b01000: n1059_o <= 3'b100;
      5'b00100: n1059_o <= n1037_o;
      5'b00010: n1059_o <= n1011_o;
      5'b00001: n1059_o <= n972_o;
      default: n1059_o <= 3'bX;
    endcase
  /* ni/packet_manager.vhd:174:3  */
  always @*
    case (n1049_o)
      5'b10000: n1061_o <= count_reg;
      5'b01000: n1061_o <= count_reg;
      5'b00100: n1061_o <= n1018_o;
      5'b00010: n1061_o <= n994_o;
      5'b00001: n1061_o <= n973_o;
      default: n1061_o <= 14'bX;
    endcase
  /* ni/packet_manager.vhd:174:3  */
  always @*
    case (n1049_o)
      5'b10000: n1063_o <= n874_o;
      5'b01000: n1063_o <= n874_o;
      5'b00100: n1063_o <= n874_o;
      5'b00010: n1063_o <= n874_o;
      5'b00001: n1063_o <= n974_o;
      default: n1063_o <= 2'bX;
    endcase
  /* ni/packet_manager.vhd:174:3  */
  always @*
    case (n1049_o)
      5'b10000: n1065_o <= read_ptr_reg;
      5'b01000: n1065_o <= read_ptr_reg;
      5'b00100: n1065_o <= n1038_o;
      5'b00010: n1065_o <= n1012_o;
      5'b00001: n1065_o <= n975_o;
      default: n1065_o <= 14'bX;
    endcase
  /* ni/packet_manager.vhd:174:3  */
  always @*
    case (n1049_o)
      5'b10000: n1068_o <= 1'b0;
      5'b01000: n1068_o <= 1'b0;
      5'b00100: n1068_o <= 1'b0;
      5'b00010: n1068_o <= 1'b0;
      5'b00001: n1068_o <= n977_o;
      default: n1068_o <= 1'bX;
    endcase
  assign n1070_o = dmatbl_data[13:0];
  /* ni/packet_manager.vhd:174:3  */
  always @*
    case (n1049_o)
      5'b10000: n1072_o <= n1070_o;
      5'b01000: n1072_o <= n1070_o;
      5'b00100: n1072_o <= n1070_o;
      5'b00010: n1072_o <= n1070_o;
      5'b00001: n1072_o <= n979_o;
      default: n1072_o <= 14'bX;
    endcase
  assign n1073_o = dmatbl_data[43:16];
  assign n1074_o = {1'b0, n1073_o};
  /* ni/packet_manager.vhd:174:3  */
  always @*
    case (n1049_o)
      5'b10000: n1076_o <= n1074_o;
      5'b01000: n1076_o <= n1074_o;
      5'b00100: n1076_o <= n1074_o;
      5'b00010: n1076_o <= n1074_o;
      5'b00001: n1076_o <= n982_o;
      default: n1076_o <= 29'bX;
    endcase
  assign n1078_o = dmatbl_data[15:14];
  /* ni/packet_manager.vhd:174:3  */
  always @*
    case (n1049_o)
      5'b10000: n1080_o <= n873_o;
      5'b01000: n1080_o <= n873_o;
      5'b00100: n1080_o <= n1016_o;
      5'b00010: n1080_o <= n992_o;
      5'b00001: n1080_o <= n983_o;
      default: n1080_o <= 4'bX;
    endcase
  assign n1081_o = n990_o[1:0];
  /* ni/packet_manager.vhd:174:3  */
  always @*
    case (n1049_o)
      5'b10000: n1084_o <= 2'b00;
      5'b01000: n1084_o <= 2'b00;
      5'b00100: n1084_o <= 2'b00;
      5'b00010: n1084_o <= n1081_o;
      5'b00001: n1084_o <= n985_o;
      default: n1084_o <= 2'bX;
    endcase
  assign n1085_o = n990_o[15:2];
  /* ni/packet_manager.vhd:174:3  */
  always @*
    case (n1049_o)
      5'b10000: n1088_o <= 14'b00000000000000;
      5'b01000: n1088_o <= 14'b00000000000000;
      5'b00100: n1088_o <= 14'b00000000000000;
      5'b00010: n1088_o <= n1085_o;
      5'b00001: n1088_o <= 14'b00000000000000;
      default: n1088_o <= 14'bX;
    endcase
  assign n1089_o = n990_o[17:16];
  /* ni/packet_manager.vhd:174:3  */
  always @*
    case (n1049_o)
      5'b10000: n1092_o <= 2'b00;
      5'b01000: n1092_o <= 2'b00;
      5'b00100: n1092_o <= 2'b00;
      5'b00010: n1092_o <= n1089_o;
      5'b00001: n1092_o <= n987_o;
      default: n1092_o <= 2'bX;
    endcase
  assign n1093_o = n990_o[31:18];
  /* ni/packet_manager.vhd:174:3  */
  always @*
    case (n1049_o)
      5'b10000: n1096_o <= 14'b00000000000000;
      5'b01000: n1096_o <= 14'b00000000000000;
      5'b00100: n1096_o <= 14'b00000000000000;
      5'b00010: n1096_o <= n1093_o;
      5'b00001: n1096_o <= 14'b00000000000000;
      default: n1096_o <= 14'bX;
    endcase
  /* ni/packet_manager.vhd:256:29  */
  assign n1103_o = n855_o[6:1];
  /* ni/packet_manager.vhd:259:52  */
  assign n1105_o = n855_o[47];
  /* ni/packet_manager.vhd:262:26  */
  assign n1106_o = n855_o[43:16];
  /* ni/packet_manager.vhd:264:48  */
  assign n1107_o = n855_o[31:16];
  /* ni/packet_manager.vhd:266:17  */
  assign n1108_o = n855_o[0];
  /* ni/packet_manager.vhd:272:28  */
  assign n1109_o = n855_o[15];
  /* ni/packet_manager.vhd:272:31  */
  assign n1110_o = n1109_o & sel;
  /* ni/packet_manager.vhd:273:20  */
  assign n1111_o = n855_o[0];
  /* ni/packet_manager.vhd:273:24  */
  assign n1112_o = ~n1111_o;
  /* ni/packet_manager.vhd:277:28  */
  assign n1113_o = n855_o[15];
  /* ni/packet_manager.vhd:277:31  */
  assign n1114_o = n1113_o & sel;
  /* ni/packet_manager.vhd:273:3  */
  assign n1116_o = n1112_o ? n1114_o : 1'b0;
  /* ni/packet_manager.vhd:266:3  */
  assign n1118_o = n1108_o ? n1110_o : 1'b0;
  /* ni/packet_manager.vhd:266:3  */
  assign n1121_o = n1108_o ? 1'b0 : n1116_o;
  /* ni/packet_manager.vhd:280:28  */
  assign n1123_o = n855_o[0];
  /* ni/packet_manager.vhd:282:50  */
  assign n1124_o = port_a_dout[44];
  /* ni/packet_manager.vhd:284:32  */
  assign n1125_o = port_a_dout[43:16];
  /* ni/packet_manager.vhd:287:48  */
  assign n1126_o = port_a_dout[15:0];
  assign n1127_o = n1125_o[15:0];
  /* ni/packet_manager.vhd:281:3  */
  assign n1128_o = hi_lo_reg ? n1127_o : n1126_o;
  assign n1129_o = n1125_o[27:16];
  assign n1130_o = n1104_o[27:16];
  /* ni/packet_manager.vhd:281:3  */
  assign n1131_o = hi_lo_reg ? n1129_o : n1130_o;
  assign n1132_o = n1104_o[31];
  /* ni/packet_manager.vhd:281:3  */
  assign n1133_o = hi_lo_reg ? n1124_o : n1132_o;
  assign n1136_o = n1104_o[30:28];
  /* ni/packet_manager.vhd:297:3  */
  assign n1140_o = dma_en ? 1'b0 : dma_update_en;
  /* ni/packet_manager.vhd:297:3  */
  assign n1141_o = dma_en ? dma_num : dma_update_addr;
  /* ni/packet_manager.vhd:308:1  */
  tdp_ram_29_6 dmatbl1 (
    .a_clk(clk),
    .a_wr(port_a_wr_hi),
    .a_addr(port_a_addr),
    .a_din(n1143_o),
    .b_clk(clk),
    .b_wr(port_b_wr),
    .b_addr(port_b_addr),
    .b_din(n1145_o),
    .a_dout(dmatbl1_a_dout),
    .b_dout(dmatbl1_b_dout));
  /* ni/packet_manager.vhd:317:26  */
  assign n1143_o = port_a_din[44:16];
  /* ni/packet_manager.vhd:322:26  */
  assign n1145_o = port_b_din[44:16];
  /* ni/packet_manager.vhd:327:3  */
  tdp_ram_16_6 dmatbl2 (
    .a_clk(clk),
    .a_wr(port_a_wr_lo),
    .a_addr(port_a_addr),
    .a_din(n1147_o),
    .b_clk(clk),
    .b_wr(port_b_wr),
    .b_addr(port_b_addr),
    .b_din(n1149_o),
    .a_dout(dmatbl2_a_dout),
    .b_dout(dmatbl2_b_dout));
  /* ni/packet_manager.vhd:336:26  */
  assign n1147_o = port_a_din[15:0];
  /* ni/packet_manager.vhd:341:26  */
  assign n1149_o = port_b_din[15:0];
  /* ni/packet_manager.vhd:348:31  */
  assign n1152_o = n855_o[10:7];
  /* ni/packet_manager.vhd:348:77  */
  assign n1154_o = n1152_o != 4'b0000;
  /* ni/packet_manager.vhd:348:16  */
  assign n1155_o = sel & n1154_o;
  /* ni/packet_manager.vhd:348:3  */
  assign n1158_o = n1155_o ? 1'b1 : 1'b0;
  /* ni/packet_manager.vhd:357:5  */
  assign n1164_o = reset ? 1'b0 : dma_en;
  /* ni/packet_manager.vhd:356:3  */
  always @(posedge clk)
    n1167_q <= n1164_o;
  /* ni/packet_manager.vhd:368:5  */
  assign n1171_o = reset ? 1'b0 : hi_lo_next;
  /* ni/packet_manager.vhd:367:3  */
  always @(posedge clk)
    n1174_q <= n1171_o;
  /* ni/packet_manager.vhd:379:5  */
  assign n1178_o = reset ? 1'b0 : config_slv_error_next;
  /* ni/packet_manager.vhd:378:3  */
  always @(posedge clk)
    n1182_q <= n1178_o;
  /* ni/packet_manager.vhd:390:5  */
  assign n1186_o = reset ? 3'b000 : next_state;
  /* ni/packet_manager.vhd:389:3  */
  always @(posedge clk)
    n1189_q <= n1186_o;
  /* ni/packet_manager.vhd:401:3  */
  always @(posedge clk)
    n1199_q <= count_next;
  /* ni/packet_manager.vhd:401:3  */
  always @(posedge clk)
    n1200_q <= read_ptr_next;
  /* ni/packet_manager.vhd:401:3  */
  always @(posedge clk)
    n1201_q <= dma_num;
  /* ni/packet_manager.vhd:401:3  */
  always @(posedge clk)
    n1202_q <= pkt_len_next;
  /* ni/packet_manager.vhd:401:3  */
  always @(posedge clk)
    n1203_q <= route;
  /* ni/packet_manager.vhd:401:3  */
  always @(posedge clk)
    n1204_q <= payload_data_next;
  /* ni/packet_manager.vhd:401:3  */
  assign n1205_o = {dmatbl1_b_dout, dmatbl2_b_dout};
  assign n1206_o = {n1076_o, n1078_o, n1072_o};
  assign n1207_o = {n1105_o, n1106_o, n1107_o};
  assign n1208_o = {dmatbl1_a_dout, dmatbl2_a_dout};
  assign n1209_o = {n1096_o, n1092_o, n1088_o, n1084_o};
  assign n1210_o = {n1182_q, n1133_o, n1136_o, n1131_o, n1128_o};
  assign n1211_o = {64'b0000000000000000000000000000000000000000000000000000000000000000, 1'b0, n1052_o};
endmodule

module schedule_table
  (input  clk,
   input  reset,
   input  [13:0] config_addr,
   input  config_en,
   input  config_wr,
   input  [31:0] config_wdata,
   input  sel,
   input  [7:0] stbl_idx,
   input  stbl_idx_en,
   output [31:0] config_slv_rdata,
   output config_slv_error,
   output [15:0] route,
   output [3:0] pkt_len,
   output [3:0] t2n,
   output [5:0] dma_num,
   output dma_en);
  wire [47:0] n783_o;
  wire [31:0] n785_o;
  wire n786_o;
  wire [29:0] stbl_data;
  wire stbl_idx_en_reg;
  wire config_slv_error_next;
  wire [5:0] dma_num_sig;
  wire [29:0] port_a_din;
  wire [29:0] port_a_dout;
  wire a_wr;
  wire n792_o;
  wire n793_o;
  wire [29:0] stbl_a_dout;
  wire [29:0] stbl_b_dout;
  wire [7:0] n794_o;
  localparam n796_o = 1'b0;
  localparam [29:0] n797_o = 30'b000000000000000000000000000000;
  localparam [31:0] n800_o = 32'b00000000000000000000000000000000;
  wire [15:0] n801_o;
  wire [5:0] n803_o;
  wire [1:0] n804_o;
  wire [3:0] n806_o;
  wire [3:0] n808_o;
  wire [15:0] n809_o;
  wire [5:0] n812_o;
  wire [3:0] n814_o;
  wire [3:0] n816_o;
  wire [2:0] n819_o;
  wire n821_o;
  wire n822_o;
  wire n825_o;
  wire [15:0] n828_o;
  wire [5:0] n829_o;
  wire [3:0] n830_o;
  wire [3:0] n831_o;
  wire n835_o;
  reg n838_q;
  wire n841_o;
  wire n843_o;
  wire n848_o;
  reg n852_q;
  wire [29:0] n853_o;
  wire [32:0] n854_o;
  assign config_slv_rdata = n785_o;
  assign config_slv_error = n786_o;
  assign route = n828_o;
  assign pkt_len = n830_o;
  assign t2n = n831_o;
  assign dma_num = dma_num_sig;
  assign dma_en = n843_o;
  /* ni/MC_controller.vhd:258:32  */
  assign n783_o = {config_wdata, config_wr, config_en, config_addr};
  /* ni/MC_controller.vhd:101:40  */
  assign n785_o = n854_o[31:0];
  /* ni/MC_controller.vhd:101:24  */
  assign n786_o = n854_o[32];
  /* ni/schedule_table.vhd:78:8  */
  assign stbl_data = stbl_b_dout; // (signal)
  /* ni/schedule_table.vhd:80:8  */
  assign stbl_idx_en_reg = n838_q; // (signal)
  /* ni/schedule_table.vhd:82:8  */
  assign config_slv_error_next = n825_o; // (signal)
  /* ni/schedule_table.vhd:84:8  */
  assign dma_num_sig = n829_o; // (signal)
  /* ni/schedule_table.vhd:86:8  */
  assign port_a_din = n853_o; // (signal)
  /* ni/schedule_table.vhd:86:20  */
  assign port_a_dout = stbl_a_dout; // (signal)
  /* ni/schedule_table.vhd:88:8  */
  assign a_wr = n793_o; // (signal)
  /* ni/schedule_table.vhd:91:18  */
  assign n792_o = n783_o[15];
  /* ni/schedule_table.vhd:91:21  */
  assign n793_o = n792_o & sel;
  /* ni/schedule_table.vhd:93:1  */
  tdp_ram_30_8 stbl (
    .a_clk(clk),
    .a_wr(a_wr),
    .a_addr(n794_o),
    .a_din(port_a_din),
    .b_clk(clk),
    .b_wr(n796_o),
    .b_addr(stbl_idx),
    .b_din(n797_o),
    .a_dout(stbl_a_dout),
    .b_dout(stbl_b_dout));
  /* ni/schedule_table.vhd:101:27  */
  assign n794_o = n783_o[7:0];
  /* ni/schedule_table.vhd:117:33  */
  assign n801_o = port_a_dout[29:14];
  /* ni/schedule_table.vhd:121:33  */
  assign n803_o = port_a_dout[13:8];
  assign n804_o = n800_o[15:14];
  /* ni/schedule_table.vhd:125:33  */
  assign n806_o = port_a_dout[7:4];
  /* ni/schedule_table.vhd:129:33  */
  assign n808_o = port_a_dout[3:0];
  /* ni/schedule_table.vhd:135:34  */
  assign n809_o = n783_o[47:32];
  /* ni/schedule_table.vhd:140:34  */
  assign n812_o = n783_o[29:24];
  /* ni/schedule_table.vhd:143:34  */
  assign n814_o = n783_o[23:20];
  /* ni/schedule_table.vhd:146:34  */
  assign n816_o = n783_o[19:16];
  /* ni/schedule_table.vhd:154:31  */
  assign n819_o = n783_o[10:8];
  /* ni/schedule_table.vhd:154:73  */
  assign n821_o = n819_o != 3'b000;
  /* ni/schedule_table.vhd:154:16  */
  assign n822_o = sel & n821_o;
  /* ni/schedule_table.vhd:154:3  */
  assign n825_o = n822_o ? 1'b1 : 1'b0;
  /* ni/schedule_table.vhd:159:21  */
  assign n828_o = stbl_data[29:14];
  /* ni/schedule_table.vhd:161:34  */
  assign n829_o = stbl_data[13:8];
  /* ni/schedule_table.vhd:164:30  */
  assign n830_o = stbl_data[7:4];
  /* ni/schedule_table.vhd:166:30  */
  assign n831_o = stbl_data[3:0];
  /* ni/schedule_table.vhd:172:5  */
  assign n835_o = reset ? 1'b0 : stbl_idx_en;
  /* ni/schedule_table.vhd:171:3  */
  always @(posedge clk)
    n838_q <= n835_o;
  /* ni/schedule_table.vhd:183:18  */
  assign n841_o = dma_num_sig == 6'b111111;
  /* ni/schedule_table.vhd:183:3  */
  assign n843_o = n841_o ? 1'b0 : stbl_idx_en_reg;
  /* ni/schedule_table.vhd:193:5  */
  assign n848_o = reset ? 1'b0 : config_slv_error_next;
  /* ni/schedule_table.vhd:192:3  */
  always @(posedge clk)
    n852_q <= n848_o;
  /* ni/schedule_table.vhd:192:3  */
  assign n853_o = {n809_o, n812_o, n814_o, n816_o};
  assign n854_o = {n852_q, n801_o, n804_o, n803_o, n806_o, n808_o};
endmodule

module mc_controller_5ba93c9db0cff93f52b521d7420e43f6eda2784f
  (input  clk,
   input  reset,
   input  run,
   input  [13:0] config_addr,
   input  config_en,
   input  config_wr,
   input  [31:0] config_wdata,
   input  sel,
   input  period_boundary,
   input  [1:0] mc_p_cnt,
   output [31:0] config_slv_rdata,
   output config_slv_error,
   output [7:0] stbl_min,
   output [7:0] stbl_maxp1,
   output mc,
   output [1:0] mc_idx,
   output [1:0] mc_p);
  wire [47:0] n544_o;
  wire [31:0] n546_o;
  wire n547_o;
  wire [7:0] stbl_min_next;
  wire [7:0] stbl_maxp1_next;
  wire [1:0] mode_change_idx_reg;
  wire [1:0] mode_change_idx_next;
  wire [1:0] mode_idx_reg;
  wire [1:0] mode_change_cnt_reg;
  wire [1:0] mode_change_cnt_next;
  wire [1:0] mode_change_cnt_int;
  wire [63:0] mode_reg;
  wire [63:0] mode_next;
  wire global_mode_change_idx;
  wire local_mode_change_idx;
  wire config_slv_error_next;
  wire [31:0] read_reg;
  wire [31:0] read_next;
  wire mode_changed_reg;
  wire [7:0] stbl_min_reg;
  wire [10:0] mc_tbl_addr;
  wire [10:0] n556_o;
  wire [10:0] n558_o;
  wire n559_o;
  wire n560_o;
  wire n561_o;
  wire n562_o;
  wire [10:0] n563_o;
  wire n565_o;
  reg n568_o;
  wire [1:0] n569_o;
  reg [1:0] n570_o;
  wire [10:0] n571_o;
  wire [1:0] n572_o;
  wire n574_o;
  wire n576_o;
  wire [1:0] n577_o;
  reg [1:0] n578_o;
  reg [1:0] n579_o;
  reg n582_o;
  reg n585_o;
  wire n587_o;
  wire [1:0] n589_o;
  wire [7:0] n591_o;
  wire [1:0] n594_o;
  wire [7:0] n596_o;
  wire [63:0] n598_o;
  wire n600_o;
  wire [1:0] n601_o;
  wire [1:0] n602_o;
  wire [63:0] n603_o;
  wire n605_o;
  wire n606_o;
  wire [1:0] n607_o;
  wire [1:0] n608_o;
  wire [1:0] n609_o;
  wire [1:0] n610_o;
  wire [63:0] n611_o;
  wire n613_o;
  wire n616_o;
  wire n619_o;
  wire [29:0] n620_o;
  localparam n622_o = 1'b0;
  localparam [1:0] n623_o = 2'b00;
  wire [1:0] n624_o;
  localparam [1:0] n625_o = 2'b00;
  wire n629_o;
  wire n631_o;
  wire n633_o;
  reg n636_q;
  wire n638_o;
  wire n641_o;
  wire n643_o;
  wire [7:0] n649_o;
  wire [7:0] n653_o;
  wire [7:0] n655_o;
  wire n660_o;
  wire [1:0] n664_o;
  wire [31:0] n666_o;
  reg n676_q;
  reg [1:0] n678_q;
  reg [31:0] n679_q;
  wire [63:0] n684_o;
  reg [63:0] n687_q;
  wire [1:0] n690_o;
  wire [1:0] n692_o;
  reg [1:0] n695_q;
  wire [1:0] n698_o;
  wire [1:0] n700_o;
  reg [1:0] n703_q;
  wire [7:0] n706_o;
  wire [7:0] n709_o;
  reg [7:0] n715_q;
  wire [7:0] n719_o;
  wire [7:0] n721_o;
  reg [7:0] n724_q;
  wire [31:0] n726_o;
  wire [32:0] n728_o;
  wire n729_o;
  wire n730_o;
  wire n731_o;
  wire n732_o;
  wire n733_o;
  wire n734_o;
  wire n735_o;
  wire n736_o;
  wire [7:0] n737_o;
  wire [7:0] n738_o;
  wire [7:0] n739_o;
  wire [7:0] n740_o;
  wire [7:0] n741_o;
  wire [7:0] n742_o;
  wire [7:0] n743_o;
  wire [7:0] n744_o;
  wire [7:0] n745_o;
  wire [7:0] n746_o;
  wire [7:0] n747_o;
  wire [7:0] n748_o;
  wire [63:0] n749_o;
  wire n750_o;
  wire n751_o;
  wire n752_o;
  wire n753_o;
  wire n754_o;
  wire n755_o;
  wire n756_o;
  wire n757_o;
  wire [7:0] n758_o;
  wire [7:0] n759_o;
  wire [7:0] n760_o;
  wire [7:0] n761_o;
  wire [7:0] n762_o;
  wire [7:0] n763_o;
  wire [7:0] n764_o;
  wire [7:0] n765_o;
  wire [7:0] n766_o;
  wire [7:0] n767_o;
  wire [7:0] n768_o;
  wire [7:0] n769_o;
  wire [63:0] n770_o;
  wire [15:0] n771_o;
  wire [15:0] n772_o;
  wire [15:0] n773_o;
  wire [15:0] n774_o;
  wire [1:0] n775_o;
  reg [15:0] n776_o;
  wire [15:0] n777_o;
  wire [15:0] n778_o;
  wire [15:0] n779_o;
  wire [15:0] n780_o;
  wire [1:0] n781_o;
  reg [15:0] n782_o;
  assign config_slv_rdata = n546_o;
  assign config_slv_error = n547_o;
  assign stbl_min = n655_o;
  assign stbl_maxp1 = n724_q;
  assign mc = n622_o;
  assign mc_idx = n623_o;
  assign mc_p = n625_o;
  /* ni/TDM_controller.vhd:64:5  */
  assign n544_o = {config_wdata, config_wr, config_en, config_addr};
  /* ni/TDM_controller.vhd:60:5  */
  assign n546_o = n728_o[31:0];
  /* ni/TDM_controller.vhd:58:5  */
  assign n547_o = n728_o[32];
  /* ni/MC_controller.vhd:86:10  */
  assign stbl_min_next = n649_o; // (signal)
  /* ni/MC_controller.vhd:86:25  */
  assign stbl_maxp1_next = n653_o; // (signal)
  /* ni/MC_controller.vhd:87:10  */
  assign mode_change_idx_reg = n695_q; // (signal)
  /* ni/MC_controller.vhd:87:31  */
  assign mode_change_idx_next = n609_o; // (signal)
  /* ni/MC_controller.vhd:88:10  */
  assign mode_idx_reg = n703_q; // (signal)
  /* ni/MC_controller.vhd:90:10  */
  assign mode_change_cnt_reg = n678_q; // (signal)
  /* ni/MC_controller.vhd:90:31  */
  assign mode_change_cnt_next = n610_o; // (signal)
  /* ni/MC_controller.vhd:90:53  */
  assign mode_change_cnt_int = n624_o; // (signal)
  /* ni/MC_controller.vhd:92:10  */
  assign mode_reg = n687_q; // (signal)
  /* ni/MC_controller.vhd:92:20  */
  assign mode_next = n611_o; // (signal)
  /* ni/MC_controller.vhd:94:10  */
  assign global_mode_change_idx = n643_o; // (signal)
  /* ni/MC_controller.vhd:94:34  */
  assign local_mode_change_idx = n613_o; // (signal)
  /* ni/MC_controller.vhd:96:10  */
  assign config_slv_error_next = n616_o; // (signal)
  /* ni/MC_controller.vhd:98:10  */
  assign read_reg = n679_q; // (signal)
  /* ni/MC_controller.vhd:98:20  */
  assign read_next = n726_o; // (signal)
  /* ni/MC_controller.vhd:100:27  */
  assign mode_changed_reg = n636_q; // (signal)
  /* ni/MC_controller.vhd:101:10  */
  assign stbl_min_reg = n715_q; // (signal)
  /* ni/MC_controller.vhd:103:10  */
  assign mc_tbl_addr = n558_o; // (signal)
  /* ni/MC_controller.vhd:124:31  */
  assign n556_o = n544_o[10:0];
  /* ni/MC_controller.vhd:124:60  */
  assign n558_o = n556_o - 11'b00000000010;
  /* ni/MC_controller.vhd:126:30  */
  assign n559_o = n544_o[14];
  /* ni/MC_controller.vhd:126:19  */
  assign n560_o = sel & n559_o;
  /* ni/MC_controller.vhd:128:17  */
  assign n561_o = n544_o[15];
  /* ni/MC_controller.vhd:128:20  */
  assign n562_o = ~n561_o;
  /* ni/MC_controller.vhd:129:26  */
  assign n563_o = n544_o[10:0];
  /* ni/MC_controller.vhd:131:11  */
  assign n565_o = n563_o == 11'b00000000000;
  /* ni/MC_controller.vhd:129:9  */
  always @*
    case (n565_o)
      1'b1: n568_o <= 1'b0;
      default: n568_o <= 1'b1;
    endcase
  assign n569_o = read_reg[1:0];
  /* ni/MC_controller.vhd:129:9  */
  always @*
    case (n565_o)
      1'b1: n570_o <= mode_idx_reg;
      default: n570_o <= n569_o;
    endcase
  /* ni/MC_controller.vhd:144:26  */
  assign n571_o = n544_o[10:0];
  /* ni/MC_controller.vhd:147:58  */
  assign n572_o = n544_o[17:16];
  /* ni/MC_controller.vhd:146:11  */
  assign n574_o = n571_o == 11'b00000000000;
  /* ni/MC_controller.vhd:151:8  */
  assign n576_o = n571_o == 11'b00000000001;
  assign n577_o = {n576_o, n574_o};
  /* ni/MC_controller.vhd:144:9  */
  always @*
    case (n577_o)
      2'b10: n578_o <= mode_change_idx_reg;
      2'b01: n578_o <= n572_o;
      default: n578_o <= mode_change_idx_reg;
    endcase
  /* ni/MC_controller.vhd:144:9  */
  always @*
    case (n577_o)
      2'b10: n579_o <= mode_change_cnt_reg;
      2'b01: n579_o <= mode_change_cnt_int;
      default: n579_o <= mode_change_cnt_reg;
    endcase
  /* ni/MC_controller.vhd:144:9  */
  always @*
    case (n577_o)
      2'b10: n582_o <= 1'b0;
      2'b01: n582_o <= 1'b1;
      default: n582_o <= 1'b0;
    endcase
  /* ni/MC_controller.vhd:144:9  */
  always @*
    case (n577_o)
      2'b10: n585_o <= 1'b0;
      2'b01: n585_o <= 1'b0;
      default: n585_o <= 1'b1;
    endcase
  /* ni/MC_controller.vhd:158:24  */
  assign n587_o = $unsigned(mc_tbl_addr) < $unsigned(11'b00000000100);
  /* ni/MC_controller.vhd:160:22  */
  assign n589_o = mc_tbl_addr[1:0];  // trunc
  /* ni/MC_controller.vhd:160:76  */
  assign n591_o = n544_o[23:16];
  /* ni/MC_controller.vhd:161:22  */
  assign n594_o = mc_tbl_addr[1:0];  // trunc
  /* ni/MC_controller.vhd:161:76  */
  assign n596_o = n544_o[39:32];
  /* ni/MC_controller.vhd:158:9  */
  assign n598_o = n587_o ? n770_o : mode_reg;
  /* ni/MC_controller.vhd:158:9  */
  assign n600_o = n587_o ? 1'b0 : n585_o;
  /* ni/MC_controller.vhd:128:7  */
  assign n601_o = n562_o ? mode_change_idx_reg : n578_o;
  /* ni/MC_controller.vhd:128:7  */
  assign n602_o = n562_o ? mode_change_cnt_reg : n579_o;
  /* ni/MC_controller.vhd:128:7  */
  assign n603_o = n562_o ? mode_reg : n598_o;
  /* ni/MC_controller.vhd:128:7  */
  assign n605_o = n562_o ? 1'b0 : n582_o;
  /* ni/MC_controller.vhd:128:7  */
  assign n606_o = n562_o ? n568_o : n600_o;
  assign n607_o = read_reg[1:0];
  /* ni/MC_controller.vhd:126:5  */
  assign n608_o = n619_o ? n570_o : n607_o;
  /* ni/MC_controller.vhd:126:5  */
  assign n609_o = n560_o ? n601_o : mode_change_idx_reg;
  /* ni/MC_controller.vhd:126:5  */
  assign n610_o = n560_o ? n602_o : mode_change_cnt_reg;
  /* ni/MC_controller.vhd:126:5  */
  assign n611_o = n560_o ? n603_o : mode_reg;
  /* ni/MC_controller.vhd:126:5  */
  assign n613_o = n560_o ? n605_o : 1'b0;
  /* ni/MC_controller.vhd:126:5  */
  assign n616_o = n560_o ? n606_o : 1'b0;
  /* ni/MC_controller.vhd:126:5  */
  assign n619_o = n560_o & n562_o;
  assign n620_o = read_reg[31:2];
  /* ni/MC_controller.vhd:212:49  */
  assign n624_o = n544_o[33:32];
  /* ni/MC_controller.vhd:223:11  */
  assign n629_o = global_mode_change_idx ? 1'b0 : mode_changed_reg;
  /* ni/MC_controller.vhd:221:11  */
  assign n631_o = local_mode_change_idx ? 1'b1 : n629_o;
  /* ni/MC_controller.vhd:218:9  */
  assign n633_o = reset ? 1'b0 : n631_o;
  /* ni/MC_controller.vhd:217:7  */
  always @(posedge clk)
    n636_q <= n633_o;
  /* ni/MC_controller.vhd:235:32  */
  assign n638_o = mode_change_cnt_reg == mc_p_cnt;
  /* ni/MC_controller.vhd:235:9  */
  assign n641_o = n638_o ? 1'b1 : 1'b0;
  /* ni/MC_controller.vhd:234:7  */
  assign n643_o = mode_changed_reg ? n641_o : 1'b0;
  /* ni/MC_controller.vhd:257:57  */
  assign n649_o = n776_o[7:0];
  /* ni/MC_controller.vhd:258:59  */
  assign n653_o = n782_o[15:8];
  /* ni/MC_controller.vhd:268:5  */
  assign n655_o = period_boundary ? stbl_min_next : stbl_min_reg;
  /* ni/MC_controller.vhd:281:7  */
  assign n660_o = reset ? 1'b0 : config_slv_error_next;
  /* ni/MC_controller.vhd:281:7  */
  assign n664_o = reset ? 2'b00 : mode_change_cnt_next;
  /* ni/MC_controller.vhd:281:7  */
  assign n666_o = reset ? 32'b00000000000000000000000000000000 : read_next;
  /* ni/MC_controller.vhd:280:5  */
  always @(posedge clk)
    n676_q <= n660_o;
  /* ni/MC_controller.vhd:280:5  */
  always @(posedge clk)
    n678_q <= n664_o;
  /* ni/MC_controller.vhd:280:5  */
  always @(posedge clk)
    n679_q <= n666_o;
  /* ni/MC_controller.vhd:302:7  */
  assign n684_o = reset ? 64'b0000000000000000000000000000000000000000000000000000000000000000 : mode_next;
  /* ni/MC_controller.vhd:301:5  */
  always @(posedge clk)
    n687_q <= n684_o;
  /* ni/MC_controller.vhd:324:9  */
  assign n690_o = local_mode_change_idx ? mode_change_idx_next : mode_change_idx_reg;
  /* ni/MC_controller.vhd:321:7  */
  assign n692_o = reset ? 2'b00 : n690_o;
  /* ni/MC_controller.vhd:320:5  */
  always @(posedge clk)
    n695_q <= n692_o;
  /* ni/MC_controller.vhd:338:9  */
  assign n698_o = global_mode_change_idx ? mode_change_idx_reg : mode_idx_reg;
  /* ni/MC_controller.vhd:335:7  */
  assign n700_o = reset ? 2'b00 : n698_o;
  /* ni/MC_controller.vhd:334:5  */
  always @(posedge clk)
    n703_q <= n700_o;
  /* ni/MC_controller.vhd:354:9  */
  assign n706_o = period_boundary ? stbl_min_next : stbl_min_reg;
  /* ni/MC_controller.vhd:350:7  */
  assign n709_o = reset ? 8'b00000000 : n706_o;
  /* ni/MC_controller.vhd:349:5  */
  always @(posedge clk)
    n715_q <= n709_o;
  /* ni/MC_controller.vhd:373:9  */
  assign n719_o = period_boundary ? stbl_maxp1_next : n724_q;
  /* ni/MC_controller.vhd:370:7  */
  assign n721_o = reset ? 8'b00000000 : n719_o;
  /* ni/MC_controller.vhd:369:5  */
  always @(posedge clk)
    n724_q <= n721_o;
  assign n726_o = {n620_o, n608_o};
  assign n728_o = {n676_q, read_reg};
  /* ni/MC_controller.vhd:160:13  */
  assign n729_o = n589_o[1];
  /* ni/MC_controller.vhd:160:13  */
  assign n730_o = ~n729_o;
  /* ni/MC_controller.vhd:160:13  */
  assign n731_o = n589_o[0];
  /* ni/MC_controller.vhd:160:13  */
  assign n732_o = ~n731_o;
  /* ni/MC_controller.vhd:160:13  */
  assign n733_o = n730_o & n732_o;
  /* ni/MC_controller.vhd:160:13  */
  assign n734_o = n730_o & n731_o;
  /* ni/MC_controller.vhd:160:13  */
  assign n735_o = n729_o & n732_o;
  /* ni/MC_controller.vhd:160:13  */
  assign n736_o = n729_o & n731_o;
  assign n737_o = mode_reg[7:0];
  /* ni/MC_controller.vhd:160:13  */
  assign n738_o = n733_o ? n591_o : n737_o;
  /* ni/MC_controller.vhd:349:5  */
  assign n739_o = mode_reg[15:8];
  assign n740_o = mode_reg[23:16];
  /* ni/MC_controller.vhd:160:13  */
  assign n741_o = n734_o ? n591_o : n740_o;
  assign n742_o = mode_reg[31:24];
  /* ni/MC_controller.vhd:354:9  */
  assign n743_o = mode_reg[39:32];
  /* ni/MC_controller.vhd:160:13  */
  assign n744_o = n735_o ? n591_o : n743_o;
  assign n745_o = mode_reg[47:40];
  /* ni/MC_controller.vhd:332:3  */
  assign n746_o = mode_reg[55:48];
  /* ni/MC_controller.vhd:160:13  */
  assign n747_o = n736_o ? n591_o : n746_o;
  /* ni/MC_controller.vhd:318:3  */
  assign n748_o = mode_reg[63:56];
  assign n749_o = {n748_o, n747_o, n745_o, n744_o, n742_o, n741_o, n739_o, n738_o};
  /* ni/MC_controller.vhd:161:13  */
  assign n750_o = n594_o[1];
  /* ni/MC_controller.vhd:161:13  */
  assign n751_o = ~n750_o;
  /* ni/MC_controller.vhd:161:13  */
  assign n752_o = n594_o[0];
  /* ni/MC_controller.vhd:161:13  */
  assign n753_o = ~n752_o;
  /* ni/MC_controller.vhd:161:13  */
  assign n754_o = n751_o & n753_o;
  /* ni/MC_controller.vhd:161:13  */
  assign n755_o = n751_o & n752_o;
  /* ni/MC_controller.vhd:161:13  */
  assign n756_o = n750_o & n753_o;
  /* ni/MC_controller.vhd:161:13  */
  assign n757_o = n750_o & n752_o;
  assign n758_o = n749_o[7:0];
  /* ni/MC_controller.vhd:281:7  */
  assign n759_o = n749_o[15:8];
  /* ni/MC_controller.vhd:161:13  */
  assign n760_o = n754_o ? n596_o : n759_o;
  /* ni/MC_controller.vhd:278:3  */
  assign n761_o = n749_o[23:16];
  assign n762_o = n749_o[31:24];
  /* ni/MC_controller.vhd:161:13  */
  assign n763_o = n755_o ? n596_o : n762_o;
  /* ni/MC_controller.vhd:258:33  */
  assign n764_o = n749_o[39:32];
  /* ni/MC_controller.vhd:257:31  */
  assign n765_o = n749_o[47:40];
  /* ni/MC_controller.vhd:161:13  */
  assign n766_o = n756_o ? n596_o : n765_o;
  assign n767_o = n749_o[55:48];
  /* ni/MC_controller.vhd:231:5  */
  assign n768_o = n749_o[63:56];
  /* ni/MC_controller.vhd:161:13  */
  assign n769_o = n757_o ? n596_o : n768_o;
  /* ni/MC_controller.vhd:215:5  */
  assign n770_o = {n769_o, n767_o, n766_o, n764_o, n763_o, n761_o, n760_o, n758_o};
  /* ni/MC_controller.vhd:161:23  */
  assign n771_o = mode_reg[15:0];
  /* ni/MC_controller.vhd:161:13  */
  assign n772_o = mode_reg[31:16];
  assign n773_o = mode_reg[47:32];
  assign n774_o = mode_reg[63:48];
  /* ni/MC_controller.vhd:257:30  */
  assign n775_o = mode_idx_reg[1:0];
  /* ni/MC_controller.vhd:257:30  */
  always @*
    case (n775_o)
      2'b00: n776_o <= n771_o;
      2'b01: n776_o <= n772_o;
      2'b10: n776_o <= n773_o;
      2'b11: n776_o <= n774_o;
    endcase
  /* ni/MC_controller.vhd:257:31  */
  assign n777_o = mode_reg[15:0];
  /* ni/MC_controller.vhd:257:30  */
  assign n778_o = mode_reg[31:16];
  /* ni/MC_controller.vhd:161:23  */
  assign n779_o = mode_reg[47:32];
  /* ni/MC_controller.vhd:160:23  */
  assign n780_o = mode_reg[63:48];
  /* ni/MC_controller.vhd:258:32  */
  assign n781_o = mode_idx_reg[1:0];
  /* ni/MC_controller.vhd:258:32  */
  always @*
    case (n781_o)
      2'b00: n782_o <= n777_o;
      2'b01: n782_o <= n778_o;
      2'b10: n782_o <= n779_o;
      2'b11: n782_o <= n780_o;
    endcase
endmodule

module tdm_controller_5ba93c9db0cff93f52b521d7420e43f6eda2784f
  (input  clk,
   input  reset,
   input  run,
   input  [13:0] config_addr,
   input  config_en,
   input  config_wr,
   input  [31:0] config_wdata,
   input  sel,
   input  [3:0] t2n,
   input  [7:0] stbl_min,
   input  [7:0] stbl_maxp1,
   output master_run,
   output [31:0] config_slv_rdata,
   output config_slv_error,
   output [7:0] stbl_idx,
   output stbl_idx_en,
   output period_boundary,
   output [1:0] mc_p_cnt);
  wire [47:0] n383_o;
  wire [31:0] n385_o;
  wire n386_o;
  wire [9:0] tdm_s_cnt_reg;
  wire [31:0] tdm_p_cnt_reg;
  wire [7:0] stbl_idx_reg;
  wire [7:0] stbl_idx_next;
  wire [3:0] time2next_reg;
  wire [31:0] clock_cnt_lo_reg;
  wire [1:0] mc_p_cnt_reg;
  wire [31:0] read_reg;
  wire [31:0] read_next;
  wire [31:0] clock_delay_reg;
  wire period_boundary_sig;
  wire stbl_idx_reset;
  wire stbl_idx_en_sig;
  wire t2n_ld_reg;
  wire [7:0] stbl_idx_inc;
  wire config_slv_error_next;
  wire run_reg;
  localparam n391_o = 1'b0;
  wire n396_o;
  wire n397_o;
  wire n398_o;
  wire n399_o;
  wire [10:0] n400_o;
  wire [30:0] n401_o;
  wire n403_o;
  wire n405_o;
  wire n407_o;
  wire n409_o;
  localparam [31:0] n410_o = 32'b00000000000000000000000000000000;
  wire [30:0] n411_o;
  wire n413_o;
  wire [4:0] n414_o;
  wire n415_o;
  wire n416_o;
  wire n417_o;
  wire n418_o;
  wire n419_o;
  reg n420_o;
  wire [8:0] n421_o;
  wire [8:0] n422_o;
  wire [8:0] n423_o;
  wire [8:0] n424_o;
  wire [8:0] n425_o;
  wire [8:0] n426_o;
  reg [8:0] n427_o;
  wire [21:0] n428_o;
  wire [21:0] n429_o;
  wire [21:0] n430_o;
  wire [21:0] n431_o;
  wire [21:0] n432_o;
  reg [21:0] n433_o;
  reg n439_o;
  wire [10:0] n440_o;
  wire [30:0] n441_o;
  wire n443_o;
  reg n446_o;
  wire [31:0] n447_o;
  wire [31:0] n448_o;
  wire n451_o;
  wire n452_o;
  wire n457_o;
  wire [7:0] n461_o;
  wire n464_o;
  wire n466_o;
  wire [4:0] n467_o;
  wire n469_o;
  wire n470_o;
  wire n472_o;
  wire n473_o;
  wire n474_o;
  wire n475_o;
  wire n476_o;
  wire n477_o;
  wire n478_o;
  wire n481_o;
  wire n482_o;
  wire n483_o;
  wire n484_o;
  wire n485_o;
  wire n487_o;
  wire n488_o;
  wire [7:0] n489_o;
  wire n493_o;
  wire [31:0] n495_o;
  wire n497_o;
  wire n498_o;
  reg n505_q;
  reg [31:0] n506_q;
  reg n507_q;
  reg n508_q;
  wire [1:0] n517_o;
  wire [1:0] n518_o;
  wire [1:0] n520_o;
  reg [1:0] n523_q;
  wire [3:0] n527_o;
  wire [3:0] n528_o;
  wire [3:0] n530_o;
  reg [3:0] n533_q;
  wire [7:0] n536_o;
  wire [7:0] n538_o;
  reg [7:0] n541_q;
  wire [32:0] n543_o;
  assign master_run = n391_o;
  assign config_slv_rdata = n385_o;
  assign config_slv_error = n386_o;
  assign stbl_idx = stbl_idx_next;
  assign stbl_idx_en = stbl_idx_en_sig;
  assign period_boundary = period_boundary_sig;
  assign mc_p_cnt = mc_p_cnt_reg;
  /* routers/synchronous/router.vhd:97:97  */
  assign n383_o = {config_wdata, config_wr, config_en, config_addr};
  /* routers/synchronous/router.vhd:96:9  */
  assign n385_o = n543_o[31:0];
  /* routers/synchronous/router.vhd:96:9  */
  assign n386_o = n543_o[32];
  /* ni/TDM_controller.vhd:84:10  */
  assign tdm_s_cnt_reg = 10'b0000000000; // (signal)
  /* ni/TDM_controller.vhd:85:10  */
  assign tdm_p_cnt_reg = 32'b00000000000000000000000000000000; // (signal)
  /* ni/TDM_controller.vhd:87:10  */
  assign stbl_idx_reg = n541_q; // (signal)
  /* ni/TDM_controller.vhd:88:10  */
  assign stbl_idx_next = n489_o; // (signal)
  /* ni/TDM_controller.vhd:89:10  */
  assign time2next_reg = n533_q; // (signal)
  /* ni/TDM_controller.vhd:165:42  */
  assign clock_cnt_lo_reg = 32'b00000000000000000000000000000000; // (signal)
  /* ni/TDM_controller.vhd:95:10  */
  assign mc_p_cnt_reg = n523_q; // (signal)
  /* ni/TDM_controller.vhd:105:10  */
  assign read_reg = n506_q; // (signal)
  /* ni/TDM_controller.vhd:105:20  */
  assign read_next = n448_o; // (signal)
  /* ni/TDM_controller.vhd:106:10  */
  assign clock_delay_reg = 32'b00000000000000000000000000000000; // (signal)
  /* ni/TDM_controller.vhd:108:10  */
  assign period_boundary_sig = n487_o; // (signal)
  /* ni/TDM_controller.vhd:109:10  */
  assign stbl_idx_reset = n485_o; // (signal)
  /* ni/TDM_controller.vhd:109:26  */
  assign stbl_idx_en_sig = n478_o; // (signal)
  /* ni/TDM_controller.vhd:109:43  */
  assign t2n_ld_reg = n507_q; // (signal)
  /* ni/TDM_controller.vhd:110:10  */
  assign stbl_idx_inc = n461_o; // (signal)
  /* ni/TDM_controller.vhd:112:10  */
  assign config_slv_error_next = n457_o; // (signal)
  /* ni/TDM_controller.vhd:117:10  */
  assign run_reg = n508_q; // (signal)
  /* ni/TDM_controller.vhd:154:30  */
  assign n396_o = n383_o[14];
  /* ni/TDM_controller.vhd:154:19  */
  assign n397_o = sel & n396_o;
  /* ni/TDM_controller.vhd:156:17  */
  assign n398_o = n383_o[15];
  /* ni/TDM_controller.vhd:156:20  */
  assign n399_o = ~n398_o;
  /* ni/TDM_controller.vhd:157:37  */
  assign n400_o = n383_o[10:0];
  /* ni/TDM_controller.vhd:157:15  */
  assign n401_o = {20'b0, n400_o};  //  uext
  /* ni/TDM_controller.vhd:158:11  */
  assign n403_o = n401_o == 31'b0000000000000000000000000000000;
  /* ni/TDM_controller.vhd:160:11  */
  assign n405_o = n401_o == 31'b0000000000000000000000000000001;
  /* ni/TDM_controller.vhd:162:11  */
  assign n407_o = n401_o == 31'b0000000000000000000000000000010;
  /* ni/TDM_controller.vhd:164:11  */
  assign n409_o = n401_o == 31'b0000000000000000000000000000011;
  assign n411_o = n410_o[31:1];
  /* ni/TDM_controller.vhd:167:11  */
  assign n413_o = n401_o == 31'b0000000000000000000000000000100;
  assign n414_o = {n413_o, n409_o, n407_o, n405_o, n403_o};
  assign n415_o = tdm_s_cnt_reg[0];
  assign n416_o = tdm_p_cnt_reg[0];
  assign n417_o = clock_delay_reg[0];
  assign n418_o = clock_cnt_lo_reg[0];
  assign n419_o = tdm_p_cnt_reg[0];
  /* ni/TDM_controller.vhd:157:9  */
  always @*
    case (n414_o)
      5'b10000: n420_o <= run;
      5'b01000: n420_o <= n418_o;
      5'b00100: n420_o <= n417_o;
      5'b00010: n420_o <= n416_o;
      5'b00001: n420_o <= n415_o;
      default: n420_o <= n419_o;
    endcase
  assign n421_o = tdm_s_cnt_reg[9:1];
  assign n422_o = tdm_p_cnt_reg[9:1];
  assign n423_o = clock_delay_reg[9:1];
  assign n424_o = clock_cnt_lo_reg[9:1];
  assign n425_o = n411_o[8:0];
  assign n426_o = tdm_p_cnt_reg[9:1];
  /* ni/TDM_controller.vhd:157:9  */
  always @*
    case (n414_o)
      5'b10000: n427_o <= n425_o;
      5'b01000: n427_o <= n424_o;
      5'b00100: n427_o <= n423_o;
      5'b00010: n427_o <= n422_o;
      5'b00001: n427_o <= n421_o;
      default: n427_o <= n426_o;
    endcase
  assign n428_o = tdm_p_cnt_reg[31:10];
  assign n429_o = clock_delay_reg[31:10];
  assign n430_o = clock_cnt_lo_reg[31:10];
  assign n431_o = n411_o[30:9];
  assign n432_o = tdm_p_cnt_reg[31:10];
  /* ni/TDM_controller.vhd:157:9  */
  always @*
    case (n414_o)
      5'b10000: n433_o <= n431_o;
      5'b01000: n433_o <= n430_o;
      5'b00100: n433_o <= n429_o;
      5'b00010: n433_o <= n428_o;
      5'b00001: n433_o <= n432_o;
      default: n433_o <= n432_o;
    endcase
  /* ni/TDM_controller.vhd:157:9  */
  always @*
    case (n414_o)
      5'b10000: n439_o <= 1'b0;
      5'b01000: n439_o <= 1'b0;
      5'b00100: n439_o <= 1'b0;
      5'b00010: n439_o <= 1'b0;
      5'b00001: n439_o <= 1'b0;
      default: n439_o <= 1'b1;
    endcase
  /* ni/TDM_controller.vhd:174:37  */
  assign n440_o = n383_o[10:0];
  /* ni/TDM_controller.vhd:174:15  */
  assign n441_o = {20'b0, n440_o};  //  uext
  /* ni/TDM_controller.vhd:175:11  */
  assign n443_o = n441_o == 31'b0000000000000000000000000000100;
  /* ni/TDM_controller.vhd:174:9  */
  always @*
    case (n443_o)
      1'b1: n446_o <= 1'b0;
      default: n446_o <= 1'b1;
    endcase
  assign n447_o = {n433_o, n427_o, n420_o};
  /* ni/TDM_controller.vhd:154:5  */
  assign n448_o = n452_o ? n447_o : tdm_p_cnt_reg;
  /* ni/TDM_controller.vhd:156:7  */
  assign n451_o = n399_o ? n439_o : n446_o;
  /* ni/TDM_controller.vhd:154:5  */
  assign n452_o = n397_o & n399_o;
  /* ni/TDM_controller.vhd:154:5  */
  assign n457_o = n397_o ? n451_o : 1'b0;
  /* ni/TDM_controller.vhd:194:32  */
  assign n461_o = stbl_idx_reg + 8'b00000001;
  /* ni/TDM_controller.vhd:198:49  */
  assign n464_o = time2next_reg == 4'b0001;
  /* ni/TDM_controller.vhd:198:74  */
  assign n466_o = time2next_reg == 4'b0000;
  /* ni/TDM_controller.vhd:198:97  */
  assign n467_o = {1'b0, time2next_reg};  //  uext
  /* ni/TDM_controller.vhd:198:97  */
  assign n469_o = n467_o == 5'b11111;
  /* ni/TDM_controller.vhd:198:79  */
  assign n470_o = n466_o | n469_o;
  /* ni/TDM_controller.vhd:198:118  */
  assign n472_o = t2n == 4'b0000;
  /* ni/TDM_controller.vhd:198:109  */
  assign n473_o = n470_o & n472_o;
  /* ni/TDM_controller.vhd:198:54  */
  assign n474_o = n464_o | n473_o;
  /* ni/TDM_controller.vhd:198:134  */
  assign n475_o = run != run_reg;
  /* ni/TDM_controller.vhd:198:125  */
  assign n476_o = n474_o | n475_o;
  /* ni/TDM_controller.vhd:198:147  */
  assign n477_o = n476_o & run;
  /* ni/TDM_controller.vhd:198:26  */
  assign n478_o = n477_o ? 1'b1 : 1'b0;
  /* ni/TDM_controller.vhd:201:46  */
  assign n481_o = stbl_idx_inc == stbl_maxp1;
  /* ni/TDM_controller.vhd:201:69  */
  assign n482_o = run != run_reg;
  /* ni/TDM_controller.vhd:201:60  */
  assign n483_o = n481_o | n482_o;
  /* ni/TDM_controller.vhd:201:82  */
  assign n484_o = n483_o & run;
  /* ni/TDM_controller.vhd:201:25  */
  assign n485_o = n484_o ? 1'b1 : 1'b0;
  /* ni/TDM_controller.vhd:205:41  */
  assign n487_o = stbl_idx_reset & stbl_idx_en_sig;
  /* ni/TDM_controller.vhd:208:53  */
  assign n488_o = ~stbl_idx_reset;
  /* ni/TDM_controller.vhd:208:33  */
  assign n489_o = n488_o ? stbl_idx_inc : stbl_min;
  /* ni/TDM_controller.vhd:220:7  */
  assign n493_o = reset ? 1'b0 : config_slv_error_next;
  /* ni/TDM_controller.vhd:220:7  */
  assign n495_o = reset ? 32'b00000000000000000000000000000000 : read_next;
  /* ni/TDM_controller.vhd:220:7  */
  assign n497_o = reset ? 1'b1 : stbl_idx_en_sig;
  /* ni/TDM_controller.vhd:220:7  */
  assign n498_o = reset ? run_reg : run;
  /* ni/TDM_controller.vhd:219:5  */
  always @(posedge clk)
    n505_q <= n493_o;
  /* ni/TDM_controller.vhd:219:5  */
  always @(posedge clk)
    n506_q <= n495_o;
  /* ni/TDM_controller.vhd:219:5  */
  always @(posedge clk)
    n507_q <= n497_o;
  /* ni/TDM_controller.vhd:219:5  */
  always @(posedge clk)
    n508_q <= n498_o;
  /* ni/TDM_controller.vhd:336:40  */
  assign n517_o = mc_p_cnt_reg + 2'b01;
  /* ni/TDM_controller.vhd:335:9  */
  assign n518_o = period_boundary_sig ? n517_o : mc_p_cnt_reg;
  /* ni/TDM_controller.vhd:332:7  */
  assign n520_o = reset ? 2'b00 : n518_o;
  /* ni/TDM_controller.vhd:331:5  */
  always @(posedge clk)
    n523_q <= n520_o;
  /* ni/TDM_controller.vhd:354:42  */
  assign n527_o = time2next_reg - 4'b0001;
  /* ni/TDM_controller.vhd:351:9  */
  assign n528_o = t2n_ld_reg ? t2n : n527_o;
  /* ni/TDM_controller.vhd:348:7  */
  assign n530_o = reset ? 4'b0000 : n528_o;
  /* ni/TDM_controller.vhd:347:5  */
  always @(posedge clk)
    n533_q <= n530_o;
  /* ni/TDM_controller.vhd:369:9  */
  assign n536_o = stbl_idx_en_sig ? stbl_idx_next : stbl_idx_reg;
  /* ni/TDM_controller.vhd:365:7  */
  assign n538_o = reset ? 8'b00000000 : n536_o;
  /* ni/TDM_controller.vhd:364:5  */
  always @(posedge clk)
    n541_q <= n538_o;
  assign n543_o = {n505_q, read_reg};
endmodule

module router
  (input  clk,
   input  reset,
   input  [179:0] inport_f,
   input  [4:0] outport_b,
   output [4:0] inport_b,
   output [179:0] outport_f);
  wire [3:0] sel0;
  wire [3:0] sel1;
  wire [3:0] sel2;
  wire [3:0] sel3;
  wire [3:0] sel4;
  wire [19:0] xbarsel;
  wire [19:0] xbarselnext;
  wire [179:0] xbarout;
  wire [179:0] xbaroutnext;
  wire [179:0] hpuout;
  wire [179:0] hpuoutnext;
  wire [179:0] hpuin;
  wire [35:0] n264_o;
  wire [35:0] port0_n265;
  wire [3:0] port0_n266;
  wire port0_outline_req;
  wire [34:0] port0_outline_data;
  wire [3:0] port0_sel;
  wire n267_o;
  wire [34:0] n268_o;
  wire [35:0] n269_o;
  wire [35:0] n274_o;
  wire [35:0] port1_n275;
  wire [3:0] port1_n276;
  wire port1_outline_req;
  wire [34:0] port1_outline_data;
  wire [3:0] port1_sel;
  wire n277_o;
  wire [34:0] n278_o;
  wire [35:0] n279_o;
  wire [35:0] n284_o;
  wire [35:0] port2_n285;
  wire [3:0] port2_n286;
  wire port2_outline_req;
  wire [34:0] port2_outline_data;
  wire [3:0] port2_sel;
  wire n287_o;
  wire [34:0] n288_o;
  wire [35:0] n289_o;
  wire [35:0] n294_o;
  wire [35:0] port3_n295;
  wire [3:0] port3_n296;
  wire port3_outline_req;
  wire [34:0] port3_outline_data;
  wire [3:0] port3_sel;
  wire n297_o;
  wire [34:0] n298_o;
  wire [35:0] n299_o;
  wire [35:0] n304_o;
  wire [35:0] port4_n305;
  wire [3:0] port4_n306;
  wire port4_outline_req;
  wire [34:0] port4_outline_data;
  wire [3:0] port4_sel;
  wire n307_o;
  wire [34:0] n308_o;
  wire [35:0] n309_o;
  wire [7:0] n314_o;
  wire [11:0] n315_o;
  wire [15:0] n316_o;
  wire [19:0] n317_o;
  wire [179:0] xbarinst_n318;
  wire [179:0] xbarinst_outport;
  wire [179:0] n369_o;
  wire [179:0] n371_o;
  wire [179:0] n373_o;
  reg [19:0] n376_q;
  reg [179:0] n377_q;
  reg [179:0] n378_q;
  reg [179:0] n379_q;
  wire [179:0] n380_o;
  localparam [4:0] n381_o = 5'bZ;
  assign inport_b = n381_o;
  assign outport_f = xbarout;
  /* routers/synchronous/router.vhd:78:8  */
  assign sel0 = port0_n266; // (signal)
  /* routers/synchronous/router.vhd:78:14  */
  assign sel1 = port1_n276; // (signal)
  /* routers/synchronous/router.vhd:78:20  */
  assign sel2 = port2_n286; // (signal)
  /* routers/synchronous/router.vhd:78:26  */
  assign sel3 = port3_n296; // (signal)
  /* routers/synchronous/router.vhd:78:32  */
  assign sel4 = port4_n306; // (signal)
  /* routers/synchronous/router.vhd:81:8  */
  assign xbarsel = n376_q; // (signal)
  /* routers/synchronous/router.vhd:81:17  */
  assign xbarselnext = n317_o; // (signal)
  /* routers/synchronous/router.vhd:82:8  */
  assign xbarout = n377_q; // (signal)
  /* routers/synchronous/router.vhd:82:17  */
  assign xbaroutnext = xbarinst_n318; // (signal)
  /* routers/synchronous/router.vhd:83:8  */
  assign hpuout = n378_q; // (signal)
  /* routers/synchronous/router.vhd:84:8  */
  assign hpuoutnext = n380_o; // (signal)
  /* routers/synchronous/router.vhd:85:8  */
  assign hpuin = n379_q; // (signal)
  /* routers/synchronous/router.vhd:89:63  */
  assign n264_o = hpuin[35:0];
  /* routers/synchronous/router.vhd:89:77  */
  assign port0_n265 = n269_o; // (signal)
  /* routers/synchronous/router.vhd:89:97  */
  assign port0_n266 = port0_sel; // (signal)
  /* routers/synchronous/router.vhd:88:9  */
  hpu port0 (
    .clk(clk),
    .reset(reset),
    .inline_req(n267_o),
    .inline_data(n268_o),
    .outline_req(port0_outline_req),
    .outline_data(port0_outline_data),
    .sel(port0_sel));
  /* ni/network_interface.vhd:362:32  */
  assign n267_o = n264_o[0];
  /* ni/network_interface.vhd:360:31  */
  assign n268_o = n264_o[35:1];
  /* ni/network_interface.vhd:354:9  */
  assign n269_o = {port0_outline_data, port0_outline_req};
  /* routers/synchronous/router.vhd:91:63  */
  assign n274_o = hpuin[71:36];
  /* routers/synchronous/router.vhd:91:77  */
  assign port1_n275 = n279_o; // (signal)
  /* routers/synchronous/router.vhd:91:97  */
  assign port1_n276 = port1_sel; // (signal)
  /* routers/synchronous/router.vhd:90:9  */
  hpu port1 (
    .clk(clk),
    .reset(reset),
    .inline_req(n277_o),
    .inline_data(n278_o),
    .outline_req(port1_outline_req),
    .outline_data(port1_outline_data),
    .sel(port1_sel));
  /* ni/network_interface.vhd:341:9  */
  assign n277_o = n274_o[0];
  /* ni/network_interface.vhd:341:9  */
  assign n278_o = n274_o[35:1];
  /* ni/network_interface.vhd:341:9  */
  assign n279_o = {port1_outline_data, port1_outline_req};
  /* routers/synchronous/router.vhd:93:63  */
  assign n284_o = hpuin[107:72];
  /* routers/synchronous/router.vhd:93:77  */
  assign port2_n285 = n289_o; // (signal)
  /* routers/synchronous/router.vhd:93:97  */
  assign port2_n286 = port2_sel; // (signal)
  /* routers/synchronous/router.vhd:92:9  */
  hpu port2 (
    .clk(clk),
    .reset(reset),
    .inline_req(n287_o),
    .inline_data(n288_o),
    .outline_req(port2_outline_req),
    .outline_data(port2_outline_data),
    .sel(port2_sel));
  /* ni/network_interface.vhd:317:28  */
  assign n287_o = n284_o[0];
  /* ni/network_interface.vhd:316:24  */
  assign n288_o = n284_o[35:1];
  /* ni/network_interface.vhd:315:28  */
  assign n289_o = {port2_outline_data, port2_outline_req};
  /* routers/synchronous/router.vhd:95:63  */
  assign n294_o = hpuin[143:108];
  /* routers/synchronous/router.vhd:95:77  */
  assign port3_n295 = n299_o; // (signal)
  /* routers/synchronous/router.vhd:95:97  */
  assign port3_n296 = port3_sel; // (signal)
  /* routers/synchronous/router.vhd:94:9  */
  hpu port3 (
    .clk(clk),
    .reset(reset),
    .inline_req(n297_o),
    .inline_data(n298_o),
    .outline_req(port3_outline_req),
    .outline_data(port3_outline_data),
    .sel(port3_sel));
  /* ni/network_interface.vhd:301:25  */
  assign n297_o = n294_o[0];
  /* ni/network_interface.vhd:300:27  */
  assign n298_o = n294_o[35:1];
  /* ni/network_interface.vhd:299:23  */
  assign n299_o = {port3_outline_data, port3_outline_req};
  /* routers/synchronous/router.vhd:97:63  */
  assign n304_o = hpuin[179:144];
  /* routers/synchronous/router.vhd:97:77  */
  assign port4_n305 = n309_o; // (signal)
  /* routers/synchronous/router.vhd:97:97  */
  assign port4_n306 = port4_sel; // (signal)
  /* routers/synchronous/router.vhd:96:9  */
  hpu port4 (
    .clk(clk),
    .reset(reset),
    .inline_req(n307_o),
    .inline_data(n308_o),
    .outline_req(port4_outline_req),
    .outline_data(port4_outline_data),
    .sel(port4_sel));
  /* ni/network_interface.vhd:284:9  */
  assign n307_o = n304_o[0];
  /* ni/network_interface.vhd:279:29  */
  assign n308_o = n304_o[35:1];
  /* ni/network_interface.vhd:278:36  */
  assign n309_o = {port4_outline_data, port4_outline_req};
  /* routers/synchronous/router.vhd:99:29  */
  assign n314_o = {sel4, sel3};
  /* routers/synchronous/router.vhd:99:36  */
  assign n315_o = {n314_o, sel2};
  /* routers/synchronous/router.vhd:99:43  */
  assign n316_o = {n315_o, sel1};
  /* routers/synchronous/router.vhd:99:50  */
  assign n317_o = {n316_o, sel0};
  /* routers/synchronous/router.vhd:102:74  */
  assign xbarinst_n318 = xbarinst_outport; // (signal)
  /* routers/synchronous/router.vhd:101:9  */
  xbar xbarinst (
    .func(xbarsel),
    .inport(hpuout),
    .outport(xbarinst_outport));
  assign n369_o = {35'b00000000000000000000000000000000000, 1'b0, 35'b00000000000000000000000000000000000, 1'b0, 35'b00000000000000000000000000000000000, 1'b0, 35'b00000000000000000000000000000000000, 1'b0, 35'b00000000000000000000000000000000000, 1'b0};
  assign n371_o = {35'b00000000000000000000000000000000000, 1'b0, 35'b00000000000000000000000000000000000, 1'b0, 35'b00000000000000000000000000000000000, 1'b0, 35'b00000000000000000000000000000000000, 1'b0, 35'b00000000000000000000000000000000000, 1'b0};
  assign n373_o = {35'b00000000000000000000000000000000000, 1'b0, 35'b00000000000000000000000000000000000, 1'b0, 35'b00000000000000000000000000000000000, 1'b0, 35'b00000000000000000000000000000000000, 1'b0, 35'b00000000000000000000000000000000000, 1'b0};
  /* routers/synchronous/router.vhd:113:17  */
  always @(posedge clk or posedge reset)
    if (reset)
      n376_q <= 20'b00000000000000000000;
    else
      n376_q <= xbarselnext;
  /* routers/synchronous/router.vhd:113:17  */
  always @(posedge clk or posedge reset)
    if (reset)
      n377_q <= n369_o;
    else
      n377_q <= xbaroutnext;
  /* routers/synchronous/router.vhd:113:17  */
  always @(posedge clk or posedge reset)
    if (reset)
      n378_q <= n371_o;
    else
      n378_q <= hpuoutnext;
  /* routers/synchronous/router.vhd:113:17  */
  always @(posedge clk or posedge reset)
    if (reset)
      n379_q <= n373_o;
    else
      n379_q <= inport_f;
  /* routers/synchronous/router.vhd:108:17  */
  assign n380_o = {port4_n305, port3_n295, port2_n285, port1_n275, port0_n265};
endmodule

module network_interface_5ba93c9db0cff93f52b521d7420e43f6eda2784f
  (input  clk,
   input  reset,
   input  run,
   input  supervisor,
   input  [2:0] ocp_config_m_mcmd,
   input  [31:0] ocp_config_m_maddr,
   input  [31:0] ocp_config_m_mdata,
   input  [3:0] ocp_config_m_mbyteen,
   input  ocp_config_m_mrespaccept,
   input  [63:0] spm_slv_rdata,
   input  spm_slv_error,
   input  [34:0] pkt_in,
   output master_run,
   output [1:0] ocp_config_s_sresp,
   output [31:0] ocp_config_s_sdata,
   output ocp_config_s_scmdaccept,
   output data_irq,
   output config_irq,
   output [13:0] spm_addr,
   output [1:0] spm_en,
   output spm_wr,
   output [63:0] spm_wdata,
   output [34:0] pkt_out);
  wire [71:0] n71_o;
  wire [1:0] n73_o;
  wire [31:0] n74_o;
  wire n75_o;
  wire [64:0] n78_o;
  wire [13:0] n80_o;
  wire [1:0] n81_o;
  wire n82_o;
  wire [63:0] n83_o;
  wire [47:0] config;
  wire [32:0] tdm_ctrl;
  wire [32:0] sched_tbl;
  wire [32:0] dma_tbl;
  wire [32:0] mc_ctrl;
  wire tdm_ctrl_sel;
  wire sched_tbl_sel;
  wire dma_tbl_sel;
  wire mc_ctrl_sel;
  wire [7:0] stbl_idx;
  wire stbl_idx_en;
  wire [3:0] t2n;
  wire [15:0] route;
  wire [3:0] pkt_len;
  wire [5:0] dma_num;
  wire dma_en;
  wire period_boundary;
  wire [7:0] stbl_min;
  wire [7:0] stbl_maxp1;
  wire [80:0] tx_spm;
  wire [80:0] rx_spm;
  wire [64:0] tx_spm_slv;
  wire [13:0] irq_fifo_data;
  wire irq_fifo_data_valid;
  wire irq_fifo_irq_valid;
  wire [47:0] config_unit_master;
  wire [32:0] irq_if_fifo;
  wire irq_if_fifo_sel;
  wire mc;
  wire [1:0] mc_idx;
  wire [1:0] mc_p_cnt;
  wire [1:0] mc_p;
  wire tdmctrl_n85;
  wire [32:0] tdmctrl_n86;
  wire [7:0] tdmctrl_n87;
  wire tdmctrl_n88;
  wire tdmctrl_n89;
  wire [1:0] tdmctrl_n90;
  wire tdmctrl_master_run;
  wire [31:0] tdmctrl_config_slv_rdata;
  wire tdmctrl_config_slv_error;
  wire [7:0] tdmctrl_stbl_idx;
  wire tdmctrl_stbl_idx_en;
  wire tdmctrl_period_boundary;
  wire [1:0] tdmctrl_mc_p_cnt;
  wire [13:0] n92_o;
  wire n93_o;
  wire n94_o;
  wire [31:0] n95_o;
  wire [32:0] n96_o;
  wire [32:0] mcctrl_n108;
  wire [7:0] mcctrl_n109;
  wire [7:0] mcctrl_n110;
  wire mcctrl_n111;
  wire [1:0] mcctrl_n112;
  wire [1:0] mcctrl_n113;
  wire [31:0] mcctrl_config_slv_rdata;
  wire mcctrl_config_slv_error;
  wire [7:0] mcctrl_stbl_min;
  wire [7:0] mcctrl_stbl_maxp1;
  wire mcctrl_mc;
  wire [1:0] mcctrl_mc_idx;
  wire [1:0] mcctrl_mc_p;
  wire [13:0] n114_o;
  wire n115_o;
  wire n116_o;
  wire [31:0] n117_o;
  wire [32:0] n118_o;
  wire [32:0] schedtbl_n131;
  wire [15:0] schedtbl_n132;
  wire [3:0] schedtbl_n133;
  wire [3:0] schedtbl_n134;
  wire [5:0] schedtbl_n135;
  wire schedtbl_n136;
  wire [31:0] schedtbl_config_slv_rdata;
  wire schedtbl_config_slv_error;
  wire [15:0] schedtbl_route;
  wire [3:0] schedtbl_pkt_len;
  wire [3:0] schedtbl_t2n;
  wire [5:0] schedtbl_dma_num;
  wire schedtbl_dma_en;
  wire [13:0] n137_o;
  wire n138_o;
  wire n139_o;
  wire [31:0] n140_o;
  wire [32:0] n141_o;
  wire [32:0] pktman_n154;
  wire [80:0] pktman_n155;
  wire [34:0] pktman_n156;
  wire [31:0] pktman_config_slv_rdata;
  wire pktman_config_slv_error;
  wire [13:0] pktman_spm_addr;
  wire [1:0] pktman_spm_en;
  wire pktman_spm_wr;
  wire [63:0] pktman_spm_wdata;
  wire [34:0] pktman_pkt_out;
  wire [13:0] n157_o;
  wire n158_o;
  wire n159_o;
  wire [31:0] n160_o;
  wire [32:0] n161_o;
  wire [80:0] n163_o;
  wire [63:0] n165_o;
  wire n166_o;
  wire [80:0] rxunit_n171;
  wire [47:0] rxunit_n172;
  wire [13:0] rxunit_n173;
  wire rxunit_n174;
  wire rxunit_n175;
  wire [13:0] rxunit_spm_addr;
  wire [1:0] rxunit_spm_en;
  wire rxunit_spm_wr;
  wire [63:0] rxunit_spm_wdata;
  wire [13:0] rxunit_config_addr;
  wire rxunit_config_en;
  wire rxunit_config_wr;
  wire [31:0] rxunit_config_wdata;
  wire [13:0] rxunit_irq_fifo_data;
  wire rxunit_irq_fifo_data_valid;
  wire rxunit_irq_fifo_irq_valid;
  wire [80:0] n176_o;
  wire [47:0] n178_o;
  wire [32:0] irqfifo_n188;
  wire irqfifo_n189;
  wire irqfifo_n190;
  wire [31:0] irqfifo_config_slv_rdata;
  wire irqfifo_config_slv_error;
  wire irqfifo_irq_irq_sig;
  wire irqfifo_irq_data_sig;
  wire [13:0] n191_o;
  wire n192_o;
  wire n193_o;
  wire [31:0] n194_o;
  wire [32:0] n195_o;
  wire [80:0] spmbus_n202;
  wire [64:0] spmbus_n203;
  wire [13:0] spmbus_spm_addr;
  wire [1:0] spmbus_spm_en;
  wire spmbus_spm_wr;
  wire [63:0] spmbus_spm_wdata;
  wire [63:0] spmbus_tx_spm_slv_rdata;
  wire spmbus_tx_spm_slv_error;
  wire [63:0] n204_o;
  wire n205_o;
  wire [80:0] n206_o;
  wire [64:0] n208_o;
  wire [13:0] n210_o;
  wire [1:0] n211_o;
  wire n212_o;
  wire [63:0] n213_o;
  wire [13:0] n214_o;
  wire [1:0] n215_o;
  wire n216_o;
  wire [63:0] n217_o;
  wire [34:0] configbus_n220;
  wire [47:0] configbus_n221;
  wire configbus_n222;
  wire configbus_n223;
  wire configbus_n224;
  wire configbus_n225;
  wire configbus_n226;
  wire [1:0] configbus_ocp_config_s_sresp;
  wire [31:0] configbus_ocp_config_s_sdata;
  wire configbus_ocp_config_s_scmdaccept;
  wire [13:0] configbus_config_addr;
  wire configbus_config_en;
  wire configbus_config_wr;
  wire [31:0] configbus_config_wdata;
  wire configbus_tdm_ctrl_sel;
  wire configbus_sched_tbl_sel;
  wire configbus_dma_tbl_sel;
  wire configbus_mc_ctrl_sel;
  wire configbus_irq_unit_fifo_sel;
  wire [2:0] n227_o;
  wire [31:0] n228_o;
  wire [31:0] n229_o;
  wire [3:0] n230_o;
  wire n231_o;
  wire [34:0] n232_o;
  wire [13:0] n234_o;
  wire n235_o;
  wire n236_o;
  wire [31:0] n237_o;
  wire [47:0] n238_o;
  wire [31:0] n240_o;
  wire n241_o;
  wire [31:0] n243_o;
  wire n244_o;
  wire [31:0] n246_o;
  wire n247_o;
  wire [31:0] n249_o;
  wire n250_o;
  wire [31:0] n252_o;
  wire n253_o;
  assign master_run = tdmctrl_n85;
  assign ocp_config_s_sresp = n73_o;
  assign ocp_config_s_sdata = n74_o;
  assign ocp_config_s_scmdaccept = n75_o;
  assign data_irq = irqfifo_n190;
  assign config_irq = irqfifo_n189;
  assign spm_addr = n80_o;
  assign spm_en = n81_o;
  assign spm_wr = n82_o;
  assign spm_wdata = n83_o;
  assign pkt_out = pktman_n156;
  /* noc/synchronous/noc_node.vhd:127:18  */
  assign n71_o = {ocp_config_m_mrespaccept, ocp_config_m_mbyteen, ocp_config_m_mdata, ocp_config_m_maddr, ocp_config_m_mcmd};
  /* noc/synchronous/noc_node.vhd:117:22  */
  assign n73_o = configbus_n220[1:0];
  /* noc/synchronous/noc_node.vhd:116:20  */
  assign n74_o = configbus_n220[33:2];
  /* noc/synchronous/noc_node.vhd:115:23  */
  assign n75_o = configbus_n220[34];
  /* noc/synchronous/noc_node.vhd:82:5  */
  assign n78_o = {spm_slv_error, spm_slv_rdata};
  /* noc/synchronous/noc_node.vhd:78:5  */
  assign n80_o = spmbus_n202[13:0];
  /* noc/synchronous/noc_node.vhd:75:5  */
  assign n81_o = spmbus_n202[15:14];
  /* noc/synchronous/noc_node.vhd:73:5  */
  assign n82_o = spmbus_n202[16];
  /* noc/synchronous/noc_node.vhd:71:5  */
  assign n83_o = spmbus_n202[80:17];
  /* ni/network_interface.vhd:227:8  */
  assign config = configbus_n221; // (signal)
  /* ni/network_interface.vhd:229:8  */
  assign tdm_ctrl = tdmctrl_n86; // (signal)
  /* ni/network_interface.vhd:229:18  */
  assign sched_tbl = schedtbl_n131; // (signal)
  /* ni/network_interface.vhd:229:29  */
  assign dma_tbl = pktman_n154; // (signal)
  /* ni/network_interface.vhd:229:38  */
  assign mc_ctrl = mcctrl_n108; // (signal)
  /* ni/network_interface.vhd:230:8  */
  assign tdm_ctrl_sel = configbus_n222; // (signal)
  /* ni/network_interface.vhd:230:22  */
  assign sched_tbl_sel = configbus_n223; // (signal)
  /* ni/network_interface.vhd:230:37  */
  assign dma_tbl_sel = configbus_n224; // (signal)
  /* ni/network_interface.vhd:230:50  */
  assign mc_ctrl_sel = configbus_n225; // (signal)
  /* ni/network_interface.vhd:231:8  */
  assign stbl_idx = tdmctrl_n87; // (signal)
  /* ni/network_interface.vhd:232:8  */
  assign stbl_idx_en = tdmctrl_n88; // (signal)
  /* ni/network_interface.vhd:233:8  */
  assign t2n = schedtbl_n134; // (signal)
  /* ni/network_interface.vhd:235:8  */
  assign route = schedtbl_n132; // (signal)
  /* ni/network_interface.vhd:236:8  */
  assign pkt_len = schedtbl_n133; // (signal)
  /* ni/network_interface.vhd:237:8  */
  assign dma_num = schedtbl_n135; // (signal)
  /* ni/network_interface.vhd:238:8  */
  assign dma_en = schedtbl_n136; // (signal)
  /* ni/network_interface.vhd:240:8  */
  assign period_boundary = tdmctrl_n89; // (signal)
  /* ni/network_interface.vhd:241:8  */
  assign stbl_min = mcctrl_n109; // (signal)
  /* ni/network_interface.vhd:242:8  */
  assign stbl_maxp1 = mcctrl_n110; // (signal)
  /* ni/network_interface.vhd:244:8  */
  assign tx_spm = pktman_n155; // (signal)
  /* ni/network_interface.vhd:244:16  */
  assign rx_spm = rxunit_n171; // (signal)
  /* ni/network_interface.vhd:245:8  */
  assign tx_spm_slv = spmbus_n203; // (signal)
  /* ni/network_interface.vhd:247:8  */
  assign irq_fifo_data = rxunit_n173; // (signal)
  /* ni/network_interface.vhd:248:8  */
  assign irq_fifo_data_valid = rxunit_n174; // (signal)
  /* ni/network_interface.vhd:248:29  */
  assign irq_fifo_irq_valid = rxunit_n175; // (signal)
  /* ni/network_interface.vhd:250:8  */
  assign config_unit_master = rxunit_n172; // (signal)
  /* ni/network_interface.vhd:251:8  */
  assign irq_if_fifo = irqfifo_n188; // (signal)
  /* ni/network_interface.vhd:252:8  */
  assign irq_if_fifo_sel = configbus_n226; // (signal)
  /* ni/network_interface.vhd:254:8  */
  assign mc = mcctrl_n111; // (signal)
  /* ni/network_interface.vhd:255:8  */
  assign mc_idx = mcctrl_n112; // (signal)
  /* ni/network_interface.vhd:256:8  */
  assign mc_p_cnt = tdmctrl_n90; // (signal)
  /* ni/network_interface.vhd:257:8  */
  assign mc_p = mcctrl_n113; // (signal)
  /* ni/network_interface.vhd:271:31  */
  assign tdmctrl_n85 = tdmctrl_master_run; // (signal)
  /* ni/network_interface.vhd:274:31  */
  assign tdmctrl_n86 = n96_o; // (signal)
  /* ni/network_interface.vhd:275:29  */
  assign tdmctrl_n87 = tdmctrl_stbl_idx; // (signal)
  /* ni/network_interface.vhd:276:32  */
  assign tdmctrl_n88 = tdmctrl_stbl_idx_en; // (signal)
  /* ni/network_interface.vhd:278:36  */
  assign tdmctrl_n89 = tdmctrl_period_boundary; // (signal)
  /* ni/network_interface.vhd:279:29  */
  assign tdmctrl_n90 = tdmctrl_mc_p_cnt; // (signal)
  /* ni/network_interface.vhd:263:9  */
  tdm_controller_5ba93c9db0cff93f52b521d7420e43f6eda2784f tdmctrl (
    .clk(clk),
    .reset(reset),
    .run(run),
    .config_addr(n92_o),
    .config_en(n93_o),
    .config_wr(n94_o),
    .config_wdata(n95_o),
    .sel(tdm_ctrl_sel),
    .t2n(t2n),
    .stbl_min(stbl_min),
    .stbl_maxp1(stbl_maxp1),
    .master_run(tdmctrl_master_run),
    .config_slv_rdata(tdmctrl_config_slv_rdata),
    .config_slv_error(tdmctrl_config_slv_error),
    .stbl_idx(tdmctrl_stbl_idx),
    .stbl_idx_en(tdmctrl_stbl_idx_en),
    .period_boundary(tdmctrl_period_boundary),
    .mc_p_cnt(tdmctrl_mc_p_cnt));
  assign n92_o = config[13:0];
  assign n93_o = config[14];
  assign n94_o = config[15];
  assign n95_o = config[47:16];
  assign n96_o = {tdmctrl_config_slv_error, tdmctrl_config_slv_rdata};
  /* ni/network_interface.vhd:294:31  */
  assign mcctrl_n108 = n118_o; // (signal)
  /* ni/network_interface.vhd:297:29  */
  assign mcctrl_n109 = mcctrl_stbl_min; // (signal)
  /* ni/network_interface.vhd:298:31  */
  assign mcctrl_n110 = mcctrl_stbl_maxp1; // (signal)
  /* ni/network_interface.vhd:299:23  */
  assign mcctrl_n111 = mcctrl_mc; // (signal)
  /* ni/network_interface.vhd:300:27  */
  assign mcctrl_n112 = mcctrl_mc_idx; // (signal)
  /* ni/network_interface.vhd:301:25  */
  assign mcctrl_n113 = mcctrl_mc_p; // (signal)
  /* ni/network_interface.vhd:284:9  */
  mc_controller_5ba93c9db0cff93f52b521d7420e43f6eda2784f mcctrl (
    .clk(clk),
    .reset(reset),
    .run(run),
    .config_addr(n114_o),
    .config_en(n115_o),
    .config_wr(n116_o),
    .config_wdata(n117_o),
    .sel(mc_ctrl_sel),
    .period_boundary(period_boundary),
    .mc_p_cnt(mc_p_cnt),
    .config_slv_rdata(mcctrl_config_slv_rdata),
    .config_slv_error(mcctrl_config_slv_error),
    .stbl_min(mcctrl_stbl_min),
    .stbl_maxp1(mcctrl_stbl_maxp1),
    .mc(mcctrl_mc),
    .mc_idx(mcctrl_mc_idx),
    .mc_p(mcctrl_mc_p));
  assign n114_o = config[13:0];
  assign n115_o = config[14];
  assign n116_o = config[15];
  assign n117_o = config[47:16];
  assign n118_o = {mcctrl_config_slv_error, mcctrl_config_slv_rdata};
  /* ni/network_interface.vhd:311:31  */
  assign schedtbl_n131 = n141_o; // (signal)
  /* ni/network_interface.vhd:314:26  */
  assign schedtbl_n132 = schedtbl_route; // (signal)
  /* ni/network_interface.vhd:315:28  */
  assign schedtbl_n133 = schedtbl_pkt_len; // (signal)
  /* ni/network_interface.vhd:316:24  */
  assign schedtbl_n134 = schedtbl_t2n; // (signal)
  /* ni/network_interface.vhd:317:28  */
  assign schedtbl_n135 = schedtbl_dma_num; // (signal)
  /* ni/network_interface.vhd:318:27  */
  assign schedtbl_n136 = schedtbl_dma_en; // (signal)
  /* ni/network_interface.vhd:305:9  */
  schedule_table schedtbl (
    .clk(clk),
    .reset(reset),
    .config_addr(n137_o),
    .config_en(n138_o),
    .config_wr(n139_o),
    .config_wdata(n140_o),
    .sel(sched_tbl_sel),
    .stbl_idx(stbl_idx),
    .stbl_idx_en(stbl_idx_en),
    .config_slv_rdata(schedtbl_config_slv_rdata),
    .config_slv_error(schedtbl_config_slv_error),
    .route(schedtbl_route),
    .pkt_len(schedtbl_pkt_len),
    .t2n(schedtbl_t2n),
    .dma_num(schedtbl_dma_num),
    .dma_en(schedtbl_dma_en));
  assign n137_o = config[13:0];
  assign n138_o = config[14];
  assign n139_o = config[15];
  assign n140_o = config[47:16];
  assign n141_o = {schedtbl_config_slv_error, schedtbl_config_slv_rdata};
  /* ni/network_interface.vhd:327:31  */
  assign pktman_n154 = n161_o; // (signal)
  /* ni/network_interface.vhd:328:24  */
  assign pktman_n155 = n163_o; // (signal)
  /* ni/network_interface.vhd:337:28  */
  assign pktman_n156 = pktman_pkt_out; // (signal)
  /* ni/network_interface.vhd:321:9  */
  packet_manager pktman (
    .clk(clk),
    .reset(reset),
    .config_addr(n157_o),
    .config_en(n158_o),
    .config_wr(n159_o),
    .config_wdata(n160_o),
    .sel(dma_tbl_sel),
    .spm_slv_rdata(n165_o),
    .spm_slv_error(n166_o),
    .dma_num(dma_num),
    .dma_en(dma_en),
    .route(route),
    .mc(mc),
    .mc_idx(mc_idx),
    .mc_p(mc_p),
    .pkt_len(pkt_len),
    .config_slv_rdata(pktman_config_slv_rdata),
    .config_slv_error(pktman_config_slv_error),
    .spm_addr(pktman_spm_addr),
    .spm_en(pktman_spm_en),
    .spm_wr(pktman_spm_wr),
    .spm_wdata(pktman_spm_wdata),
    .pkt_out(pktman_pkt_out));
  assign n157_o = config[13:0];
  assign n158_o = config[14];
  assign n159_o = config[15];
  assign n160_o = config[47:16];
  assign n161_o = {pktman_config_slv_error, pktman_config_slv_rdata};
  assign n163_o = {pktman_spm_wdata, pktman_spm_wr, pktman_spm_en, pktman_spm_addr};
  assign n165_o = tx_spm_slv[63:0];
  assign n166_o = tx_spm_slv[64];
  /* ni/network_interface.vhd:345:24  */
  assign rxunit_n171 = n176_o; // (signal)
  /* ni/network_interface.vhd:346:27  */
  assign rxunit_n172 = n178_o; // (signal)
  /* ni/network_interface.vhd:347:34  */
  assign rxunit_n173 = rxunit_irq_fifo_data; // (signal)
  /* ni/network_interface.vhd:348:40  */
  assign rxunit_n174 = rxunit_irq_fifo_data_valid; // (signal)
  /* ni/network_interface.vhd:349:39  */
  assign rxunit_n175 = rxunit_irq_fifo_irq_valid; // (signal)
  /* ni/network_interface.vhd:341:9  */
  rx_unit rxunit (
    .clk(clk),
    .reset(reset),
    .pkt_in(pkt_in),
    .spm_addr(rxunit_spm_addr),
    .spm_en(rxunit_spm_en),
    .spm_wr(rxunit_spm_wr),
    .spm_wdata(rxunit_spm_wdata),
    .config_addr(rxunit_config_addr),
    .config_en(rxunit_config_en),
    .config_wr(rxunit_config_wr),
    .config_wdata(rxunit_config_wdata),
    .irq_fifo_data(rxunit_irq_fifo_data),
    .irq_fifo_data_valid(rxunit_irq_fifo_data_valid),
    .irq_fifo_irq_valid(rxunit_irq_fifo_irq_valid));
  assign n176_o = {rxunit_spm_wdata, rxunit_spm_wr, rxunit_spm_en, rxunit_spm_addr};
  assign n178_o = {rxunit_config_wdata, rxunit_config_wr, rxunit_config_en, rxunit_config_addr};
  /* ni/network_interface.vhd:360:31  */
  assign irqfifo_n188 = n195_o; // (signal)
  /* ni/network_interface.vhd:362:32  */
  assign irqfifo_n189 = irqfifo_irq_irq_sig; // (signal)
  /* ni/network_interface.vhd:363:34  */
  assign irqfifo_n190 = irqfifo_irq_data_sig; // (signal)
  /* ni/network_interface.vhd:354:9  */
  irq_fifo irqfifo (
    .clk(clk),
    .reset(reset),
    .config_addr(n191_o),
    .config_en(n192_o),
    .config_wr(n193_o),
    .config_wdata(n194_o),
    .sel(irq_if_fifo_sel),
    .irq_data_fifo_data_valid(irq_fifo_data_valid),
    .irq_irq_fifo_data_valid(irq_fifo_irq_valid),
    .irq_data_fifo_data(irq_fifo_data),
    .config_slv_rdata(irqfifo_config_slv_rdata),
    .config_slv_error(irqfifo_config_slv_error),
    .irq_irq_sig(irqfifo_irq_irq_sig),
    .irq_data_sig(irqfifo_irq_data_sig));
  assign n191_o = config[13:0];
  assign n192_o = config[14];
  assign n193_o = config[15];
  assign n194_o = config[47:16];
  assign n195_o = {irqfifo_config_slv_error, irqfifo_config_slv_rdata};
  /* ni/network_interface.vhd:378:32  */
  assign spmbus_n202 = n206_o; // (signal)
  /* ni/network_interface.vhd:379:39  */
  assign spmbus_n203 = n208_o; // (signal)
  /* ni/network_interface.vhd:373:9  */
  spm_bus spmbus (
    .clk(clk),
    .reset(reset),
    .spm_slv_rdata(n204_o),
    .spm_slv_error(n205_o),
    .tx_spm_addr(n210_o),
    .tx_spm_en(n211_o),
    .tx_spm_wr(n212_o),
    .tx_spm_wdata(n213_o),
    .rx_spm_addr(n214_o),
    .rx_spm_en(n215_o),
    .rx_spm_wr(n216_o),
    .rx_spm_wdata(n217_o),
    .spm_addr(spmbus_spm_addr),
    .spm_en(spmbus_spm_en),
    .spm_wr(spmbus_spm_wr),
    .spm_wdata(spmbus_spm_wdata),
    .tx_spm_slv_rdata(spmbus_tx_spm_slv_rdata),
    .tx_spm_slv_error(spmbus_tx_spm_slv_error));
  assign n204_o = n78_o[63:0];
  assign n205_o = n78_o[64];
  assign n206_o = {spmbus_spm_wdata, spmbus_spm_wr, spmbus_spm_en, spmbus_spm_addr};
  assign n208_o = {spmbus_tx_spm_slv_error, spmbus_tx_spm_slv_rdata};
  assign n210_o = tx_spm[13:0];
  assign n211_o = tx_spm[15:14];
  assign n212_o = tx_spm[16];
  assign n213_o = tx_spm[80:17];
  assign n214_o = rx_spm[13:0];
  assign n215_o = rx_spm[15:14];
  assign n216_o = rx_spm[16];
  assign n217_o = rx_spm[80:17];
  /* ni/network_interface.vhd:389:41  */
  assign configbus_n220 = n232_o; // (signal)
  /* ni/network_interface.vhd:392:35  */
  assign configbus_n221 = n238_o; // (signal)
  /* ni/network_interface.vhd:394:41  */
  assign configbus_n222 = configbus_tdm_ctrl_sel; // (signal)
  /* ni/network_interface.vhd:396:42  */
  assign configbus_n223 = configbus_sched_tbl_sel; // (signal)
  /* ni/network_interface.vhd:398:40  */
  assign configbus_n224 = configbus_dma_tbl_sel; // (signal)
  /* ni/network_interface.vhd:400:40  */
  assign configbus_n225 = configbus_mc_ctrl_sel; // (signal)
  /* ni/network_interface.vhd:402:46  */
  assign configbus_n226 = configbus_irq_unit_fifo_sel; // (signal)
  /* ni/network_interface.vhd:384:9  */
  config_bus configbus (
    .clk(clk),
    .reset(reset),
    .ocp_config_m_mcmd(n227_o),
    .ocp_config_m_maddr(n228_o),
    .ocp_config_m_mdata(n229_o),
    .ocp_config_m_mbyteen(n230_o),
    .ocp_config_m_mrespaccept(n231_o),
    .supervisor(supervisor),
    .config_unit_addr(n234_o),
    .config_unit_en(n235_o),
    .config_unit_wr(n236_o),
    .config_unit_wdata(n237_o),
    .tdm_ctrl_rdata(n240_o),
    .tdm_ctrl_error(n241_o),
    .sched_tbl_rdata(n243_o),
    .sched_tbl_error(n244_o),
    .dma_tbl_rdata(n246_o),
    .dma_tbl_error(n247_o),
    .mc_ctrl_rdata(n249_o),
    .mc_ctrl_error(n250_o),
    .irq_unit_fifo_rdata(n252_o),
    .irq_unit_fifo_error(n253_o),
    .ocp_config_s_sresp(configbus_ocp_config_s_sresp),
    .ocp_config_s_sdata(configbus_ocp_config_s_sdata),
    .ocp_config_s_scmdaccept(configbus_ocp_config_s_scmdaccept),
    .config_addr(configbus_config_addr),
    .config_en(configbus_config_en),
    .config_wr(configbus_config_wr),
    .config_wdata(configbus_config_wdata),
    .tdm_ctrl_sel(configbus_tdm_ctrl_sel),
    .sched_tbl_sel(configbus_sched_tbl_sel),
    .dma_tbl_sel(configbus_dma_tbl_sel),
    .mc_ctrl_sel(configbus_mc_ctrl_sel),
    .irq_unit_fifo_sel(configbus_irq_unit_fifo_sel));
  assign n227_o = n71_o[2:0];
  assign n228_o = n71_o[34:3];
  assign n229_o = n71_o[66:35];
  assign n230_o = n71_o[70:67];
  assign n231_o = n71_o[71];
  assign n232_o = {configbus_ocp_config_s_scmdaccept, configbus_ocp_config_s_sdata, configbus_ocp_config_s_sresp};
  assign n234_o = config_unit_master[13:0];
  assign n235_o = config_unit_master[14];
  assign n236_o = config_unit_master[15];
  assign n237_o = config_unit_master[47:16];
  assign n238_o = {configbus_config_wdata, configbus_config_wr, configbus_config_en, configbus_config_addr};
  assign n240_o = tdm_ctrl[31:0];
  assign n241_o = tdm_ctrl[32];
  assign n243_o = sched_tbl[31:0];
  assign n244_o = sched_tbl[32];
  assign n246_o = dma_tbl[31:0];
  assign n247_o = dma_tbl[32];
  assign n249_o = mc_ctrl[31:0];
  assign n250_o = mc_ctrl[32];
  assign n252_o = irq_if_fifo[31:0];
  assign n253_o = irq_if_fifo[32];
endmodule

module noc_node
  (input  clk,
   input  reset,
   input  supervisor,
   input  run,
   input  [2:0] proc_m_MCmd,
   input  [31:0] proc_m_MAddr,
   input  [31:0] proc_m_MData,
   input  [3:0] proc_m_MByteEn,
   input  proc_m_MRespAccept,
   input  [63:0] spm_s_rdata,
   input  spm_s_error,
   input  north_in_f_req,
   input  [34:0] north_in_f_data,
   input  east_in_f_req,
   input  [34:0] east_in_f_data,
   input  south_in_f_req,
   input  [34:0] south_in_f_data,
   input  west_in_f_req,
   input  [34:0] west_in_f_data,
   input  north_out_b_ack,
   input  east_out_b_ack,
   input  south_out_b_ack,
   input  west_out_b_ack,
   output master_run,
   output [1:0] proc_s_SResp,
   output [31:0] proc_s_SData,
   output proc_s_SCmdAccept,
   output [13:0] spm_m_addr,
   output [1:0] spm_m_en,
   output spm_m_wr,
   output [63:0] spm_m_wdata,
   output [1:0] irq,
   output north_in_b_ack,
   output east_in_b_ack,
   output south_in_b_ack,
   output west_in_b_ack,
   output north_out_f_req,
   output [34:0] north_out_f_data,
   output east_out_f_req,
   output [34:0] east_out_f_data,
   output south_out_f_req,
   output [34:0] south_out_f_data,
   output west_out_f_req,
   output [34:0] west_out_f_data);
  wire [71:0] n1_o;
  wire [1:0] n3_o;
  wire [31:0] n4_o;
  wire n5_o;
  wire [13:0] n7_o;
  wire [1:0] n8_o;
  wire n9_o;
  wire [63:0] n10_o;
  wire [64:0] n11_o;
  wire [35:0] n13_o;
  wire n15_o;
  wire [35:0] n16_o;
  wire n18_o;
  wire [35:0] n19_o;
  wire n21_o;
  wire [35:0] n22_o;
  wire n24_o;
  wire n26_o;
  wire [34:0] n27_o;
  wire n29_o;
  wire [34:0] n30_o;
  wire n32_o;
  wire [34:0] n33_o;
  wire n35_o;
  wire [34:0] n36_o;
  wire [34:0] ip_to_net;
  wire [34:0] net_to_ip;
  wire ni_master_run;
  wire [1:0] ni_ocp_config_s_sresp;
  wire [31:0] ni_ocp_config_s_sdata;
  wire ni_ocp_config_s_scmdaccept;
  wire ni_data_irq;
  wire ni_config_irq;
  wire [13:0] ni_spm_addr;
  wire [1:0] ni_spm_en;
  wire ni_spm_wr;
  wire [63:0] ni_spm_wdata;
  wire [34:0] ni_pkt_out;
  wire [2:0] n38_o;
  wire [31:0] n39_o;
  wire [31:0] n40_o;
  wire [3:0] n41_o;
  wire n42_o;
  wire [34:0] n43_o;
  wire [63:0] n47_o;
  wire n48_o;
  wire [80:0] n49_o;
  wire [4:0] r_inport_b;
  wire [179:0] r_outport_f;
  wire [179:0] n53_o;
  wire n55_o;
  wire n56_o;
  wire n57_o;
  wire n58_o;
  wire [35:0] n61_o;
  wire [35:0] n62_o;
  wire [35:0] n63_o;
  wire [35:0] n64_o;
  wire [34:0] n65_o;
  wire [4:0] n68_o;
  wire [1:0] n69_o;
  assign master_run = ni_master_run;
  assign proc_s_SResp = n3_o;
  assign proc_s_SData = n4_o;
  assign proc_s_SCmdAccept = n5_o;
  assign spm_m_addr = n7_o;
  assign spm_m_en = n8_o;
  assign spm_m_wr = n9_o;
  assign spm_m_wdata = n10_o;
  assign irq = n69_o;
  assign north_in_b_ack = n15_o;
  assign east_in_b_ack = n18_o;
  assign south_in_b_ack = n21_o;
  assign west_in_b_ack = n24_o;
  assign north_out_f_req = n26_o;
  assign north_out_f_data = n27_o;
  assign east_out_f_req = n29_o;
  assign east_out_f_data = n30_o;
  assign south_out_f_req = n32_o;
  assign south_out_f_data = n33_o;
  assign west_out_f_req = n35_o;
  assign west_out_f_data = n36_o;
  assign n1_o = {proc_m_MRespAccept, proc_m_MByteEn, proc_m_MData, proc_m_MAddr, proc_m_MCmd};
  assign n3_o = n43_o[1:0];
  assign n4_o = n43_o[33:2];
  assign n5_o = n43_o[34];
  assign n7_o = n49_o[13:0];
  assign n8_o = n49_o[15:14];
  assign n9_o = n49_o[16];
  assign n10_o = n49_o[80:17];
  assign n11_o = {spm_s_error, spm_s_rdata};
  assign n13_o = {north_in_f_data, north_in_f_req};
  assign n15_o = n57_o;
  assign n16_o = {east_in_f_data, east_in_f_req};
  assign n18_o = n58_o;
  assign n19_o = {south_in_f_data, south_in_f_req};
  assign n21_o = n55_o;
  assign n22_o = {west_in_f_data, west_in_f_req};
  assign n24_o = n56_o;
  assign n26_o = n63_o[0];
  assign n27_o = n63_o[35:1];
  assign n29_o = n64_o[0];
  assign n30_o = n64_o[35:1];
  assign n32_o = n61_o[0];
  assign n33_o = n61_o[35:1];
  assign n35_o = n62_o[0];
  assign n36_o = n62_o[35:1];
  /* noc/synchronous/noc_node.vhd:95:8  */
  assign ip_to_net = ni_pkt_out; // (signal)
  /* noc/synchronous/noc_node.vhd:96:8  */
  assign net_to_ip = n65_o; // (signal)
  /* noc/synchronous/noc_node.vhd:102:1  */
  network_interface_5ba93c9db0cff93f52b521d7420e43f6eda2784f ni (
    .clk(clk),
    .reset(reset),
    .run(run),
    .supervisor(supervisor),
    .ocp_config_m_mcmd(n38_o),
    .ocp_config_m_maddr(n39_o),
    .ocp_config_m_mdata(n40_o),
    .ocp_config_m_mbyteen(n41_o),
    .ocp_config_m_mrespaccept(n42_o),
    .spm_slv_rdata(n47_o),
    .spm_slv_error(n48_o),
    .pkt_in(net_to_ip),
    .master_run(ni_master_run),
    .ocp_config_s_sresp(ni_ocp_config_s_sresp),
    .ocp_config_s_sdata(ni_ocp_config_s_sdata),
    .ocp_config_s_scmdaccept(ni_ocp_config_s_scmdaccept),
    .data_irq(ni_data_irq),
    .config_irq(ni_config_irq),
    .spm_addr(ni_spm_addr),
    .spm_en(ni_spm_en),
    .spm_wr(ni_spm_wr),
    .spm_wdata(ni_spm_wdata),
    .pkt_out(ni_pkt_out));
  assign n38_o = n1_o[2:0];
  assign n39_o = n1_o[34:3];
  assign n40_o = n1_o[66:35];
  assign n41_o = n1_o[70:67];
  assign n42_o = n1_o[71];
  assign n43_o = {ni_ocp_config_s_scmdaccept, ni_ocp_config_s_sdata, ni_ocp_config_s_sresp};
  assign n47_o = n11_o[63:0];
  assign n48_o = n11_o[64];
  assign n49_o = {ni_spm_wdata, ni_spm_wr, ni_spm_en, ni_spm_addr};
  /* noc/synchronous/noc_node.vhd:131:1  */
  router r (
    .clk(clk),
    .reset(reset),
    .inport_f(n53_o),
    .outport_b(n68_o),
    .inport_b(r_inport_b),
    .outport_f(r_outport_f));
  assign n53_o = {ip_to_net, 1'b0, n16_o, n13_o, n22_o, n19_o};
  assign n55_o = r_inport_b[0];
  assign n56_o = r_inport_b[1];
  assign n57_o = r_inport_b[2];
  assign n58_o = r_inport_b[3];
  assign n61_o = r_outport_f[35:0];
  assign n62_o = r_outport_f[71:36];
  assign n63_o = r_outport_f[107:72];
  assign n64_o = r_outport_f[143:108];
  assign n65_o = r_outport_f[179:145];
  assign n68_o = {1'b0, east_out_b_ack, north_out_b_ack, west_out_b_ack, south_out_b_ack};
  assign n69_o = {ni_config_irq, ni_data_irq};
endmodule

