-- 
-- Copyright Technical University of Denmark. All rights reserved.
-- This file is part of the T-CREST project.
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions are met:
-- 
--    1. Redistributions of source code must retain the above copyright notice,
--	 this list of conditions and the following disclaimer.
-- 
--    2. Redistributions in binary form must reproduce the above copyright
--	 notice, this list of conditions and the following disclaimer in the
--	 documentation and/or other materials provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDER ``AS IS'' AND ANY EXPRESS
-- OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES
-- OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN
-- NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY
-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF
-- THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation are
-- those of the authors and should not be interpreted as representing official
-- policies, either expressed or implied, of the copyright holder.
-- 


--------------------------------------------------------------------------------
-- A parameterized latch stage of the asynchronous noc.
--
-- Authors: Evangelia Kasapaki
--	    Rasmus Bo Sorensen
--------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.config_types.all;
use work.noc_defs.all;


entity link_pipeline is
  generic (
    -- direction: 0 north or south, 1 east or west
    constant DIRECTION : in integer := 1;
    -- disables the clock gating
    -- default: gating enabled
    constant GATING_ENABLED : integer := 0;

    -- for some cases a delayed request is needed
    -- default: request delay disabled
    constant GENERATE_REQUEST_DELAY : integer := 0;

    -- to fix hold violations: delay the acknowledge
    constant GENERATE_ACKNOWLEDGE_DELAY : integer := 0;

    -- initial state to implement
    constant init_token : latch_state := EMPTY_BUBBLE;

    -- initial data
    constant init_data : phit_t := (others => 'X')  -- Forced unknown
    );
  port (
    preset    : in  std_logic;
    left_in   : in  channel_forward;
    left_out  : out channel_backward;
    right_out : out channel_forward;
    right_in  : in  channel_backward
    );
end link_pipeline;


architecture struct of link_pipeline is
 
begin
 	  stage : entity work.channel_latch(struct)
	    generic map (
	      init_token => init_token,
	      init_data	 => init_data
	      )
	    port map (
	      preset	=> preset,
	      left_in	=> left_in,
	      left_out	=> left_out,
	      right_out => right_out,
	      right_in	=> right_in,
	      lt_enable => open
	      );
end struct;

